* LTspice Encrypted File
* 
* This encrypted file has been supplied by a 3rd
* party vendor that does not wish to publicize
* the technology used to implement this library.
* 
* Permission is granted to use this file for
* simulations but not to reverse engineer its
* contents.
* 
********************************************************************************
* ON Semiconductor T6 40V Standard Gate Model Library
* Release: Aug, 2020
* Model Version: 5.8
* Simulator: LTspice
* Process case: TYPICAL
*
********************************************************************************
* Model Contacts:
*    James Victory     James.Victory@onsemi.com
*    Scott Pearson     Scott.Pearson@onsemi.com
*    Ken He            kencanzhong.he@onsemi.com
*    Hyeongwoo Jang    Hyeongwoo.Jang@onsemi.com
*    Jie Bai           Jie.bai@onsemi.com
*    Kan Jia           Kan.Jia@onsemi.com
*
********************************************************************************
* Reversion History:
*	Vers.	Date		Brief Description
*	1.0		07/19/2017	1. Extract scalable base model from data of NVMFS5C450N. 
*                       2. Generated models for :NVMFS5C450N, NVMFS5C404N
*	1a		08/02/2017	Added NVMFS5C442N, NVMFS5C430N, NVMFS5C410N, NVMFS5C426N
*	2		03/14/2018	1. Added NVMFD5C446N, NVMFD5C462N, NVMFD5C466N, NVMFD5C470N
*						2. Fixed diode curve with ikfd=0
*	3		05/14/2018	1. Added NVD5C454N, NVD5C460N, NVD5C478N, NVD5C486N, NVMFS5C456N, NVMFS5C460N,
*						   NVMFS5C466N, NVMFS5C468N
*						2. Extracted thermal parameters using R in datasheet
*	4		06/21/2018	1. Added NTMFS5C426N, NTMFS5C410N, NTMFS5C404N
*						2. Extracted thermal parameters using R in datasheet
*   5       05/22/2019  1. Added NTMJS1D0N04C, NVMJS1D0N04C, NTTFS003N04C, NVTFS003N04C, NTMYS3D5N04C, NVMYS3D5N04C,
*						   NTMJS1D0N04C, NVMJS1D0N04C, NTTFS003N04C, NVTFS003N04C, NTMYS3D5N04C, NVMYS3D5N04C, 
*						   NTTFS004N04C, NVTFS004N04C, NTMYS5D3N04C, NVMYS5D3N04C, NTTFS005N04C, NVTFS005N04C, 
*						   NTMJS1D7N04C, NVMJS1D7N04C, NTMYS011N04C, NVMYS011N04C, NTTFS008N04C, NVTFS008N04C, 
*						   NTMJS1D3N04C, NVMJS1D3N04C, NTTFS015N04C, NVTFS015N04C, NTMTS0D4N04C, NVMTS0D4N04C, 
*						   NTMTS0D6N04C, NVMTS0D6N04C, NTMYS1D3N04C, NVMYS1D3N04C, NTMTS0D7N04C, NVMTS0D7N04C, 
*						   NTMFS5C406N, NVMFS5C406N, NTTFS002N04C, NVTFS002N04C 
*                       2. Update RGshield calculation
*                       3. Update diode reverse recovery model
*	5.1		10/18/2019	1. Update convergence capacitor
*	5.2		04/02/2020	1. Added NTMJS0D9N04C, NVMJS0D9N04C
*	5.3		04/28/2020	1. Added NVD5C434N, NVIS1D7N04C, NVIS1D9N04C
*	5.4		05/12/2020	1. Add NVIS1D5N04C, update NVIS1D7N04C
*	5.5		06/11/2020	1. Update Substrate mobility
*	5.6		08/27/2020	1. Improve temperature behavior
*   5.7     09/24/2020  1. Added NVMFSC0D9N04C
*	5.8		10/12/2020	1. Update thermal models for NTMFS5C426N_5P, NTMFS5C410N_5P, NTMTS0D7N04C_5P
********************************************************************************
* Usage:
* https://www.onsemi.com/pub/Collateral/AND9783-D.PDF
* https://www.onsemi.com/pub/Collateral/TND6330-D.PDF
* https://www.onsemi.com/pub/Collateral/TND6329-D.PDF
*
* This library contains 3 and 5 pin(or terminal) models. 
* The 3p models are isothermal with self-heating effects turned off.
* The 5p models are electro-thermal and contain 2 additional pins: 
* tj (or junction temperature)
* tcase (or device case thermal terminal).
* tj should always be left floating or can be connected to a very
* large resistor (>1meg). This terminal is meant to provide the user with
* output information on the junction temperature under operation. For model
* verification purposes against the data sheet and isothermal device simulations
* for example, tcase should be connected to a "E" voltage source with value {TEMP},
* the simulator ambient temperature. For system/module level simulations that
* include thermal effects, tcase should be connected to the device-module
* thermal interface node such as the heat sink interface point.
*
* In the case a designer wished to bypass the internal ZTH network, tj should be
* shorted to tcase and then tcase connected to the user defined ZTH network.
*
********************************************************************************
* Support devices:
*   NVMFS5C450N_3P, NVMFS5C450N_5P
*   NVMFS5C404N_3P, NVMFS5C404N_5P
*   NVMFS5C442N_3P, NVMFS5C442N_5P
*   NVMFS5C430N_3P, NVMFS5C430N_5P
*   NVMFS5C410N_3P, NVMFS5C410N_5P
*   NVMFS5C426N_3P, NVMFS5C426N_5P
*   NVMFD5C446N_6P, NVMFD5C446N_9P
*   NVMFD5C462N_6P, NVMFD5C462N_9P
*   NVMFD5C466N_6P, NVMFD5C466N_9P
*   NVMFD5C470N_6P, NVMFD5C470N_9P
*   NVMFD5C478N_6P, NVMFD5C478N_9P
*   NVD5C454N_3P,   NVD5C454N_5P  ;New 05/13/2018
*   NVD5C460N_3P,   NVD5C460N_5P  ;New 05/13/2018
*   NVD5C478N_3P,   NVD5C478N_5P  ;New 05/13/2018
*   NVD5C486N_3P,   NVD5C486N_5P  ;New 05/13/2018
*   NVMFS5C456N_3P, NVMFS5C456N_5P  ;New 05/13/2018
*   NVMFS5C460N_3P, NVMFS5C460N_5P  ;New 05/13/2018
*   NVMFS5C466N_3P, NVMFS5C466N_5P  ;New 05/13/2018
*   NVMFS5C468N_3P, NVMFS5C468N_5P  ;New 05/13/2018
*   NTMFS5C426N_3P, NTMFS5C426N_5P ; New 6/21/2018
*   NTMFS5C410N_3P, NTMFS5C410N_5P ; New 6/21/2018
*   NTMFS5C404N_3P, NTMFS5C404N_5P ; New 6/21/2018
*   NTMJS1D0N04C_3P, NTMJS1D0N04C_5P; New 05/14/2019 
*   NVMJS1D0N04C_3P, NVMJS1D0N04C_5P; New 05/14/2019 
*   NTTFS003N04C_3P, NTTFS003N04C_5P; New 05/14/2019 
*   NVTFS003N04C_3P, NVTFS003N04C_5P; New 05/14/2019 
*   NTMYS3D5N04C_3P, NTMYS3D5N04C_5P; New 05/14/2019 
*   NVMYS3D5N04C_3P, NVMYS3D5N04C_5P; New 05/14/2019 
*   NTTFS004N04C_3P, NTTFS004N04C_5P; New 05/14/2019 
*   NVTFS004N04C_3P, NVTFS004N04C_5P; New 05/14/2019 
*   NTMYS5D3N04C_3P, NTMYS5D3N04C_5P; New 05/14/2019 
*   NVMYS5D3N04C_3P, NVMYS5D3N04C_5P; New 05/14/2019 
*   NTTFS005N04C_3P, NTTFS005N04C_5P; New 05/14/2019 
*   NVTFS005N04C_3P, NVTFS005N04C_5P; New 05/14/2019 
*   NTMJS1D7N04C_3P, NTMJS1D7N04C_5P; New 05/14/2019 
*   NVMJS1D7N04C_3P, NVMJS1D7N04C_5P; New 05/14/2019 
*   NTMYS011N04C_3P, NTMYS011N04C_5P; New 05/14/2019 
*   NVMYS011N04C_3P, NVMYS011N04C_5P; New 05/14/2019 
*   NTTFS008N04C_3P, NTTFS008N04C_5P; New 05/14/2019 
*   NVTFS008N04C_3P, NVTFS008N04C_5P; New 05/14/2019 
*   NTMJS1D3N04C_3P, NTMJS1D3N04C_5P; New 05/14/2019 
*   NVMJS1D3N04C_3P, NVMJS1D3N04C_5P; New 05/14/2019 
*   NTTFS015N04C_3P, NTTFS015N04C_5P; New 05/14/2019 
*   NVTFS015N04C_3P, NVTFS015N04C_5P; New 05/14/2019 
*   NTMTS0D4N04C_3P, NTMTS0D4N04C_5P; New 05/14/2019 
*   NVMTS0D4N04C_3P, NVMTS0D4N04C_5P; New 05/14/2019 
*   NTMTS0D6N04C_3P, NTMTS0D6N04C_5P; New 05/14/2019 
*   NVMTS0D6N04C_3P, NVMTS0D6N04C_5P; New 05/14/2019 
*   NTMYS1D3N04C_3P, NTMYS1D3N04C_5P; New 05/14/2019 
*   NVMYS1D3N04C_3P, NVMYS1D3N04C_5P; New 05/14/2019 
*   NTMTS0D7N04C_3P, NTMTS0D7N04C_5P; New 05/14/2019 
*   NVMTS0D7N04C_3P, NVMTS0D7N04C_5P; New 05/14/2019 
*   NTMFS5C406N_3P, NTMFS5C406N_5P; New 05/14/2019
*   NVMFS5C406N_3P, NVMFS5C406N_5P; New 05/14/2019
*   NTTFS002N04C_3P, NTTFS002N04C_5P; New 05/14/2019 
*   NVTFS002N04C_3P, NVTFS002N04C_5P; New 05/14/2019 
************
*   NVMYS8D0N04C_3P, NVMYS8D0N04C_5P New 12/26/2019
*   NTMYS8D0N04C_3P, NTMYS8D0N04C_5P New 12/26/2019
*   NVMYS4D5N04C_3P, NVMYS4D5N04C_5P New 12/26/2019
*   NTMYS4D5N04C_3P, NTMYS4D5N04C_5P New 12/26/2019
*   NVTFWS002N04C_3P, NVTFWS002N04C_5P New 12/26/2019
*   NVMYS2D4N04C_3P, NVMYS2D4N04C_5P New 12/26/2019
*   NTMYS2D4N04C_3P, NTMYS2D4N04C_5P New 12/26/2019
*   NTMFS5C430N_3P, NTMFS5C430N_5P New 12/26/2019
*   FDBL9401_F085T6_3P, FDBL9401_F085T6_5P New 12/26/2019
*   FDBL9403_F085T6_3P, FDBL9403_F085T6_5P New 12/26/2019
*   NTMJS0D9N04C_3P, NTMJS0D9N04C_5P New 04/02/2020
*   NVMJS0D9N04C_3P, NVMJS0D9N04C_5P New 04/02/2020
*   NVD5C434N_3P, NVD5C434N_5P New 04/28/2020
*   NVIS1D7N04C_3P, NVIS1D7N04C_5P New 04/28/2020
*   NVIS1D9N04C_3P, NVIS1D9N04C_5P New 04/28/2020
*   NVIS1D5N04C_3P, NVIS1D5N04C_5P New 05/12/2020
*   NVMFSC0D9N04C_3P, NVMFSC0D9N04C_5P New 09/24/2020
********************************************************************************
*
* Begin:
 31 6B 4B FE 88 B3 ED A2 F8 66 30 06 10 BB C8 77
 F4 84 0C A0 CF AF D7 E4 92 92 45 B6 57 14 A4 9E
 BE C7 B0 7B 97 D3 AA 69 80 17 92 EA 2A 11 59 9B
 04 D8 F5 62 71 C5 DE 00 7C 40 96 DB 98 DE 42 C4
 F7 4D A7 60 E7 0C F4 52 C1 4C 9B A2 6E 75 70 2E
 7E F7 72 FA 6C C3 65 22 DC 91 98 84 DB 96 E6 CE
 5F 5F 81 89 76 A6 5B 69 F0 7A 88 FA 34 08 F9 82
 3D F3 F7 90 22 20 E2 C2 69 60 2D EE AA 49 45 28
 1E B0 1E 37 1E 72 77 06 E4 DE 6A 70 E8 CD 66 8F
 BC 46 54 08 57 2A D5 D5 12 5C 22 DE BB 17 BD 68
 A3 B0 9F 0A D9 81 49 E2 74 43 61 53 09 26 82 53
 A3 1B 82 97 F4 87 B0 02 34 9B A9 09 18 08 9A 54
 03 1F A4 0D 07 B3 50 83 27 C5 F9 33 F7 9A 08 CB
 32 8C 20 41 8C 55 CD 9F C2 36 ED B5 9E 51 40 AB
 7D 24 FF 2E BA 92 E0 3E 01 FC 28 AB 84 8B 99 E2
 C6 44 92 ED 2C C1 6D 19 83 06 15 C9 4A 1A F7 36
 88 6F 02 2A 25 09 13 AA 9A 6C A5 ED 61 54 C4 B1
 CF D0 C8 A0 53 80 B1 E7 DA B1 7C 9D 98 23 75 88
 B4 46 CB 48 A4 E8 DB 6E 0A D0 4F 5F DF A4 97 67
 91 B3 84 3C F9 43 E4 FE 23 86 07 D5 22 73 80 8C
 FD 00 B6 70 76 37 76 0F 55 47 C0 39 B3 FF 8D 4E
 30 99 98 B3 86 6E 27 B7 39 1C 44 F8 0C 5C FC 7A
 B5 8E CA 83 C1 D7 B0 57 5F 28 4B B3 A2 31 7E 32
 D4 F1 D4 B0 D1 43 E5 57 6E FF 41 2E 0D 47 FE DA
 8B 7B E1 8A 15 52 3E E7 F9 B3 3D 77 AB 46 98 EB
 8E 69 BA 67 DC 2B E3 34 A9 D4 4E 4E B4 B3 8E CD
 13 38 00 17 32 10 DD 6F B8 80 69 D7 6E 02 35 68
 B2 80 57 01 EA 1E 41 7A 29 7D 84 DC C3 D8 18 E8
 27 49 62 51 BD B6 EF 3A 73 17 18 8F FD 5E B4 F3
 F1 C2 10 6D 0F 82 37 3B 0A BE 69 84 8D 96 B6 74
 4E 8D 8A 06 4C 97 95 A1 EA 38 8B D5 AD CA 7F 31
 B9 A4 40 F6 54 F7 2E 2A 81 F3 E4 3C F9 68 58 15
 B2 FD 04 09 33 93 2C 11 CE FD 38 9D 62 EC EA 05
 B5 A7 F4 4E 8D 85 04 E6 11 55 ED D4 6B 19 C0 62
 A6 74 04 53 7E 78 B3 93 49 40 F8 37 CF C0 9F A0
 CD AC 3F 07 09 12 77 1D 71 34 5F C0 9D E6 E8 09
 C5 F6 74 8E B6 51 CD 62 6B A1 18 E4 24 F3 74 32
 1B 24 4B CF DE 1E 81 F3 9A 95 B5 E9 0C A2 19 CC
 D3 AC 21 B0 1F E0 39 42 CE A1 3B 15 40 F6 01 D5
 6A 5E 98 C8 9A 41 3E D2 92 DC FC DE 1F A3 A8 8F
 EB FD 8E AA AC 75 57 B2 AC D4 4C 79 5F D7 A3 29
 2D 05 A6 2C 1D 1F 48 64 93 1E 42 09 EA E5 9C AF
 DA 63 25 5D E6 4C CD B9 18 FB A7 38 E3 DE 1F 0E
 6C A4 0A F8 1C 85 47 3E 26 60 B2 13 F9 DB 3B 5F
 CE 86 47 41 90 1F 8F 81 E1 10 F3 EE 4E 07 34 37
 82 0B FC 4E 61 35 0D 66 7F BB 79 A4 68 85 06 76
 F9 95 20 9D 28 D1 B3 A8 04 F9 DD 63 3D AE B0 FC
 AC 6B 6D D9 F3 7E 0B 0F 8A 87 EF 1F 1A A7 FF 13
 8A CD 42 0A 6C 0B 30 E3 1E C5 AB C1 9F 25 54 6E
 B7 84 56 00 08 AC 9B F1 90 84 7D F6 89 C7 20 05
 31 5F 7B EA 92 73 CB B9 8C 0C 5C 93 B5 2B B9 5F
 3F 81 85 A3 24 17 96 AD 6A 26 7C 56 D1 66 DC 3C
 3D 76 D1 EE BE C6 26 4D CA 8F 86 22 E0 E4 B8 87
 F7 3F 78 C5 20 F7 30 DA 63 64 8E 4F 6C 56 39 D6
 F3 22 36 35 B8 D5 2C 63 0F C0 92 13 03 21 15 38
 36 8F 81 2B BC 45 B3 E8 8E 55 07 91 73 6D E6 54
 38 AB EC 87 CF 8A F1 DC 8D 41 FD C5 D6 8C F7 19
 59 26 A0 68 2B 97 19 82 3B B1 44 ED 6A B0 FA A2
 DC 6D D6 B3 2A C5 81 C6 A1 FB BC 0A AD D2 5C 6F
 73 3B BC 5F AF 28 93 74 C5 81 7A 38 5A FE 72 2B
 B0 F8 2A 21 6D 1C A8 5E 47 59 98 D9 98 32 B2 A4
 47 C6 A6 50 13 DC 98 E7 71 F6 E8 47 89 DA 1D 49
 A1 A9 61 A4 91 5D E5 B7 E9 F0 83 2A B6 B1 B4 6A
 54 B6 66 FD 75 8E 26 9C 68 31 CD 39 2D 9F 5A 8F
 F3 89 26 0F 0E 66 41 68 EA 94 84 46 DD 55 7A 54
 4A 32 40 4E 4C 33 20 83 B2 8A A0 8E 7F 77 72 65
 78 7B 07 5B 43 EE 96 E6 24 3B 9D 06 60 5C 99 FA
 AB AC EB 7B 5F 53 9D FC DE D4 A5 86 47 B3 FF 0C
 D3 39 38 5B D3 C2 27 B4 63 62 DE 1D 0F 05 96 17
 45 54 31 51 99 46 D2 01 1C 24 F2 D2 75 58 57 31
 03 F6 2C 4E 5C 87 AD 8C 42 31 C1 B0 0D D1 30 3A
 6E D3 72 FA 28 6A 79 75 79 FA CA 93 14 C2 D3 29
 DA F9 D5 17 2C B8 D6 5E 57 42 41 EA 5B 8C B3 A7
 F3 09 83 E5 9F 9A 44 CA 98 F0 51 AF 65 EF F3 47
 BA 8A 28 AC 81 50 A3 3E 3E 11 AF 97 E1 43 67 E4
 C9 74 E7 4E C0 D2 9F 0D FF F2 B3 2F 7F 74 55 B9
 ED 57 66 38 04 D7 BB 45 50 9C 52 96 C6 C0 54 B3
 C7 F6 5E A1 5A 9E 34 8B 72 F0 94 44 78 AE 05 C4
 E1 5E D6 CD 30 18 58 0C C2 8E A0 6B 61 30 A0 9A
 3C E6 44 42 F2 A6 C1 E2 68 A7 BC 61 5F EF 52 1F
 0B C3 25 D6 BB B2 27 74 FF B9 59 F2 96 14 1B E1
 56 D7 37 C8 31 73 1B 27 D0 45 FA 8B 35 77 A0 EC
 D7 2B D3 4D 3A 08 AD 3D B8 95 D6 D6 28 74 A3 24
 90 91 A1 A4 BA 73 22 00 BB B0 C1 88 32 46 93 1E
 9B 48 EC 0B 37 CB 20 BA B4 0C AE D2 D6 7F 69 7A
 DA CE 1E D9 2F D4 08 E8 DB 78 AD FB 95 A6 CD 23
 04 8B 77 3E 0A 3A 69 08 C0 D6 ED 0D 62 38 EB 33
 73 3F D1 CC F2 18 9B 1E 27 99 C5 53 CC 98 39 9E
 40 A4 59 45 B3 03 43 16 96 66 A4 3C 4B 5D 96 68
 EC E8 A5 A0 61 A7 BD F6 CA 76 2C 42 F6 90 DE C3
 DF 67 70 86 91 6C E1 2C 4A F2 E4 FF B3 EB D3 5F
 9C F3 CE 4F 2B CD 1F AF 07 86 6E A5 0E 69 10 A8
 63 6C 5A 24 D9 14 BC 70 63 C7 52 7F 30 A0 1A 4C
 35 B2 03 0C 97 68 C4 55 9D 93 0E A6 9C B5 66 48
 98 94 DB 08 56 1E D4 9A 03 97 E9 9D C3 AF E5 A9
 DD FA DA C4 DF 1B 44 B4 0C 62 77 86 00 4A 91 EF
 22 2F B6 70 EF 1A A7 E2 FB 6B 43 68 77 9A 5E C9
 50 44 DE 25 38 84 A2 A0 80 0D 95 14 42 D8 21 CD
 60 C8 EB 0F AC F0 0C EA 2A 2F 63 58 1A 1D 2E 2C
 1A 85 89 51 15 F8 AE 92 D8 BF E4 28 A3 33 B4 C8
 B0 E9 CE 49 94 53 C8 88 78 F2 26 79 0F 16 FD D5
 2A AA D2 A0 51 EF C2 8F 5C 1D 23 70 CD D6 C9 21
 A2 6B 9F 2E 36 6F E4 DB B5 B2 B3 D9 A9 53 8C AF
 B2 36 F5 5B 1C 41 2F 46 BB BB 60 46 21 FF 80 70
 81 04 87 14 AB AA 4C 6B A8 8B 24 01 1A 1C 4B 7D
 34 20 DF 79 0F 14 AC DA 8E 7B 9A A1 E6 C7 F0 BF
 64 AC 4D 8F 35 33 1C 15 35 53 0B 9C 6A 73 E4 C4
 AD C2 15 8E 50 66 80 50 A9 7E EF 1D E9 5C D1 63
 ED 73 92 AA C1 2B 2E FE 12 F1 79 C6 1B 32 38 8C
 08 37 C0 96 4A 1A 07 8F 27 47 3C 9C 7A 0E 34 1E
 55 4A 8B 88 AD EE B9 EE 17 C4 3B C0 0C 52 46 FE
 19 4F 5C 74 07 42 EA 72 54 35 9B 27 B9 58 3D 11
 1F 8E 45 7B 97 04 7A 33 9F 54 77 93 CB 1A FF 89
 21 12 50 18 CA 54 84 5F 80 1D 75 59 A1 A9 9D 3F
 9B F0 56 3A 28 BE A9 BA 41 BB 2F 8E 0B 98 BF 66
 68 9E 3F 52 CE 80 CD 06 1A 00 71 BF 41 80 DB 00
 FE 26 4F AD 04 04 D4 BD E8 23 FC A8 64 CA EB 79
 ED AC B9 04 EB BE 8B 19 30 0B F1 7F CA BA 9A B1
 A8 CD D3 A0 CA EE D9 91 34 B8 8E 06 78 DF 33 29
 33 05 7A 8E D0 E8 66 F2 05 C6 6C 87 1E A9 7C D7
 58 92 C1 17 EC 76 FE F8 72 75 52 D3 D6 AD 9D 08
 54 F1 03 FA 8F 29 36 0B 22 7F 84 B0 AE 15 F5 73
 F0 90 4B C0 DB A1 F6 CF C5 F6 A6 D3 ED 83 2D 20
 45 ED 0B 34 C6 C4 0D 40 3F 4B A7 55 6D BE DF F5
 A1 B9 55 28 64 C8 3E C2 9E 6F F4 D8 72 B2 46 B8
 12 7B 81 67 6F 98 51 46 E5 56 C4 62 4D 97 F2 94
 46 FC 7F 45 60 15 05 09 B6 B7 60 15 0A D8 4A 21
 AC B3 38 22 C6 1A FB 53 EE AE 1C FC 47 8D DC CC
 EB E0 2A 4D 35 AF 3E F7 A2 92 32 79 0D 06 26 1D
 78 BF EC 54 D7 AD 0A 78 0E 85 5F 4A 9F C0 BE FA
 6C BC 81 9D C1 E4 7A 0F F7 2B A8 76 4F BA 8C 4F
 4B 2F 83 AC BE EB 42 48 B4 37 05 5A CC 07 B8 A5
 8A 06 23 91 47 FA 64 5E AE 79 F8 93 59 FF 26 50
 67 BD 27 AD 5A 56 2E 27 FF 5F 5F D6 6E A3 2C 6B
 6F 27 54 F4 D9 06 D0 87 0B 33 01 83 0A F0 2B 87
 FD 3C 2A 3D 9C 74 58 00 68 63 DA FC 4D 4C 47 46
 E9 1D 75 9E 4F D4 C0 BD B3 70 3C 68 F4 C1 80 63
 87 F0 C7 E2 90 22 74 77 75 34 39 08 F3 A3 83 D6
 2A 62 05 E3 CC E5 40 9D 9D 2B 96 28 4A 1F 79 8E
 7D 6C 80 A3 F2 1E A4 40 3F 1D 76 06 30 2F B2 75
 21 80 1E 08 B8 BE 50 1D 86 2C 6C 82 D6 5D D9 A3
 E9 2C 6A 82 31 32 BB A3 83 3D 3F 5A 4B 10 40 E4
 2E 87 0F AC 02 C8 51 63 F3 70 FF C5 3A 15 08 C1
 E9 19 FB 6D 45 03 AC 64 AA 25 6D 94 FD 87 00 CD
 68 9F 41 60 DA A7 18 F6 D8 62 78 8F 9C 01 97 16
 6C 0F A3 CB C9 A5 DA FC F4 8A FD 11 95 B1 19 DF
 D7 C9 8D 41 D1 AB 99 40 03 93 24 FF FB D4 49 08
 8B DB 3B E9 FA 36 25 0B 14 DF 9C 8E 7E 86 F6 6B
 6D 11 DA D2 71 C8 B0 84 21 8F C8 59 7D DE 22 8E
 07 21 C2 93 45 50 2B 6B 54 41 87 40 26 81 5A BB
 C9 F4 21 DF 90 CC EC 65 68 99 90 CE CB 83 A5 60
 1E 5D 07 61 88 AB 51 20 6A 15 10 71 26 87 B4 A2
 81 4A FE C6 3D A7 96 57 16 82 EE 76 72 68 02 28
 F6 D4 2F 81 75 35 1B A3 18 15 E1 CE A4 D2 F3 08
 4D AC 9C BD 10 45 EA B9 F3 0D 02 0E 2B C0 E8 44
 CF 5F 15 CE 64 66 EA DF 00 47 E4 2C B8 D6 58 DF
 67 07 52 EF F2 4B 57 6A 08 04 49 71 C2 73 F2 EC
 5E 1C ED 3D 5C 05 C1 42 9B B5 52 7E 8F 7F 7C 43
 B3 AE ED DD FA CC 8D 0E 31 86 AA 02 36 76 E6 8D
 1F 8F 75 4F BC 4D 31 EB 77 F4 DB 92 99 68 EE 62
 3A 65 F2 DD 87 4B 46 FD 9A 1F 5C EB 30 0F 66 3E
 78 F2 36 40 E1 A4 45 18 5A F9 72 B0 55 3E C7 55
 8E 02 88 A3 1E BF 7D B8 C5 25 E2 31 56 81 5E 33
 8E 71 00 9D A3 53 E9 4E 16 F1 58 BD 31 86 19 63
 65 A5 95 D5 7D 4E BD AD 3E EC F1 20 06 B9 D8 FA
 3E 79 FA 35 1C 8E DD CB 3C 84 77 2A 73 1B 55 55
 CF D3 E2 85 9B 40 37 4C 2F 43 7F 9F E9 59 E5 0D
 94 8D 0D 2C C5 49 A3 A9 A7 22 04 8A 92 F6 35 1B
 13 82 B4 41 8A 66 4F 95 DB F0 2A BB C9 F4 D1 4F
 12 1D FA 30 F1 9F 8A 18 56 72 98 98 52 CE C7 1C
 A3 9A F9 57 17 D8 EA 67 8F 55 7B A5 F2 D8 9E F8
 B9 FD DC 27 FE 80 16 E5 86 5A E5 B3 86 03 7B 2D
 CB 13 D0 BB 4D AB 6B 4C D1 24 AB A6 46 B2 2C E0
 6E 5C 96 C8 7E B7 79 20 49 B6 AA 9D E5 FA EB 2C
 A7 B8 3A CA 07 EE FB 88 2D 0F 8E 4D 8E 00 41 9D
 23 52 A8 C8 37 9F 49 42 66 FE FD 87 1A C9 9A 90
 98 6B 78 61 EF 83 2A F9 A5 78 CF 61 77 94 EC 6C
 D4 28 54 F9 02 9C 7A 9E AA 1A 7C FD 5C A6 A0 9E
 D4 E2 EF 35 19 1A 69 8A C6 9F 77 92 0E DB 14 ED
 6E 89 F8 B3 9E 09 8F 79 D4 CA CB 57 C9 7A AA 3B
 9F 54 D6 C9 09 AE E2 21 C5 BB E4 34 8E 35 AA A3
 1E 8C 94 96 05 FB 4E 12 48 C2 D7 BD 15 72 42 A2
 6B 5D 3C 32 53 93 6C 56 CD 63 15 E2 57 DD DE 31
 9F E8 F1 CA 48 E3 73 6F 52 94 E5 F6 F4 D6 86 5B
 2D 3B 99 62 E2 76 82 52 3F 06 13 14 5F 40 34 A2
 1E 4B 14 CE 73 1B B8 D8 4F 8C EF 57 32 71 D1 A5
 EB 9F D0 F5 18 77 8B F6 2F AC 09 13 42 F9 DB 46
 EC 13 41 E1 A2 EB 50 8D 4D 22 C0 DC CB 6D 76 05
 5D 11 E9 15 53 FD C8 1D A1 51 23 95 EA E3 9C 29
 28 E5 E8 7C CE 08 26 AD B6 8E 2D 24 9C F7 93 83
 01 C5 B5 C0 B7 96 4B B8 FD D5 18 8E 43 49 83 60
 6C 6D 90 26 FA 66 E1 89 F3 E0 78 83 93 DE 75 3A
 E7 EA A3 7E 02 CB DD 5E 62 02 4B 30 AA 55 A9 B7
 67 49 8A F1 86 F0 75 64 20 DF 6D 78 39 77 E6 95
 EA EF E2 F7 2D B3 A4 DD C9 E1 17 74 D6 4E A2 61
 AC C0 4B AA 73 53 5B 1F F3 B0 82 B5 7F 3F C7 D0
 09 3A 1F 38 9D 1D B8 F8 73 8A DF B9 80 35 82 8E
 0D 8A EF 98 55 A1 46 29 8F 83 B2 17 94 74 16 6C
 9F 10 83 A7 56 99 33 B5 5C F6 D6 51 27 C1 4C 7D
 BC 54 CD FF 2B 2B 1A 56 83 04 FC EC B8 37 07 6B
 06 05 38 D2 26 EC B9 7E 24 01 40 82 73 9E 68 35
 7A AB 24 EC 8C 34 E3 8A 21 CD 47 7F 71 C3 54 8E
 2A B7 B6 AB 20 D5 F7 31 4B 73 78 D8 F8 37 0E 2A
 26 8B E9 65 50 C2 A1 4E 8C 2B C0 9A B2 A9 FA 97
 91 1C 4F 02 04 75 3A D9 97 F9 66 E3 EB 5C F0 32
 9C B0 9A BA 6F 94 99 17 F1 7C 51 2B 6B A0 EE 90
 EA BE 23 20 BE CF 5B 25 61 1D 5B FF B9 84 97 D0
 A3 F4 13 8A 1F A3 13 BD 9F 11 64 E6 FD 8A A3 00
 1D EC F2 F7 5C FE 76 E7 0C F9 37 C1 AE D0 AD A4
 5E E1 45 C8 6E 83 F0 94 43 6B 75 64 DF 9F 07 19
 F5 EC 31 A2 46 3D CD 20 E8 F5 10 39 AF E6 1E 20
 02 83 25 72 E9 7D 86 FD E6 7B B1 05 0F 83 2F D6
 46 9A E6 60 97 07 91 16 74 31 69 C1 30 01 EA CA
 B1 36 61 F9 BE A0 0C 2B 82 29 F8 0C 2A 39 B7 DF
 C9 8C E3 E3 66 02 9B 2E A0 CA FC AA 1F E3 B7 F1
 01 18 36 57 80 A7 FC 40 8B DC BC C6 6A 4C 86 7A
 EC 11 29 A6 91 F1 85 79 05 4A 68 FA 89 71 3C C5
 F2 29 04 57 76 98 F6 25 7F C6 B4 BC 61 20 A1 58
 B0 AF EF 6B 99 B6 07 67 0C C4 4E 9E A9 08 7E 14
 45 32 F6 0D 34 58 17 E6 FD 8B AC 65 8D 74 14 10
 89 3F B0 8D D8 E1 9F 27 82 34 D2 61 D8 9E 2A 4A
 79 51 A3 BA 18 6C 55 40 92 7A 5E 56 CD E7 91 14
 98 F8 50 58 53 BC F7 FE E0 60 CD 50 80 65 D2 3A
 51 A1 EC F9 3B 51 11 7E 68 CE E8 7C C9 30 92 02
 FA AF 73 A6 B7 14 9E B7 0B 94 83 C5 55 24 87 73
 01 8F FB 2B D2 85 45 5E 02 41 E5 97 59 3C D3 05
 32 C9 92 41 EA 95 1C 7F BE EB E2 F1 BA A5 9B A8
 EA B0 BD CD A5 28 23 C0 4C AC F2 4C 51 AF 6B 38
 6A 4A BC 64 9F EB A3 19 E8 3F 7E 91 5D 58 83 86
 CA 5C 60 84 D5 22 1D A1 B4 A6 24 32 D9 87 2F B5
 FD C7 85 77 06 2C 5F 41 AE FA 9B 34 EA BE B7 1E
 AD 43 B1 31 8D 66 D9 BE 8F 0A E4 95 3F 30 8C E5
 EE EC 3B BE AF E1 F5 AA B6 1B 12 43 20 EC 07 80
 BB 4B ED 77 43 E1 70 88 C2 7A 1C 16 50 B0 DB C8
 EB B8 A6 24 6B 32 D3 6C BB 88 39 FF 91 EF 9E A6
 94 83 A1 5E 3D 02 94 0B 79 C0 93 71 F1 83 1F 3B
 10 49 D8 B5 F4 1D 64 D6 7E 24 FB 7A 6A 61 62 A7
 80 62 DF EA EA F4 0D BF 5E 46 E5 A2 8A E2 09 6A
 4E E6 21 A1 D1 49 3C 20 DB 89 4A 7A 77 61 8B FC
 79 AF C3 96 FA 1E E8 17 EC 25 76 98 45 85 1A 23
 E8 32 96 E1 DF A2 5B 90 99 24 98 0B 20 07 ED 8A
 8C BE D3 A8 4B F0 1A BE 0A 34 E9 85 08 78 B2 0E
 EE E2 4E DA 8B 64 65 80 63 12 99 DC A5 03 F2 26
 CE 48 56 89 28 60 8F 46 CC A5 E0 46 1A D4 F8 B9
 74 14 76 2A C3 77 BB F8 5D 3A 23 E7 15 A7 6C 6A
 F1 DE 16 94 F5 64 E8 B7 EC 0F DE AA D4 F2 32 E2
 5A 1B D5 8C 63 A1 E1 05 52 AB 8E 2D EE 2D 4F 89
 49 7C A2 E5 BB FE A4 8D 7B 2B 5B 86 99 BB CE 98
 13 A9 84 F4 12 03 07 89 51 D5 0F DE 04 20 71 E9
 5C FF 66 41 61 28 D0 DF EC 89 E0 72 A2 A8 6A 02
 C1 4F 2A 51 26 74 BC 7E EF DE BF FE AB 28 CA 8B
 D2 C1 EC C4 0E 57 3B E4 BF 91 36 AA B0 69 E5 54
 32 F8 F7 46 C8 71 24 E7 55 37 17 37 02 BD FB CA
 19 7A 5C 5C 7F FF 46 AE 46 75 77 25 5C 28 45 DB
 FD 9B 80 82 85 8E 60 E1 0C FB 99 31 5B 47 8C 79
 88 71 2D AA 0C FA 6C B1 2D B9 B6 54 4C 46 0A 2E
 38 59 10 D0 F9 93 A3 DD 7B 1C 76 A0 A7 58 6F 37
 F3 42 5F B2 C2 E1 0C 2E 9E 1A 9C 7D AB F9 D7 F6
 84 CC 2B 92 02 3A BC A4 4E 60 D0 92 38 16 13 72
 B8 00 C7 3F 29 2B CC 29 C0 91 C2 EE C3 0F 78 37
 B3 E8 1D 6D 27 67 3E 50 D6 E3 D3 52 56 45 97 A5
 F3 8A 83 46 27 3A C5 3D 9D F7 62 6F E0 2B F6 85
 F3 7C 50 5D 86 13 2D 91 FD 5D A9 B7 CB 8E 58 D7
 8C 02 5C 38 A4 35 78 94 D4 B1 2C 3E DB 23 50 4B
 83 B6 B0 78 A8 4C B3 64 28 FA 3E 76 D6 90 B1 B0
 FA 50 12 65 2F AC 39 32 63 6F CF 2B 3C 1F F3 12
 86 9A 38 E2 18 0D C9 1A 92 FF B2 76 32 81 4B 11
 9C 40 CF 02 06 CF F4 E8 E7 06 3B ED D6 AE 0B 2C
 7E 51 52 70 C1 F7 15 B2 31 96 3C 0B 99 C4 03 0B
 AC 91 F3 DE 83 DC 50 D7 06 55 0D BD 1B 69 CD EE
 D9 D8 75 7B DE 94 13 35 48 21 67 83 EA 19 33 1D
 4D 99 D0 0A F2 D1 7D B2 FC D1 59 5C AE A0 BD A3
 36 C4 96 DF B4 C3 AD 70 E3 7A 01 CD 85 E7 10 CC
 20 89 A1 95 89 42 77 5D 02 DE D4 62 12 B9 53 AA
 62 5F 7E 8F 6D 42 EC B7 85 71 80 F8 15 DB 06 FD
 7B CC AA 6D A1 A4 2F 37 67 8E 70 CA CF 73 3D EC
 51 FD 02 34 CC 42 7F 6F 51 86 48 6F 34 2B D7 83
 E9 A4 BE 44 B1 6A D3 82 D1 6E 58 60 81 A8 5F 86
 8C 2F 66 A2 BE 7A 6E 78 27 C3 E3 E5 01 5E 5E 3C
 F2 A6 AD 30 C9 38 AC 86 39 F3 20 1C 06 DE 67 81
 91 BB C0 8B CC 37 A7 23 96 78 36 D0 98 11 0E 80
 DE 42 0B DE AA 51 80 26 1F 33 9C C9 DF 93 51 EB
 D6 73 2B 68 FF 74 D9 3E 31 30 BF EA 61 94 20 22
 AA 51 70 58 B3 21 89 A8 1C 37 11 DE C8 E9 83 E4
 A5 2E 2F 15 5B EE DF 2F 91 50 03 D4 44 5A 19 25
 AB 46 77 D5 B5 87 0A ED 9D 72 B0 81 4E 4A A9 51
 5A CD 6E E1 6A 5C FF D5 8E 65 61 A2 B4 7B C4 C0
 43 4B B2 1D 1C 24 1E DB 78 6A 28 DA A9 12 14 2E
 DC DA 12 4D 23 49 40 BE BB 87 05 C9 70 10 F1 21
 31 A1 A4 53 6E 3D 21 2D 4B 99 DE E1 E7 58 E4 7F
 02 3E D6 49 C1 E4 E9 06 14 9F 56 CB 83 48 CA 33
 9D D0 73 20 0F 2E BD 63 AD 75 6F B0 98 D8 06 CD
 8A C6 70 DE 8A 49 BF E7 47 31 56 1A 4B 55 D8 16
 0D 3A 7D 40 D9 D0 C3 E4 2A 22 D7 EE 2F D2 04 03
 A8 2B B9 0F 26 B2 67 2C 55 28 10 60 01 57 B5 FD
 57 DB 54 B5 86 67 59 76 6A AC 9D C7 B7 51 0E 18
 DB D5 61 0C CA 89 CA E4 79 9C F5 2A FA 80 81 73
 E2 5F DD 3F D1 FD CE 2B 55 D8 1E 23 93 C6 35 AA
 EB 98 0E D8 68 F4 4D F5 8B 41 FC E4 32 55 F6 D5
 7D DC B8 59 B7 B6 43 23 D9 58 50 A3 0E 5D 30 FF
 E4 8C 89 63 09 D4 C1 C6 BC 2A 76 EB 6F 77 86 4D
 91 FA F4 61 43 C7 E2 75 97 10 76 B1 C6 E4 20 10
 69 D4 4F 9F 17 99 EE 06 81 6A 93 87 D0 45 1B 55
 2A 5C 23 22 6A FD B1 68 2F B8 74 EB A4 A9 A0 5D
 8D 18 72 B5 38 ED DB D5 F8 6D 8D AE F3 AB 60 62
 1B 16 0F E7 75 43 98 EE B4 72 46 F1 D3 C3 42 02
 8A B3 DA 81 D6 34 E0 E8 91 90 62 10 06 87 BF 8F
 74 11 11 2D 08 02 46 55 44 F7 A8 0B ED D7 9B EF
 0A CA 88 BA 9A E0 12 4E 92 E2 20 4D AB BC 3F A6
 82 79 65 16 BB 47 41 A6 19 C6 27 C8 93 EC AB DE
 0B 5F 74 67 68 E2 55 14 D8 2A F1 29 C4 98 B9 1B
 07 02 F2 0C D1 48 27 17 01 6D AC E7 B5 BC 0D 16
 31 5B 17 11 3A 39 30 C9 59 A3 EF 4E 7B 1C FB 23
 8B 21 1C 38 7E 3F 7E C1 5F 6E 29 B7 CC 24 55 BA
 2C 54 BC DB C4 FB 6C 06 27 54 99 FF 40 41 46 2D
 32 12 45 58 9E ED E1 86 3D 18 0B 14 44 D8 13 53
 F9 8F 34 CC 7E 45 CE FA 12 AE 7B 60 ED 41 A3 7C
 87 2C 9B F7 61 87 4D 9E A8 01 66 0E EB D4 F4 8B
 25 26 E3 C6 50 BA ED 5F F8 C7 6F 1A A4 A1 91 F1
 40 E4 71 18 33 1D EE 8D 1A 6B E8 4D 7F D3 E8 35
 26 A2 3B DD 10 00 3A 6E CC 05 4F 0C 0B 70 EC DC
 F6 95 88 A3 55 4A 0E FD AC 2D E3 2F 6A 5D B0 6C
 4C 85 0F C6 2A 57 04 20 6D D0 3A 41 F5 22 12 A3
 20 AF CB 25 54 CE CF FB 2A 89 D1 9D 9B B5 07 F0
 F0 02 49 DD 40 FD 11 83 78 74 E3 F4 E7 31 0A C5
 68 8E BF 05 52 7D C7 AB 01 A4 38 D5 B7 63 B3 B9
 01 3C 8A A0 4C 7D E3 B6 26 24 1C A2 A1 38 9A 93
 67 10 59 C9 47 8D 22 08 6B AD 5D 24 6E C9 EA 0E
 2A 2D BE 10 1E DA BF B2 E1 74 66 CD 9E D9 6F 83
 15 8C E1 D9 8D 14 C7 20 9F F4 1D 2A 99 C6 E8 7E
 EB 1B C7 2C 39 F7 A5 1E 96 55 FD 66 24 79 DB 96
 D4 E8 83 8B 1C 19 5E 6D 50 FB B3 96 4B C6 EE 77
 1C DF 15 53 54 19 9C 61 57 69 08 0D FF F3 F4 02
 01 6C 90 60 D7 F3 48 28 6D 19 84 41 FB 7C 61 05
 45 F6 99 96 6D 41 86 08 C2 83 78 7C CB 8A 24 21
 40 A0 C4 68 13 48 F6 22 34 08 50 E5 98 EB 17 15
 7A D9 CC F7 D2 10 04 C8 CE 8B 97 29 26 10 85 11
 0D 0C C1 8D FB 48 60 1B 20 12 54 25 75 F7 70 74
 73 5C 81 6F 87 0E CF 77 CD FB AE AE EF E2 E5 26
 72 69 B9 7A D7 E4 82 E6 B9 41 E4 0E CA 41 3B 37
 10 54 D1 C6 5E 41 A1 73 66 63 0D 4C AF 2D EA 7F
 14 33 79 4D 89 D2 DD D6 70 AC 89 46 BD 4C 22 78
 5D 0F F9 82 25 CC CF 20 DE 20 63 F5 A4 FA 3D A6
 44 1B 45 09 72 91 40 23 1F DD FC 09 25 EC 45 A0
 56 06 62 B4 93 4E A4 DC D0 67 10 31 4C 64 90 5C
 9D FC 19 1B 40 18 D7 EB BE 86 A5 C4 AF 2F 92 CE
 5E 7B 58 9F 11 DF 8D 45 7A 82 66 56 1D E5 29 E6
 D3 86 CE 3A BE 79 3B 33 37 AE 3B E2 2C A6 A6 CC
 F8 AC 69 E8 3F CE BC 85 EF A9 97 A1 25 51 18 F7
 11 36 39 BB 53 2C 74 4E F0 12 17 09 9B 7A E1 23
 36 A7 DD 02 24 34 79 6E BB A7 8A 5C CD 56 A7 A6
 C1 DE B6 54 A5 AA 1D 7E 47 AE FB F3 B4 1D C4 59
 3A 94 16 A3 F3 45 F2 35 BC 1A 6B 5D 2A D1 3D 42
 33 24 B9 5D F8 45 23 96 45 00 40 98 0B 1A 9C 13
 2C A2 B0 62 B1 20 BB C8 C1 40 1D F0 F0 BC CE 0D
 5E 02 77 31 F3 6A 58 F7 62 4F 70 37 18 5D B6 23
 AA DF 86 98 8B AF 39 20 92 18 D4 F3 34 13 CA 44
 A9 30 92 A3 8C 0A 62 3B 2F AA 23 F7 13 51 A6 CC
 05 C7 EA 5D FB DB FC 53 33 BD 14 F0 AE 39 91 E7
 8F 00 2B 52 A9 62 99 67 92 FF 47 B3 76 F7 43 BE
 AD 2A 4B D8 2D C2 05 BF BC 52 D0 75 6A 11 76 1A
 A4 D5 3A F2 4D 76 72 EA 11 74 27 E9 38 18 23 DE
 BF 85 D3 0D 94 80 24 65 BE 60 76 38 C6 54 BE E5
 14 C9 A5 0A 13 B5 F1 8A 0F D7 81 EB BB 1A B4 B0
 5A E9 29 76 05 37 A3 22 48 6E BE A3 B0 BD 54 E3
 D0 D4 70 97 30 92 F7 DA ED 9E 23 D8 67 F0 44 7F
 B7 EA EE 01 5F 31 DC 06 06 E9 BD E5 BE DD F4 7A
 33 C6 DE 14 25 F0 04 DD B7 89 EE 09 62 DF 21 B1
 25 C7 AE C4 33 D9 C9 A8 E0 5B B9 E2 70 4F AE E4
 46 EC 87 BB 02 37 86 A1 11 1D 1A 61 A5 5D 37 2F
 CD FE 21 10 78 E8 1E DC DB EE 9C 50 47 6B 94 7E
 D2 3D 23 BE 39 5F 60 C8 D0 61 B2 9A 41 F9 D8 C3
 69 6C A8 1B A7 A2 64 9A 6F E3 AC F9 5E 4B C8 4F
 1D 99 85 9B 57 E8 E1 B3 47 A7 F5 B4 D8 EC 0D CE
 D1 67 A8 5B 80 0F 7C 7B 43 35 23 71 1D 5A E6 AB
 CA 0C 23 F6 A0 47 A2 EE 82 FB BF 5C 89 4C 56 7C
 F3 C3 40 3C F4 0B E4 EB 24 1C 2C 3B 6F C2 85 87
 16 8C DB 86 AD 8C 9C F3 3F C1 E5 BA E1 37 25 8B
 D1 4A 6A 7E 1A 33 83 CB 60 B7 3A C3 21 77 B9 F6
 32 79 72 28 0D 1E 8E C3 5D 47 24 30 F5 43 B5 8A
 03 AE BA 06 BF 02 6E AB AA 6B 31 C2 C1 84 AB 15
 D0 EB 76 13 42 2B 37 1D 7F D4 6A 3F 9F A4 17 23
 63 22 D2 6F C8 B8 2F B9 C1 87 AE DE 3D 6C 21 00
 1B E6 CF 54 2C 8D 34 D2 E8 22 81 96 1A 5C D1 B5
 3B 2A 32 BA 58 BE 61 62 90 42 D1 63 27 1C 53 08
 9C FC 66 B3 89 5A DA 95 9B 05 A2 AA 22 A4 7A 53
 27 9B 0C 26 C0 35 92 C4 A2 0E 11 D5 4B 7D 20 0C
 85 86 BE 85 66 1A 71 DD AC A6 52 BC 26 C1 CC B8
 38 A0 B7 B5 2A 11 55 F6 1F F0 98 8E 32 F2 5C 9D
 BF 67 8F 19 83 9E 3B 69 EB C4 B5 43 C6 AF 39 89
 A8 30 B9 9D 99 33 6A BE AF 6F 96 A1 5E CC 86 1C
 E2 34 09 96 FA 49 39 D9 F0 73 79 99 7E AE 35 61
 1D 9C 18 15 13 80 C7 92 76 0E 86 19 17 BE FB 2D
 51 DB AD 4A 6C 3B BC 83 54 FA 05 28 65 1E A8 3B
 70 89 3C FE 58 87 C2 34 8B 89 06 4A D1 B1 F3 47
 2A C5 33 A2 7A A5 5C 46 5B 4D 0C A2 1C 7F 1E EB
 06 9D CE 3C 97 92 70 32 BC DD 4B C6 9E 72 17 8B
 29 31 53 07 1E 9B F4 33 05 AC E6 B9 13 71 0A 54
 0A 26 ED 71 D4 6F 78 51 02 FA 4E 29 7A 7E 2F 47
 6B 2B B0 24 D9 32 EE B1 90 05 3A 49 E6 6F 21 C3
 F1 DF 1C 70 DE 8C A0 9F DA 69 5A 07 9C A8 FC A7
 AE 89 FA 22 E9 53 4F 43 34 5A 32 1E DE 22 13 0A
 DB 9B 62 F9 82 F5 E5 8D 73 DF BB A7 97 1B 2A 50
 B1 A1 BC 40 F0 CD 5E 25 46 AD CD 54 D7 BC 3E AF
 AB 35 A1 27 8B AA 63 A2 06 3B C7 72 5B FF 38 A1
 B2 93 5E 85 2E 6D 52 BC B1 F1 28 5B 87 5F CA F9
 06 4E E1 9E 26 4A FA 25 13 17 37 23 A9 85 BE 36
 5F 9C 55 D6 B8 19 C6 5D 60 14 BF 50 DE A1 41 1A
 11 5A 03 E6 6A A7 DC B5 32 71 E9 F2 0E 09 CD 87
 44 3C E1 B9 0D 05 73 4E 69 47 99 A9 F4 17 C1 F9
 2F E5 85 16 63 5A CE 04 26 C9 05 4D B7 A1 7A 6E
 64 68 5A 93 E2 99 E9 3B 95 9C 78 02 FC D5 A4 A8
 1D 55 29 F7 14 33 B0 D9 98 15 46 C7 78 C9 6B 52
 67 DF 2C 5B 8B 49 9B 12 69 94 D9 38 D9 D5 20 F9
 F0 28 85 D8 18 81 96 57 C5 4E 9C E1 B6 B9 9A 3C
 5E 73 32 7E 20 25 BC 82 97 AB 12 14 78 56 7F DD
 4D 95 36 4A 13 14 FD 13 66 55 FA 5D 4E E7 AF B9
 41 76 F0 BA AB AE 84 7F 90 EE 39 36 5E 86 1C E7
 66 BC B1 52 BF 54 45 EE F2 ED 26 BA 14 10 7F 5D
 78 51 82 DD B9 37 E3 69 31 93 2E CB DF 58 64 23
 3D C7 B1 CB E9 A3 F6 D3 B2 F4 44 4B 5A 48 B0 22
 B7 C5 47 CD 4E 0D 4E 35 CE 7B 96 E7 E1 1C 5E D6
 EB F7 00 65 17 0F D9 37 00 10 EA 0E 44 5C 84 9A
 57 DE E8 FA 13 0A 87 D8 93 12 5B 34 EF 4A 58 1E
 E6 DD B8 80 BB C3 3A 4B 9E 7E D6 38 0B E4 96 06
 40 3D 11 10 24 BE 32 A4 9A 01 6E 34 64 96 62 5E
 FC BE 54 13 84 1A 55 78 2F F5 BD 1B 99 41 8A BD
 61 9F 0C 20 CB 25 3A 12 1E C7 3E 0B FE 60 03 3D
 65 64 CD 5A 59 79 F6 65 D3 FA A0 00 AF 87 CA 66
 9F 42 6A 06 65 B7 D9 5E C0 BC 6D 00 98 97 6F 4A
 F7 85 00 0E 8F D8 52 FE C7 1C 40 8E 77 03 02 22
 E0 36 5E AA 05 C7 B6 16 1E 6B 69 54 17 13 D8 93
 1D 06 80 44 E8 C6 76 9B 68 13 C3 DF 7F F4 EA 18
 89 50 F9 A2 94 89 16 54 CB C2 50 1D B9 24 73 3D
 B0 36 D3 1B 76 49 36 F5 E1 0D D3 5A DB E4 70 51
 9F E3 D9 A0 16 32 91 4C 31 9E 0B 48 84 1A D8 7A
 B8 E3 7A 22 E6 43 81 1C AB A3 60 BD C2 23 A5 53
 31 C0 70 C2 81 91 37 24 95 C4 14 CA 3D ED 46 95
 DF B1 6E BD 79 9E 75 6F DD C7 42 BF 8F 64 A6 B2
 8D 21 31 92 3E E0 65 01 2B 53 85 EF EF 35 16 0A
 C5 FD 82 4A 3B 45 FC 0F D7 04 4E BC D1 57 73 E0
 B2 ED 5A B8 1E 41 45 56 8B D6 27 BD 7F A6 07 C4
 FE F6 8D 46 DE 9D E2 04 69 A1 04 85 30 91 B4 E4
 2B F5 93 FD D5 2B B0 B2 0E 62 84 EE DA 30 FA 07
 4A 7F 9F 1D 0F 22 11 5E 51 2C 7D 27 2B EA F9 EE
 0B 62 EC B6 AF 5D 7C DE EB 68 5F 2A A3 9F 65 21
 75 0D 57 C4 36 47 9C 40 9D A2 FF AB CD FB C4 93
 75 B9 50 2B D4 51 9D 25 57 05 86 5D AA 86 36 49
 D5 7B 61 57 68 B3 4A AD DD 71 1F B5 6D 43 9D D1
 E6 0B 31 8B 90 78 55 7F 8C 5E 49 CA CA A1 47 9B
 85 8A B0 DE 25 E6 B9 70 0B B4 63 78 B6 08 F3 B5
 A8 66 90 47 E3 93 EF 30 21 E0 D2 BF A8 9F 1F 89
 6D 22 DC 44 42 DA 16 A3 03 79 20 8F AB 69 40 02
 5E 4E BB 6B 62 9E 49 36 2D CD 4C 88 DC 36 41 D7
 8C 51 1D B5 94 FA 12 3B A7 7E 31 42 8B D8 9A 0A
 CF FE DB 30 D0 2B 6C 5E 33 74 95 14 18 21 C9 D5
 68 7F CF 17 43 AF F2 0C F2 EC 8F C0 E6 64 61 D3
 09 87 57 F1 E5 BF EA C5 7E EA 34 2B 29 D7 7C 0A
 92 44 5F E4 C6 82 E7 A8 B6 AC 64 13 A4 03 A1 EF
 7A 55 B2 3A 77 11 04 27 81 36 98 CE 2D CE CA 94
 81 A5 F6 19 86 A9 C3 0C B1 3B FC 52 86 22 14 ED
 53 9F 1D 64 BC F0 8C D0 F6 F2 DC 79 9A A1 DC 38
 26 E8 88 B3 94 A0 1C 0F 9B 6A 6C 8F F0 95 0E 8C
 58 A4 DC 21 6A 8A 0D 17 33 AE A2 1B 7C 68 05 BD
 CE 05 DD 7C D4 62 B8 32 94 3C 4F 3C CF 08 5C 9F
 8A E4 3B 2A B2 AF F1 34 16 1A E7 64 F4 E8 55 F9
 46 13 21 37 4B EB F3 68 2D 70 A1 E7 F2 9C E4 CA
 2A 7F 06 F0 41 95 12 16 8D EF C5 93 4E C1 EC 10
 B6 87 AA 28 4F 93 71 4B 33 A4 68 46 DE C6 D0 E1
 83 29 38 CA 40 86 4A F8 86 D4 08 64 71 23 9B 1F
 EC F3 29 76 1F 4F 8C D1 F5 3F 53 43 61 00 AB 44
 93 BE 77 7D 99 F9 DC B7 18 7E 9F D2 BF 84 2B A6
 B3 9E 2D AA 1A 6A A1 C8 87 52 D6 CE 36 82 07 B4
 99 AE FF BD DF AB CB FC E9 1A EF 77 9D CD 45 B3
 52 07 78 76 22 94 5D B8 D3 72 65 77 2F 02 C3 18
 14 F6 9E 15 1B 10 D1 B6 E8 20 34 9F 1C 62 1E 8E
 52 53 97 35 34 AA 8D C4 BE 0B 04 F1 AD AB 48 6E
 ED FA 71 89 E7 3D 94 8C 7E 14 A4 84 DE A5 9A 0E
 A7 6C 12 19 67 A8 FA 55 BB C9 BE 0D 5D AC 0E 94
 A6 25 7B 8C BE 90 C5 AF 30 E1 17 F2 CF 61 A2 69
 F6 7B 0F FE 70 C2 BC D4 0F 85 90 C2 69 9B 44 31
 D6 D0 36 99 FF B7 E4 98 1A 9F BF 91 51 B1 8C E7
 EF 73 22 DC 21 FB A5 DB 30 F3 98 A4 C9 13 5B 0E
 C0 3A A7 6A 4B 3E 0C FA D6 80 01 30 D6 EE DE 75
 D6 61 22 0D 8D BC 09 CD CD FC 43 48 56 78 E8 4B
 B5 23 0F 76 C9 3B A3 BA C6 8D F3 76 63 D3 C6 41
 1D 8D 60 B4 0B 2A 0C EC AF 29 AC 94 6F 23 5B E4
 7F 72 6D 61 F9 E2 94 C8 56 AF C5 5C AC D4 A6 B9
 82 4F 94 00 EB 3A 31 7C C5 9E 65 EA 45 77 5D 35
 25 90 27 EF 73 BC 86 4E 39 85 92 5A 13 77 EF 29
 FD DF BF CD 3B 5B CE 60 BE DE 45 F3 16 40 76 D5
 96 F6 EE A7 36 EA F2 89 5C 00 33 35 76 79 36 7C
 48 8A 8C B4 77 BB 88 F8 EB A9 B4 26 F3 1D FD E1
 05 5E 79 24 4E 2D 04 E4 3D 8F DD 4A 65 FB 1F 54
 A8 7E EC F5 91 6A 53 C4 82 0D 62 28 56 F5 51 4E
 B7 C7 91 08 92 05 6C B7 4E 26 4D AD 10 09 08 BD
 34 9A 64 BE 30 C7 23 09 54 73 04 2B 88 22 81 98
 6E 13 8A C0 2C 14 E6 A2 5F C6 C1 6B 7B 21 11 F2
 B3 3A 32 29 F3 90 F2 19 A0 77 7D A3 37 B1 F6 B5
 4C A3 11 3D 07 6C 28 39 C3 4D 0A AB EA E1 B0 C3
 3C 60 7A 6A F7 3A 26 7E 78 34 6E 4B CA 82 4D F8
 B5 39 8B C6 AA FB 39 C6 6D F8 E6 63 3B 03 93 7F
 B4 42 A8 AA 4D 21 3D AD 3B 11 43 91 9E 30 F2 0C
 72 FB 87 A6 D5 FB 5A C4 2F 43 10 B7 92 5B F5 54
 BC 44 69 D2 3A 74 23 EF 0E B9 34 FF AF BB F6 F5
 9E 4B 0C 7F 31 52 B2 95 83 AC 0D A0 61 F1 B1 24
 38 8B 78 A9 B3 EA 98 0D D2 68 BE 4F EA 31 29 E8
 EF DF 5D 0E 31 B2 BE F9 8C E5 5C 1D 17 C4 D0 AA
 6A 1B E1 B2 1F 25 25 6B E3 1E B5 F8 15 E0 38 BC
 4A DE 1F B1 F0 74 04 58 0F A4 58 1F A0 F3 28 21
 28 24 42 E0 F2 83 AA 97 55 F8 F4 19 C8 E8 D1 01
 E8 65 AC BF 9E 00 0B 3A 98 50 78 D8 FA D8 0E BF
 7A 06 80 62 8A D9 86 48 80 D0 17 C1 99 1C 8F 02
 83 2C 52 20 03 A9 91 06 4B 4A 14 87 D3 E4 8D 45
 6F E3 B1 67 72 9E 0A 57 56 28 E1 15 75 BF 58 EB
 36 ED A9 2C 9B 4A 8A B3 20 9E D1 E1 6C DC 50 71
 0F 20 B6 E0 A0 06 72 26 B4 CF 30 40 D8 8C 34 37
 D7 29 9B 48 FD AC 9A B2 6A A9 30 6A C1 ED CB F8
 1F 78 AF D9 C0 19 DF A9 DE AC B9 BF 39 D3 03 15
 0A 14 F3 BF B3 78 13 BF 4D C0 45 3A A8 93 EA 9E
 10 32 BB 95 23 33 58 AC 62 2C C1 8B 2F 13 5C 0C
 20 26 23 B3 84 D9 23 09 C2 6B 47 43 72 13 F6 49
 D5 25 E1 B0 BE BF 8D 70 5C 2F E3 7F 10 8C 7B 5C
 48 D9 BF 2F B3 D9 BC B4 D5 3C ED 92 BD C6 38 C3
 75 D1 1C DC 42 50 98 61 6E C2 A1 6C 8E 18 21 1C
 9E 2D BF 4C F7 70 EF F7 EE 1E E1 2F 8F 14 60 C7
 95 00 B0 B9 60 0C 73 85 76 AB 4B C4 E0 EE 14 11
 5D 88 DE 9E 59 48 61 D0 1F 1E E5 2B 16 E4 53 2A
 BD 9A 47 BC F6 73 96 60 22 42 72 79 2D 00 D2 78
 B8 D5 55 C5 3B 1F B0 EC 77 2C A9 7E AE 2D 2F 68
 16 C5 2D BE AE 5C DB A3 6F 38 04 9C 7E 99 64 DC
 F5 8F CA 6B 18 98 85 39 27 FA D2 10 EA 78 02 F7
 9F 4D 0F F9 B7 F7 77 62 E2 C8 CE 13 AD 4B 11 07
 4B F9 8B 4B CF 8A EE 68 C5 0A B3 A4 28 45 80 BB
 41 DA 69 B9 F7 E5 E4 0D 3A 81 3E 45 AF 5F FC C0
 E0 D8 31 FF CF 57 1C E0 B9 5D F4 16 3B 14 4D F2
 AB D8 4B 34 4E 93 24 24 37 3A 8B CF 5F 37 2C 25
 CE 4F F9 8B BF 83 18 0A 6E 6A D7 A7 30 8B E3 9E
 76 6C 12 8B 28 48 E5 D8 B8 D9 32 E5 4C 85 AF B6
 91 DB B3 07 4D 08 74 A1 4E D2 CD EF 1F DA 1B BF
 4D EE A0 6A 2C 33 A2 D6 E2 76 38 97 5F AE 65 EB
 05 A0 3C 93 36 74 15 AF 00 07 50 B5 7D 54 C4 1C
 7A AB FE 2E 22 B7 82 93 76 2A 42 46 D8 EF 30 72
 D2 E9 76 90 48 24 3D FF B8 50 EE 29 75 39 7F 01
 E2 E7 13 2A D9 04 03 CD A4 16 09 C5 94 04 48 D0
 3F 09 C7 73 07 8D 21 3C 66 BD 04 EB 89 30 D6 60
 8B 49 C2 47 FD 75 29 83 7F BE 81 EF 73 45 20 A8
 04 34 13 80 35 EC EC C0 95 E3 65 C5 A6 B9 B2 EB
 41 B4 26 18 B0 D7 F8 BA 32 A8 F1 70 38 8F 3D AA
 1E EE 97 FD 28 56 5E 79 26 58 71 03 F4 FE 2A 3C
 7D C6 F2 0F 87 2B 32 77 51 C8 04 6F DF FD 21 7D
 FB 89 40 F8 F4 47 68 4A F7 59 1F 6F 03 A3 87 85
 73 88 FD BD EE 68 D7 CE 31 76 A9 CD 46 22 23 F1
 A6 95 EE 26 E9 E2 36 C2 AD 72 94 98 EF A7 74 C7
 A1 A2 75 94 1A 8E FB 96 AE 11 87 F4 95 47 5F A4
 E0 52 03 6A 09 B1 D7 C0 22 2C A4 7B 7F E9 24 CC
 39 50 19 72 A2 DA 88 98 F7 63 86 E1 BE 2C DC 7E
 C8 94 C3 E6 60 80 97 0A C9 32 66 C4 D1 E0 67 58
 50 E8 4D B9 CE A8 0F 34 73 8F 04 09 C5 38 8A EA
 85 A4 42 EE 66 F0 E5 FF 86 35 B5 86 F3 FF 5D 8C
 D3 87 E4 C2 1E 21 66 1D 9C 96 AA EA FF C0 B4 9E
 7B 6E 87 67 6C FB 2B BB 2F 1E 65 B5 4E 50 FE 04
 9F 75 DA 25 A6 49 10 70 84 2A A5 E4 3C 0F C0 70
 9D 14 AD 50 77 7C BA 08 DF 23 40 B8 4A 3D 7D 11
 F5 21 6C 59 5B 7D 80 BD 92 F0 10 C4 14 A9 49 60
 B1 09 E2 6F D4 49 F3 82 05 CC 16 58 F9 61 AB 22
 BB 4A 8E 01 DF 04 E3 41 64 04 E7 9D A0 B7 8B 2F
 69 26 77 E1 10 85 E1 E3 11 F9 EE 2D 97 65 29 26
 55 2E AF F4 D1 F5 26 20 57 96 1D 9F 73 21 DD A0
 28 FF 67 D1 FA 68 20 EC 57 AF 20 1A C5 59 3B 99
 69 EC 96 C7 3E 3C 43 1B 01 88 C5 89 B6 E3 C4 E6
 9C B0 85 88 72 06 51 6F A4 EB 5C 0A 73 70 FD 88
 39 94 74 3B D4 14 5E D1 99 8E D7 E3 21 E4 C1 C8
 BD D7 CC CA 11 2D 1C 29 3F B8 B8 3C D5 6C 0B 6B
 5D 94 5A 38 2A BD DD 3F 4B 2B 81 AF 06 29 9B 89
 69 5B D8 B3 2B EA 14 FC 65 C7 BD D9 01 20 62 A6
 8E 19 CB 4E 82 87 69 DC FB 7A B8 43 80 74 FF AB
 6A B0 4D 84 3F 53 1A 9B A5 71 B3 2B A2 06 F8 5C
 7A BB B0 E2 46 EB 32 7C DE 3E AE 00 A6 0D 6C 44
 DF 30 6C 2F 87 9A 5D AA 1A CC CA ED FB B0 C9 A5
 4D 9E 2D 04 A9 94 2E 3F B9 E8 4D 7D AE 46 55 B9
 94 C9 10 CB 21 3C B1 7C 57 C7 7C DB 3A 0E 24 1D
 C5 6E CC A7 4F 09 EA 10 FF 3E 42 78 AF 73 F9 2C
 74 AB 47 CC 86 04 A7 F2 23 99 63 CB 2C 9D AF 61
 AC EC 18 5E C5 52 57 0A F1 9C 37 B3 7F 3C 70 49
 4A 5B 2A 53 B7 0F B5 73 B8 23 BA C8 FD 22 0A F6
 0D AB A0 A8 02 36 72 4B 84 E5 3D F0 84 BA 02 BF
 18 E2 42 76 F8 70 3B C3 AB D1 B1 8A 8D 8C 02 AE
 0B E4 38 E4 51 11 AC 27 C6 17 48 28 0F 41 C3 FD
 4A 3A 81 69 76 63 28 AB FE FA CF B6 B7 D2 40 F0
 F3 8A 01 79 A0 AB 0C 58 B9 6A 15 93 D9 0A 88 15
 76 78 DF A7 A6 D5 85 01 36 DC D2 43 69 44 2E 25
 1A 5B 45 D6 B8 12 40 4E EA 47 F0 A5 C6 91 94 EA
 1A 45 5C C0 F9 3A C3 61 C7 34 72 5A FC 3E 71 11
 EF 2E A4 3F 10 AA EF EB 09 F1 73 19 F0 72 A3 E5
 4C D1 04 4F 3D 65 3A 3B 81 55 E8 1C A3 B7 00 31
 54 8D D6 F1 30 E4 B3 F9 3E A4 94 09 FB DE 8A 01
 35 41 2D 3A B2 C4 B0 46 1F BD 70 78 FB 44 1E 7F
 90 99 A0 1B 8E 13 93 9C 92 F8 D6 B0 14 EB BA A7
 97 76 E3 2A 6C 2F D4 47 F5 5A 35 F3 C3 39 18 F3
 CF 44 1F 1D FA 5C 51 6A EE 3B ED 8E 61 92 A6 BA
 23 4E FD 80 57 AD 9C D3 C2 B0 BC 55 F3 26 C8 6F
 8E C1 56 DF 49 D3 37 03 4D E2 9A 4C 4F 43 73 04
 8C F1 60 4A 78 26 D3 FA 69 87 CA 0F 3B 00 DB AE
 23 D0 7F 30 4A D4 FA 91 2D B2 FA C3 07 8E 67 67
 25 F6 2C C9 11 BF 6D B5 AE 73 95 C7 85 00 DD 62
 36 C9 2F 13 D3 A1 3F 5D CA 3C 25 BD E6 C2 0C 4C
 F5 3C 9F 44 DF 42 24 85 E1 80 3E 48 15 05 56 56
 64 B8 44 04 4C 45 06 C5 6F 4F 9F 4B 6C 3E F1 D5
 98 01 D2 BC 26 EC 66 DC 92 C4 20 51 05 CC F4 93
 DC 2C E9 A3 C0 26 F5 21 90 18 5E C4 94 7F 36 50
 A7 15 99 8D 94 DE 68 F7 1D 23 66 4D 30 EB F4 FB
 9D DB 53 FA E7 28 F6 48 A7 5C BE 14 82 56 ED 93
 75 E1 EF FE 19 46 B2 7D 74 6E A7 93 80 B2 26 68
 E4 47 B2 70 E4 ED E6 9F AA 4D 9A 5E 76 BE 52 16
 36 C3 47 B8 12 BD 2D 01 A6 91 E4 A2 4A 4F 46 D6
 DB B8 62 BB 03 9F 9E 72 27 CB F7 48 77 C1 0C ED
 58 EE B9 FC D2 E1 A4 F0 F0 64 1A 09 39 A3 8A 75
 17 96 04 8E 6A 73 28 78 41 2F D4 C2 22 2A CE B1
 E7 80 C5 C9 77 F2 11 4E 01 C1 DB B1 45 AE BF 1A
 25 72 8B 2C A8 4A 35 66 CE 38 6E 0F 59 BD AE B8
 DE C3 90 90 9B C0 9D D2 CF EE CE 44 F5 31 B8 40
 EF A4 8C 6B 01 1F D9 32 FC C7 60 5F 28 23 E0 2B
 C3 23 FA 9D 0C 86 BD 56 89 74 6C B3 37 68 54 84
 D8 5A 66 EC 3C 34 A7 BA A4 4B B4 5D B9 29 3B 83
 97 2D 44 86 60 C0 0E 90 75 F0 80 99 DD 77 D1 2F
 B1 C1 A6 1E 1C CA B0 6B DF 40 EA 89 81 88 2E 51
 0D E0 ED 04 D0 A7 CA 57 A3 56 BC 96 0F F7 1A 31
 02 16 FC 6D E9 75 B8 CC 8F F0 08 B8 15 45 58 BA
 EB BE E5 06 A3 C0 84 AE 65 59 87 D3 8E A4 C5 8E
 9F 58 29 E3 F6 25 8C 6D 08 24 E3 D7 33 C9 6F 65
 BB 13 B0 DF 3B 54 39 8F 7A 33 6D 70 1B 8E 2E ED
 7F 7E 05 60 8A 35 D4 03 32 50 14 35 71 26 D9 A9
 0F BE A4 A0 A5 74 16 B5 BF 7C C7 37 64 FC D7 29
 3A 2C 5A 55 42 9F 77 C6 E8 62 66 72 B8 38 9C 85
 2A F5 FA 23 DA 48 6E 5E 79 0C 2E C3 A6 CA 29 A9
 A5 1F 57 BE 99 1A 5D 14 38 54 6B 3D EE F1 0C 53
 B3 62 5F 87 07 5E C1 EF A4 00 2D 5E 1A 24 A5 7D
 3A 94 71 37 AC 54 03 FD 59 43 82 A3 F7 67 1E 9B
 66 F0 BD F0 BE CF 42 11 3C 7E 75 F6 14 CF 80 CB
 B6 4E 35 11 6F 12 80 7E 6B 02 2E DB EF 44 8D 63
 F9 B1 AC 0C 43 CF 17 D7 08 BF 19 C1 E3 9C 84 E1
 50 5B A1 3C 6A FB 85 E0 AE 14 CE F0 F3 90 FB 1B
 91 8C DB F5 C6 DB A9 2D 37 20 B0 1C B6 28 5F AD
 BF 1E CF 34 69 7A D0 A1 30 70 1A 7A A1 77 05 F5
 28 67 0B C6 11 2D D6 11 CB 1A 67 2F 71 07 8F 95
 39 05 77 73 27 5D 6C 19 DA 3F 41 2E EF 68 9C A8
 6A 36 06 43 95 A6 73 30 40 40 4E 23 28 AF 91 96
 6B 1F 77 79 3D 95 2D 20 CA 5D 81 24 E9 A2 6C F5
 91 9C D0 48 4A 4E 06 61 81 12 01 22 C7 56 82 FF
 EA A5 3A 86 07 BD 03 30 CA CD A5 A2 6A D8 DD 05
 64 EF 77 BB 12 C2 36 74 14 28 38 ED 82 52 41 70
 B3 74 A4 86 A8 5E E7 79 D2 98 EE F6 85 32 1F 4B
 60 E8 34 BE C5 39 8A B3 24 7C 39 1C 8B BD 3E DB
 D5 AF BE F8 87 9B 6B 54 C4 8A 7B 67 5E 8C C0 02
 A9 8B 66 6C 48 34 DC D4 57 99 5B DA CE BD 17 A0
 FA 95 F7 A4 E8 67 3B EC 14 95 5D 0C F2 DD 22 D5
 20 EF 08 92 AE BD E5 C0 C4 D2 BC 52 FC C9 C0 DA
 E2 52 AF 1E 13 4D 89 7D 57 3E 56 56 70 C0 BE 1B
 D2 79 0F C0 A0 91 B6 48 D1 BD CA F9 BB 92 EE 56
 7E 7E F4 AA 95 97 E6 AB BD BE 3C 38 D9 99 CF 20
 0B 68 30 38 F6 10 45 D6 F1 B9 E9 2F EF 6B 6B 92
 FB 6F 86 41 C9 C0 EB F8 EC B3 D7 75 4A 39 53 F5
 C7 6D 37 39 90 B4 D9 80 A6 A3 2D D2 33 3B B1 AE
 EC CF 3C EF C5 18 37 39 CA 41 48 8A A2 C6 2E 9A
 69 CF 0E 14 D6 8B 4B BA 90 0D BC FB 6E 11 82 73
 6A 72 5C 49 5E 6C 0A 4D 37 47 56 C1 41 3F F1 7E
 A6 63 ED CA D2 47 23 96 43 81 2A CE 32 79 C8 7F
 FB 15 38 FC 8E EE B0 C0 55 18 A3 AF C4 91 14 80
 7B A6 33 8E D7 D9 45 20 29 BA 7D 28 0D E0 11 7F
 90 B0 8C EF 82 30 9D 98 BE B3 03 8D CC A3 1C B9
 99 AF B1 EE 4C 50 5D B1 76 45 0D A6 48 8F 23 74
 F5 4D 63 45 6C C2 55 50 A2 A4 FF 85 5F 04 43 E0
 AF 55 43 87 15 88 88 84 95 3C B0 36 4D F3 C1 D4
 E6 B3 43 DD AB 7B 3D C5 3A D0 78 F0 E9 1B B0 55
 2E 74 F9 52 B6 C6 04 20 A9 1D B3 96 C9 AB 81 5C
 CF 4F 21 4A FE 00 FA 41 99 03 EF E9 54 0D 2C 07
 FF 0E 1C 2B D7 D0 D2 C6 51 FF 36 B1 08 5E 88 BE
 A4 F1 83 4B FB 1D A3 75 E2 59 76 9F 78 1F 84 EA
 45 AA 35 2F BC E8 F3 6F A6 A4 8F 19 A3 0A 32 5F
 22 0B 2E 11 42 B6 44 A4 F5 96 1D 6D 89 89 0F 90
 9E FA 3B 08 E8 7B 93 6F 7F 6E 0F 99 59 45 DD AE
 B7 AF A2 F2 45 3C E2 0C 2E 82 77 FD D5 33 EB 75
 47 D2 52 92 3E 76 6B E3 D0 2F 3A B8 2A 60 31 8F
 E4 32 2F C1 B5 64 04 4A 3C 64 61 61 96 75 BA EC
 FF DD 77 75 7F 61 D5 66 F6 A4 5C 71 DF 23 74 DC
 23 F9 8B A5 D1 0D B3 F4 69 10 83 1B 36 16 DA 62
 E4 66 C5 0F 26 1E 8F 64 CC 11 F1 EF 1E 13 75 99
 0F 6A 67 F6 40 B6 9F 7A 7B 77 89 02 22 4C 02 91
 B2 72 AE DA B3 03 48 5B 89 B8 1C 7F 15 C1 E1 75
 CD EB CD D5 F4 1B AC EB 8D FF 7D 5C 75 39 18 0C
 75 45 82 46 83 20 F3 16 27 3F DF 27 F7 C9 3A F2
 C7 EF DD 19 7F F8 D9 42 0D 32 0C 57 4A 18 3E C8
 44 4B B4 24 A5 29 82 6E 0D 3E 65 8E B8 F3 B5 DA
 17 26 DC F3 7C 9B 9F F7 15 E7 D9 FF AA 53 FD 33
 97 B6 16 90 DE E7 E3 B9 BB 9A 3C 5F EF FE 68 9C
 EB 5C CC 31 32 5F 2F 62 45 9A 41 9D 21 BC 63 DB
 83 76 84 FE 74 B7 06 43 99 A1 16 FA FE CA A4 25
 06 B8 6C 2C 67 AF D1 70 32 D1 71 26 D1 8F A7 99
 27 07 BF 42 9A 7A 5F 17 27 73 BA F7 A5 A2 CB 0E
 1E E0 B8 4A 0B 05 65 E1 3E B4 D2 92 7C 39 20 07
 AB E7 DC 81 66 31 B5 E2 C4 8A C0 0C 24 56 D4 19
 AD 0F AB 9C 90 14 4F 42 B6 41 E5 47 70 7E 51 A5
 AC C5 25 CB DC 75 F7 13 EA 6B 73 65 2E 5C 46 9B
 30 88 2C E4 78 7C 9B 76 53 95 7E 16 9D 1A 95 94
 90 41 C2 59 40 EF 9A 34 45 5C 1B 7B 86 6F B2 4D
 F1 9C B7 81 64 6D 90 98 42 23 56 A9 5C 32 10 82
 1E 5F 67 BF 00 72 7D 08 ED 65 B8 D8 8D CB A0 BF
 5F F8 32 9B 84 F3 94 27 4D 9F 23 FC ED ED 35 A2
 BA 2B 85 CD 47 B7 C5 A3 97 20 08 3F 5C D7 EE A6
 CE 6F 9D 77 EC 8F DA FB B7 BE 79 52 A7 69 9E 36
 EF EC 87 B3 B2 83 57 7E 52 F9 99 44 86 39 D2 1D
 AE 2B 0D 0A 4D 0E 72 4C 3A 44 58 9A 34 E0 0E 9C
 84 0D 9D 16 AA 95 EB 4F 3F C3 79 19 F4 D9 7D D7
 97 03 57 70 9A 1A E7 14 E6 B4 E4 63 0C E6 94 93
 89 3B EF 2E F9 F1 06 40 2F 79 CA 4A F7 3A B8 C9
 10 87 2B 2D DE 4D 19 D9 81 AF F3 7B D8 FE 3B 8C
 0C 1A 48 A0 4B 56 6F BA 56 67 3E BB 77 17 16 8E
 CC 09 9D 3E 61 82 F1 E8 6A D1 EA 98 29 80 A2 7B
 BD 16 D4 0F 54 73 4A 80 BB 57 71 A9 CC 8B EC D5
 0A D0 41 09 32 1E D2 6F 14 28 B6 07 16 DF 49 18
 7D 7B 41 ED 84 95 5D 84 57 69 15 F4 0C 53 E9 7E
 F7 A5 45 78 29 2B B6 ED 89 D6 D2 A3 15 5C 8B 86
 59 A4 F0 65 AC B3 04 E4 C7 28 F1 A8 27 2D 2E 10
 AA 7A 32 D8 93 F5 13 C4 80 7B 2A AE 75 66 AC 8D
 BB BB 4D AA 98 CD B3 B4 A0 E7 F7 5A D7 97 31 F0
 8E AB B3 7D 71 A7 D5 C6 9B 10 98 B8 F9 67 73 77
 FD A5 F4 61 D9 03 55 7B 5F 0E AE 83 EC 73 13 D0
 9D BA F8 B9 D9 87 DA 9C 82 3E E9 5F 73 4D 6F E1
 AC 99 D2 55 9C AB 1C E4 9B EC 21 A9 E7 75 CF 22
 E8 A4 BD F5 C5 68 15 BA F5 B9 02 A9 8B ED DC 33
 FE 05 85 7A ED 86 6F 89 E7 09 15 94 41 0F C0 6E
 F7 A3 F2 A4 AF 4A 49 9E D5 05 1C 5E BB CE 19 CE
 8D 19 84 9D 30 BE 25 3C 52 3F 10 A6 3A 04 84 19
 B6 48 99 CE DC B6 7D CE 60 DD 2C AB E0 12 DE 34
 48 B2 96 3F C2 7C B2 5D C4 CA 3A 14 A1 E5 6E DF
 78 B0 2B 5B 91 AD E2 56 DE 76 CE 46 4C F6 21 67
 9E CD BB 8F D0 C2 3E 71 F1 11 AC F8 77 F4 A8 8E
 3C EC A6 FC 7C 1B 37 55 84 8A BC CE C8 3D 87 FA
 9B 34 AC 3F F1 D3 E1 1E 66 92 C3 AC 44 54 20 CC
 87 A5 F9 2A 6A 5D 54 8D 28 30 F0 57 18 14 50 6B
 2C 76 5B 33 4F 4A F6 23 FE F1 CC 5E E5 B8 01 21
 1F 23 11 8A 79 5E D5 C6 D2 88 4F 5A B5 43 7A 5D
 47 43 85 8D B6 7A 7C 04 A7 BB BF 3A 48 14 CC 2D
 E4 B2 DE EB 03 F7 80 97 73 3F 6F 5E 90 3E 61 1A
 F7 98 CF 31 B6 BB 10 DB 62 CC 23 20 76 62 68 1D
 9E 82 A8 88 A4 04 87 ED 46 1C 53 68 88 A7 4E DF
 29 AC CD 3A D0 6D 4D 3D 7A D9 9D 79 02 BB EA B4
 20 F9 F4 F9 B9 E1 29 3B 9A 6F 61 53 C8 2A E1 AC
 C6 6E DD 1D FC D2 EB 51 08 2A 02 62 74 2F 15 7C
 41 B4 A9 12 E4 F5 A6 5D 95 70 2B DB 14 0E 7F EC
 1F E5 86 55 46 91 D8 C9 BF F5 E6 EF C1 3D 97 D2
 2A 2B D6 19 6D 64 7C EA FB 97 9D 70 E3 AA 3B D7
 4B B2 E5 04 76 32 E3 C7 D6 F0 13 C4 C0 8C 80 D8
 BB BF 30 C5 27 4B BE 6F 21 B7 91 B8 26 77 C3 6E
 67 D8 02 40 16 D1 36 14 8F 7B 24 60 16 6E 1D A1
 C6 C8 17 DD CD 63 75 0B 8A DF EA 0D 18 DB 02 0D
 DF 7D 64 B8 8E 75 10 D4 B2 19 E1 7D DA 45 F0 6B
 6D 81 24 C2 74 8C 13 09 7F C4 B0 0D 8D 0D E5 C7
 A9 66 9A 01 7D 8B 4A CC 17 2E 35 5F 3E A3 4E 60
 D9 BE E2 9A CA 77 62 DC 7B 6B 18 A6 82 CC 82 C8
 C8 F6 28 AD 7E 3B 4A F4 83 89 99 0D 17 34 41 F9
 0B 13 E2 99 FE 8C C6 66 B9 52 65 FB 9F 60 E2 98
 12 91 AD CF 00 62 31 DD 84 D8 2D AE AA 23 3F 6C
 CD FA FB D9 83 69 1B C7 C6 45 EC 2C D0 27 68 9F
 62 17 7B 89 EE 9A A2 72 19 12 25 B8 72 8B D7 A0
 11 BF 7F DF F4 17 D4 03 66 58 D6 0D C7 20 6B 03
 B5 6D AB E1 D6 25 0B 11 FB 2D F0 F6 38 A7 10 1B
 09 F3 80 29 B2 FF D0 48 CA 48 43 92 6E 8B F0 83
 5D C5 5F CB A5 E8 40 A7 04 C6 63 63 1C 9C 7D 0E
 22 DA 2F 0D 17 D6 23 76 7C 5F 8B 01 A3 6C 33 02
 76 27 84 C4 13 A5 B9 E3 1E 69 96 BE 37 A8 52 57
 CF F4 39 E8 36 DE CD 76 11 B6 74 64 9E 62 17 DB
 3F 87 CC DA ED 03 4B 6C 3B 99 7C 66 82 47 DF 87
 9F F1 0B A0 21 8A F4 9A AE 46 2F 76 CF 34 44 77
 70 0F 7F 44 99 D6 F5 0F B2 7F BC AC 33 50 64 56
 A7 6C 29 A6 35 1B DE 2C 65 5F 69 6C 74 8F D3 A3
 62 95 AC 87 42 BD 3E 05 1F 91 6E 0F 2B 74 D2 46
 42 E8 D5 5A 64 31 D9 14 D4 E2 29 89 54 4C 55 F4
 71 6F 92 0C 36 9F BC 24 31 20 6C AD F3 B5 06 5B
 6E 23 25 B6 FD 04 D6 44 8F 16 34 A1 35 A6 19 D4
 3A 72 76 91 82 94 6D 6D DA 4D E4 80 AC AC 94 89
 C0 7B 42 F4 5D 48 55 47 5C 23 73 BA E8 86 CE 5B
 84 85 75 C0 FD 1F BD 20 1D 52 EA 27 12 E6 7D EB
 D0 92 1B B1 88 F5 3D 9E D7 7B 0E 96 E3 6A 43 98
 FB 47 C4 BC 10 7A 44 F2 B7 E2 FA 57 BF 5E 42 34
 6B 26 EF 2C 7E C4 5B 3D 1A 14 9A 21 0C B8 92 84
 5F C6 FF E4 4F 53 7C E0 C7 45 29 7B 07 16 95 67
 F3 E2 C0 07 96 A4 2F E4 C1 58 53 3E D9 B1 12 FA
 92 7D DA 87 93 ED 5A D3 0B 88 53 8F 60 D5 9E 10
 65 CF D1 46 16 F9 DC 39 3B FE 40 39 9D 65 60 A5
 C1 8A 30 4C E1 7B EC 08 E0 68 FD DC 99 FF B5 BD
 FA 2E AC DE 53 29 0C 8D D6 91 AE 07 FB BA 3B E0
 BF FC 2C 04 E1 44 25 8F 1F 5F F6 A3 77 9F 5E 0F
 CE 42 7D 69 09 65 B9 2D 03 55 A6 D9 20 CD 25 29
 CA 92 03 E9 72 7E 53 0F BA 25 79 50 64 96 74 F8
 88 26 DB 40 4F 04 33 0D 49 EC 95 41 A2 CF 6D 1D
 9E CB 66 8B F5 E3 9E 45 B1 48 F9 5E F5 DB 47 B7
 F5 1F 3C 17 A1 08 E8 E8 ED B5 89 F2 4E A2 75 DC
 79 4B D7 A1 F1 EB DB E4 E6 03 A4 39 4C E6 67 75
 A5 47 2E 39 98 C5 B5 65 B8 B8 85 10 B4 97 D5 51
 13 A3 75 0F 07 4D 93 B0 19 08 E0 77 F2 97 BD C0
 0F 26 87 C1 62 4F 5D 94 45 8A 86 29 FB 22 2D 12
 08 2A 9B AA E5 FA 1C 1E 38 FF EE D2 2B BE 22 2F
 CA C3 FC 35 9B 13 E1 DC DB 3D 1F E0 29 16 96 FD
 B9 7F 24 5B FC 17 0F 6C 1F 88 94 DA EF 8D 44 72
 08 83 FA A9 F2 43 C5 8B 4E 5D 92 76 0D 81 4E 0E
 12 A7 1A BD 93 BB A1 AA AC 44 77 64 E4 F4 E2 9B
 58 3A C0 CB 94 10 ED 13 27 32 28 9A DC BA D0 73
 4E 29 38 09 95 1B 5E 15 D4 25 E8 EE 50 E0 39 CC
 7F 88 C7 2D 3A 34 62 FE 85 E8 78 85 63 0F 74 11
 CB 3A E4 A7 0E 7C 4B 9B 53 10 D2 27 35 37 E6 CD
 E8 6D 68 DA AC 68 56 8C 04 B9 89 69 C4 90 9A EE
 18 4A FF 16 B2 0E 2C F1 BB 8F 8E E3 39 13 82 1B
 2D F6 0B 89 C6 46 6B AE 11 4C 65 FB 40 1C E3 80
 A3 18 1A 8B 7D 6E 85 77 3D 7D D0 ED 58 19 23 F2
 FF 5F 09 89 16 A6 B7 89 76 22 B7 92 D3 88 66 1F
 EE 4C 33 3D 5E 51 B9 A5 AE F1 21 89 AA 27 BE 80
 8B 63 02 96 00 94 5D 9E ED 19 E6 06 DF C2 05 56
 95 0F 5D 54 E8 0C 7C F7 0C A5 AE 17 7D 36 A7 FE
 B0 92 A9 4B CB 43 A9 F3 3B 2C 6D 3C BF 64 AD 62
 FC F6 8F AF E4 31 96 79 2D 4D C6 3B 66 DF 8D 06
 8F D5 A0 74 DD 53 B0 43 47 61 3C 9F 60 03 C9 34
 71 34 C7 EC 6A BE E0 39 3A 4E 78 66 8E 9A 75 4C
 D8 B4 B9 DB 14 4C 4D B1 3B F7 40 47 3B F9 06 55
 99 E3 A0 5E 33 64 1F 86 A1 9D A7 18 7C 99 C5 B7
 FF 8C 76 DC 1D DE 7D D3 54 86 D1 1D 61 21 4C 60
 85 33 A8 10 01 C4 3E FF EF 91 9E EE 9F 0A 35 1F
 1B 55 40 37 F2 C9 8B 94 BD B6 69 D1 6D 94 EE 57
 DC E8 C4 8B D2 9E 5F 2A 45 6A 26 3A EB A3 F3 2F
 27 5C C6 38 4B 04 93 60 86 72 FB 0E 7C 46 98 6A
 87 3F E4 DC CB 94 93 94 09 17 6A 8F 53 58 77 3B
 09 89 EA D0 93 28 78 C5 6C A7 48 CB CE 2A CB 84
 34 3D BF 87 0C AB E8 A1 02 FC E1 37 D8 8D F6 A9
 CA 0D 7E 8C 9A 90 27 DF 2C D0 0C 37 5C C9 D7 DB
 E1 DF A8 2D 97 9B AE E7 18 B4 2F 15 29 FD EF A0
 68 00 A7 C8 B1 DB A2 0E 9C B2 C0 B5 F8 90 DA 75
 A4 41 71 11 89 79 C7 18 B9 B8 9E 47 EE A9 5A 7B
 59 D4 06 55 19 F4 49 FD 3F DD E6 E0 FD CA 40 1E
 DC 56 68 0A D5 C5 BA 41 F0 73 FE 39 D0 08 5A 07
 85 3C C6 A0 F0 B8 19 17 AB 9C 41 20 59 AE A9 0D
 34 5B 90 01 02 DD 26 63 87 7F DD 44 14 2E DD 86
 36 60 AF 9D A1 3D AE 97 7D 26 76 49 E9 39 20 F5
 DA AF 2D 52 29 41 CE D2 C4 62 31 60 E4 74 2F F1
 B5 F4 4F 44 C4 0A 98 74 D2 5E 6B 01 12 A8 17 9B
 0A 84 54 7A 3F 44 09 80 38 9A A3 68 C7 10 4D 33
 53 8E 04 12 EA C2 B2 2C DD 5D C1 72 EF 5B 52 D9
 B3 A5 BC EC 5C 44 BD 5F 22 DD 8B 0E 5A 7A C8 82
 CA 9B E3 74 9C 9B 41 F6 42 B3 AC 8E 68 68 38 7B
 7E 93 22 AC 18 B9 19 78 F8 EC 82 6B 30 87 07 94
 67 3B 10 E1 25 59 13 00 04 80 A3 8B C1 AB 83 73
 67 C5 9F E8 2F A5 1B 68 21 64 35 11 85 84 B7 0D
 AB 53 0F CA FB D1 E6 F3 F1 FC E7 91 6B 73 C0 6D
 8E 79 A4 8E 95 1E BC FD 33 D6 52 53 D5 D0 7D 72
 C6 A6 F4 58 90 0B 22 3F 24 E4 7B 07 E5 8C 43 36
 F2 70 F9 BF 01 5F 76 09 B3 A3 E1 BA 90 E5 67 7D
 D8 0E FC 67 64 BB 21 68 10 55 11 01 40 27 D2 97
 35 97 CA 7B 1B FC 38 A5 8B 28 64 5D C2 6E 98 93
 D9 46 1E C8 49 47 0A B0 41 59 F8 13 1C ED 8D AC
 10 A6 F4 C8 B3 09 5D 0C 69 C8 B2 43 AB 2A C4 AA
 09 62 3A 96 F5 EC 1F 9A BD E9 2A 15 3C 3A 95 7A
 CA 38 6B 32 C6 74 C1 E0 5A 68 F9 74 02 F3 E6 67
 B3 5D 67 F2 5A CD 5A 1E DA 39 61 6C B7 49 07 D4
 5E 45 F1 47 72 BA A1 79 69 3B 8B 43 3D 05 23 9A
 ED A4 1D 1F 3E 55 D1 C0 51 23 BC FB 70 39 86 44
 8A B1 56 58 D8 85 4B 0C 41 35 1C 65 34 27 C6 41
 43 E2 92 FB 49 83 01 C3 E7 FB B1 56 44 18 32 C3
 17 27 5B 22 B6 30 C9 9D CC 0F 05 C8 9C 86 66 1D
 C6 27 F5 5A 5F 75 3B 5C 01 AF 9D DE 33 7B 84 BE
 BD 15 B1 D4 FF C7 09 1C 71 E2 61 4C 04 44 3B A0
 29 D8 99 8C D7 6E 43 5F F5 B6 D5 7F 96 79 52 29
 44 00 51 E8 03 96 D8 CE C0 CC 6B 4A DD 49 7A 5F
 CD 88 58 E6 CB 94 BB 8B AD 41 BD 57 B7 CE D3 73
 47 03 73 0C B2 CA A9 09 84 38 DC F9 14 0E 72 CA
 03 B3 27 E2 97 F3 F7 BE 52 0B F6 4A 01 1E 8E D7
 F2 7D A2 5C AE 41 90 D2 65 E7 E9 FA 39 E6 5F B7
 02 C4 85 11 D1 C8 BC D8 D2 44 93 06 D9 42 61 7E
 1F 55 1C 93 A3 4B DD F2 C5 C9 87 DB 16 A6 E8 3C
 C4 DB F7 06 AA 8E CE 06 16 0D 1A C7 C6 5F A4 01
 12 5D FA 96 98 9D 8E 58 C5 41 82 5B AB A7 D5 CA
 25 EB 6D 38 AF AC 8B 0A 67 E1 E3 52 4C D5 AC 84
 96 A9 EE BF 0A 13 1A 31 4B 77 0F 34 87 40 C7 C8
 CB 75 6F EF D9 33 A8 B3 15 3F AE D6 1A 72 24 E6
 2A 32 2B 8B E1 5C 31 3B 50 65 13 6A 31 EA D5 AC
 CA 5C 0C 4D C6 CC 9E 5D FB 57 1D C3 75 2A 0D 59
 61 7A 99 4C EA 74 54 99 C8 75 85 69 C5 FB E3 94
 CA 00 B6 71 B1 01 E9 FA 42 43 AE 5C C1 01 A8 0A
 CF 7E AF 6F D8 60 30 9E F7 A3 62 C7 F4 58 5C F5
 CF CF D5 BD B0 58 AF 95 06 AF F8 7C 5B CD 6A 38
 EE F0 26 6D CE 43 E7 54 BA EC EC 17 97 8D 3B CA
 86 0C 18 BC EE FD AE 31 AB 38 D1 53 32 CF D0 41
 4B 93 73 63 F5 97 9E 3C 0A EC 98 54 F7 04 6A 3E
 DF 6C D1 7E E9 11 43 4D A2 92 ED 9A EB E2 4E 8A
 3A 82 9F F9 3E 4C 73 08 63 A9 E6 75 7B 4E 5C E8
 18 ED 69 86 6F 57 E2 2E D5 7D F3 AE D0 91 38 DE
 09 74 81 B6 72 16 04 EF D6 3D 80 36 65 7D F0 B9
 41 F9 DA AA B4 D0 0A DE 0D 3F 50 12 B3 B4 DF B9
 38 58 AE 2F 61 37 8E AE 2D 13 76 10 90 38 12 4B
 AA A9 BC 4F 74 CD 45 52 B8 A3 EE E9 66 44 C9 8C
 66 B8 0D B0 E2 39 4E 58 54 28 6E B9 5D 1A 68 2B
 31 2D E2 FA 8B 84 28 40 EB 85 0E B2 50 2A 83 BA
 61 B1 C6 04 D4 DB BC 63 78 14 88 0B EE B4 A6 B8
 57 D7 80 A9 5E 1A 0E 70 48 21 79 53 BF AF 42 D2
 65 9F AD 1E 92 2E EB 19 4F 50 4F 2A 23 0B D9 4C
 C5 84 D4 68 E9 35 74 8D 78 11 0C BA EC 8D 57 58
 A7 1E 4B 51 DB A6 7F 75 9D A9 AE 89 ED CF E5 A1
 BE D1 B5 43 B6 E7 CD 9E 2E 62 F4 48 15 4F A6 7C
 14 3B DF C0 8F A8 17 8E 9B 3F E5 50 AE 4A 66 3F
 62 90 AC 42 DF 68 5A 44 48 60 22 10 2C CD 39 C6
 71 22 B6 5E 99 4C 79 F1 79 08 3D A8 0F A5 D5 B0
 3F 34 60 1E 83 EE E2 21 C0 38 CE 34 57 E6 B9 3A
 4D 10 97 F8 0D 22 70 DE F2 F8 7E 75 ED DF 0B 06
 8E C5 7D 3B 2A AA 01 AC 4D 59 E7 88 ED 21 AD 7D
 28 BC 67 83 B8 70 D2 BA 6D 84 CB C3 38 76 64 FC
 89 61 AB B5 A1 D7 88 20 18 E6 31 29 D4 5C 20 55
 29 25 CE 93 27 C6 A2 AF C3 4F 08 10 A2 6F 5B 6A
 05 03 AA 47 05 E8 C0 68 72 D5 E9 56 2A 65 A3 00
 96 E8 E5 B4 DB AF 7B 71 8F E4 0E 2E 2A 3B DC B0
 A4 07 23 35 65 C8 93 02 E6 38 AA 95 24 BC 95 BC
 77 EB F0 D6 77 9B 71 B9 55 02 A9 F2 94 59 A6 44
 59 69 4F 76 2A A8 64 5C 25 E0 70 D1 80 23 9D C0
 85 39 5C E8 25 F9 2B 09 21 DF 43 CE D6 CF E1 C6
 4E 64 0A 46 EF BB 65 F9 33 48 AE 58 5E AF AF CE
 0F 7D E6 DF 7B E3 AF 63 58 C5 C3 C2 29 AC B6 14
 BD 2A 63 54 9D 20 15 32 EC F5 93 A5 B8 9D F2 38
 4F 40 01 FF AC FD C6 43 79 B1 33 DF 3D 48 3E AE
 0E 9A 85 C3 57 DD D1 05 67 92 6A 2A B6 4A 1C 1E
 8B 77 B3 35 63 E3 C4 49 95 B8 7F D8 D3 0F 9D 70
 46 4E 81 34 69 CC 36 E0 B6 6D 78 D7 6E 5D A2 0B
 47 F9 C2 60 10 C7 B8 AE 2B 7A 3D 60 4D FB 16 52
 E6 59 56 63 76 E4 82 EA F8 B9 42 ED 35 E8 CB 69
 51 2C FF 2C 27 30 E9 8C 17 1A 41 DA 03 EA F1 E1
 2A D6 ED 5C 40 2B 34 AC 83 CA 92 EE C0 6A CE 15
 49 3C 6A BA 6E E4 E0 2C DD 36 10 DB 00 80 3A D6
 03 2F E7 C7 0B E0 24 D4 14 1E 81 34 AA 64 BD AA
 83 27 A7 26 8B 77 C9 62 8A 33 42 5B B2 D9 92 62
 D8 C1 4B DC 7A 58 BD E8 18 7B 5E 33 40 71 CC 20
 09 FC 98 57 60 F7 98 6D 49 30 25 43 4B 97 EA 54
 F1 EF EB 71 E2 34 1A 11 FA 48 91 92 90 CF 32 3D
 BA 04 48 91 71 7D 11 FA EC 6F C7 CB 9C 14 B0 E4
 48 51 C0 D7 DB 1E 56 0B F6 E9 C1 BA 1B F2 F0 4E
 25 40 37 AB 97 F3 63 BE ED E7 A3 77 DE D1 C5 88
 C6 56 DA 15 A4 40 18 5B 76 7C 5C 5F 47 94 B8 01
 75 AB 79 16 41 7F 21 BF 6A B4 5D 55 E2 0B 75 00
 42 F0 73 EA FB 0F FC 84 19 4B 50 7D 28 40 36 F6
 47 8F B1 64 4C CD 18 73 5D F9 AA 89 9A A1 25 F4
 CF 2D 8B FF EA 12 64 21 33 C0 B3 A2 B6 DE 93 0B
 D6 CF 8A 1C 42 51 EC EE 3C 32 B9 8A DF D1 3A 4F
 50 90 2C 17 5E A4 00 FD F0 E4 17 2A E4 33 F1 15
 8C B4 74 F3 88 9B 70 C6 23 03 66 B4 4D 63 93 E0
 F4 7E 70 36 7C 12 F4 8E E5 C1 FD A0 F6 94 0E 6E
 E8 77 69 98 7D C3 7B 0C D0 3B 70 7A 28 BC D6 CD
 3A 34 80 82 D8 76 65 34 F0 45 9E 7A F9 15 2C 2E
 4F 0A BA 9C 2C 93 82 A9 F0 63 E8 E7 BA 3D F1 6B
 CC F1 A6 81 B0 C5 A0 9E 4B E3 64 BD 23 2C 1A C3
 35 C9 26 8D FB 31 F9 13 B4 DF 50 D1 AD B3 A5 E5
 2F 8B 7B 82 96 49 CD 20 F6 1A 3B 95 2F 78 EE 4A
 0D 36 26 8B D8 D8 6C 8E 0B 29 1D 54 92 B3 C8 2D
 B8 1D 77 C8 6E 0D 34 29 29 E8 AC B7 AF CF FC 4F
 D5 94 65 DA CC 02 2E E8 88 58 18 D8 D7 E6 BD 82
 2D C6 E1 01 61 AD 6F 0F 19 9B 9F E5 21 A3 35 44
 D0 1D B0 ED E3 56 F7 EF 68 DB 9C CD 99 5E 83 88
 A3 FB C6 96 71 F5 24 6F 6B BC 17 36 C8 84 C3 0C
 96 11 E7 40 C3 F8 35 F6 37 58 1D 03 C9 94 C5 CE
 C1 55 2C 33 C2 4E 36 BD 2C 23 CA F5 DF E1 65 1E
 D5 21 5D 61 7A 0C 10 4B 4C 03 13 A3 79 E8 45 F1
 05 CA EA AB AB BF B6 C0 47 C7 D9 F8 6D 0E 19 BD
 4D 6B 97 F9 94 7B 34 F1 B5 48 A3 6A 31 FA 62 3E
 04 44 57 98 50 6F A9 AB 56 20 3D 99 A4 41 E0 A1
 A2 EB 56 28 CC F9 97 AD 76 0C 9F 52 B1 B7 98 43
 64 66 AA 61 1A EC 69 6C 09 C6 E1 39 5F 35 A1 2C
 82 88 1B 72 F1 0D 00 00 B9 91 21 41 2D BF A1 05
 2B A9 5B 67 C0 CF A2 36 52 93 91 22 88 8B 55 43
 B7 95 88 92 CC 43 BC EE B6 9B 6D 4C D3 49 CD 67
 62 C9 50 1B CB AA 40 A4 A1 45 C6 FE 99 0D 21 83
 88 7C BC 6E 7F 6D 13 EE EB 5D 03 D2 E3 4B BB E4
 18 55 B3 E7 60 44 69 4E AA AE 84 DF 2C CD 83 97
 82 BC DA AD 08 33 01 2A FC E5 BB 53 51 04 C5 24
 D6 B8 AC B8 BD 65 D8 55 A0 8A 61 0E 08 D7 FD E0
 2C EB 9A 69 A3 F8 1F 38 85 07 92 3E 2B 4D 44 81
 10 8E 43 E1 AC AF CE B6 21 D2 3A BA 59 FE 92 52
 ED 31 C6 4C 65 33 BC 84 2E 0E F8 06 86 75 0C 83
 EB 04 6D 5F 33 A8 13 82 B7 CF C6 E8 23 FA 9F 07
 8B 42 18 0D EF 93 39 17 86 FB A1 EF C2 2C F9 8E
 95 0B FE 40 53 55 D7 01 54 41 77 1C 43 43 08 BD
 98 D2 4A 40 38 BA 47 01 D0 AD CE BF 18 47 BD 37
 77 C1 B8 2E BC E8 35 CA AD 93 DD 0C 28 2E 2F 6E
 9F E8 B8 59 08 0A 46 94 A6 F5 74 20 20 A5 A0 C0
 77 96 38 3E 65 FC 9A 1B 06 7B 45 F3 FA F0 D6 89
 5C BE FE BE A2 27 65 F2 8C CE AF 62 F9 37 A4 40
 01 5B EA 34 A6 2D 38 13 53 68 A5 A7 F0 B4 C2 8F
 DF AD AA BC 48 6E E5 09 7F 91 8B 19 C3 86 16 B3
 F8 DF AE 81 A9 A2 75 8A 61 1F DF 74 AB F2 D8 7B
 91 02 66 37 B3 A4 B3 BC 5E E7 A5 09 91 BF 04 8C
 D7 54 42 84 D2 E8 5D 36 DB 58 B8 40 20 42 CE 09
 E4 94 36 A2 D0 C8 5A F0 5D 91 1F F8 D5 15 F0 75
 01 AC 49 74 18 75 C6 69 39 C2 EB C7 57 9F F1 69
 E6 95 05 DE B8 17 A9 58 81 5E 0F 7D C3 0C DC 75
 12 CE 50 F4 71 B1 0A 9A 08 6F C0 C7 46 99 B0 72
 CF AA E9 2D 9B ED 6F 5C 05 81 0B 84 7B 87 33 A8
 C9 4C 97 64 DB 6B A2 4E FC 99 25 9E 55 77 2C 20
 97 61 29 A0 49 35 BE A8 E6 D2 CD AA A1 9B 3D 8E
 D5 02 32 AF 8A E8 7E 22 42 DB AB B7 D1 98 F0 07
 66 53 37 14 A5 56 67 F8 6C E9 0A 68 2F A1 E4 7B
 0A 01 B7 2A C2 33 78 8F EF 11 6B E4 AD D0 51 A6
 53 8B BC C9 4E 10 11 21 2E A2 78 A2 AE 8B 97 48
 47 49 C8 48 8B 16 17 F8 18 B2 D5 8F 87 80 13 08
 CC 15 CB EF DA D3 92 50 EE 20 2E 9D 4C C3 06 76
 78 70 65 0D 8F B4 7B C4 DA D1 89 51 E9 2A 25 E1
 9D AE A6 A3 F0 07 49 25 E1 F7 F9 79 1A F7 00 D8
 50 E4 D1 DF 07 17 8E 43 1D 5C 5D 4C 0A CD 96 B0
 22 1A F3 96 84 87 AA 74 E8 0A F5 F0 79 D0 96 31
 2D 44 D7 85 4A 49 CE 53 1A F2 32 C8 79 1C 98 EF
 0D 46 CE 0A 5A 57 A4 51 07 10 28 DA C0 D6 21 BC
 74 70 46 69 A2 DF CF F9 1E 0F 9C 68 05 DA 4E 7E
 F0 D7 32 1F 11 CD 00 2E FF 6C 86 81 9C 68 23 A5
 D1 93 44 2E 3F AD 45 3D 14 DB AC 39 5E 7F 5E 77
 0D E4 77 5D 7E BE 0D 10 66 09 18 6A 22 6E E4 05
 00 A3 69 0A 1D EC 64 BB F9 C1 34 55 9F F6 D7 6D
 85 95 47 80 31 0C 21 6B 3F E1 AC CD 1B C6 E6 A7
 06 0B C5 CA 44 6E 35 CE AF B0 91 17 6D AC 9C 07
 47 87 A7 D1 49 A2 79 D5 7C 61 7F D6 92 3B EF 6B
 17 AA 80 B4 FD 8A 44 E6 FB 72 2D 1A 58 CC FB 0C
 A9 A8 AD 4C 7B 17 80 48 34 2C BC 5D 03 E0 53 95
 20 7E 98 CE 1F 10 18 37 BD C2 CF 73 76 F6 D6 7A
 19 C7 F0 D4 F9 87 05 7C 89 E9 34 D7 00 1C 49 82
 F9 71 F5 43 1A 10 88 84 DC DA E5 9F FB 9E 9E 18
 DF 62 EB D6 34 D4 7E 55 54 30 69 4A 6E 2C F0 24
 FC 28 04 0E 73 B4 1D 60 5A BB 37 A5 16 F8 63 FF
 5D 6E 3E 2B 10 7B 81 2B 61 53 BD 01 46 BE 85 4E
 73 35 AC C4 28 A7 70 06 3D 69 F7 26 3A 11 30 D3
 2D 06 6C DE 2E B8 67 E7 35 F0 22 94 A8 51 EA AA
 E5 39 99 88 8F 8E 41 77 EA 5B 68 EA 00 C0 B2 CB
 02 10 61 34 F7 10 5B CE B0 06 2A 86 82 61 A2 AE
 80 0B C6 A3 D7 F6 C3 DD 1A 8D 07 24 55 38 D9 6E
 7F FC 80 AD B2 0C 94 DE 13 F9 CC 31 B1 40 27 7E
 F9 3B 33 C5 23 73 79 DE 80 84 ED 8D EA 60 F0 0A
 8C 04 60 80 40 29 B4 81 4D 22 88 22 95 1D 24 65
 51 F4 14 13 EC 84 96 9C 16 D5 CB 9A C6 16 CE 58
 03 D8 1E CC 02 8E 7C 3A D2 68 A4 92 05 C0 41 6D
 AC B5 3C 27 2F 1D B9 DF D0 AC 47 E5 CF 7D FF 06
 0F E1 4A 15 A1 43 14 64 F9 F2 D5 01 4A 8D 69 63
 DB 5E E6 A5 EA FC DC 62 9D C2 60 AC 42 AC DE 33
 03 8E 22 6C 48 28 83 B8 D7 E8 D2 9F 5C 59 4D AE
 08 0C 33 D3 BA FF C3 08 B1 02 FD 71 A4 55 FB D7
 F7 5A B3 3E 8F 87 10 5E F2 4E 84 B6 F4 52 B9 6C
 98 41 8B 44 5D 8A A4 B7 21 67 CC 8B C4 8B 53 CB
 6F A1 CE E6 C7 57 5C 42 BB 12 DA FF 56 0C 55 9C
 3B B4 CB 93 A1 5C 34 A2 BA 2F 72 F4 F3 FD 3F 49
 2D E6 C6 40 4D A8 31 1E C2 32 28 50 80 9D F6 87
 AA 0B 4E 7B 4D 99 F9 A1 BE 72 EC 47 66 7B B0 34
 56 13 C9 35 8A 0C 52 13 5C 3F 7A 88 FA 58 AD BA
 33 37 9D 90 7D 30 D2 8E FF 92 3F FB A0 ED CA CA
 64 99 BA ED FC F9 07 37 68 7E 06 12 A1 FE B7 D3
 9F A1 3A 3A 94 3E 61 EC 36 5E C1 62 28 19 BD 69
 EA 41 4A E7 29 44 AC B6 23 E5 6E DD 15 F9 87 91
 9E 83 1B B0 F9 21 D7 75 31 F9 BB DC 72 43 94 B4
 B2 64 49 8F 4B 59 33 6B 58 7C 10 1F 98 84 B1 0B
 8A 13 A0 CC 87 EF 42 3D 48 14 DA 27 60 53 0A DC
 19 4F 3D D0 7F 52 52 E0 97 A3 BA 09 A4 8B 58 48
 7C E2 1C 88 B9 83 8D 7B C3 C0 A8 3F D8 61 81 82
 B4 C5 33 15 E1 C4 81 FF 8A 06 AD 03 8D 76 C6 45
 65 7D DB 10 9B D7 B7 17 20 FE AA E2 83 6B CF 9F
 D7 93 0D 26 87 56 25 87 51 A4 C5 A4 BF 87 15 D2
 F5 CA 8B 7D 5F 03 0B 81 61 30 84 41 F7 0F 78 2F
 96 71 B5 C5 94 A4 FC 4C 35 05 C0 1E C2 34 FA 7B
 98 4C C0 5D 90 E3 E6 7F A9 35 FA 51 9C 23 C1 33
 4D 77 28 82 60 AD 6D 4D 80 15 29 B9 7B 83 65 8A
 8C DB E6 B7 77 07 13 72 97 23 B7 54 D2 33 A6 6F
 69 D5 25 CB 97 A6 85 0F 44 35 C9 DA DA 51 E7 4B
 4C 79 B3 59 B3 AA BD 36 9F 9B A8 32 E3 95 68 AD
 04 4C D9 B8 FB C9 14 CD B9 A1 D0 DA 21 3E 18 D1
 66 EF 4C 3C 8A 78 2B 22 D4 2F FB 9D 3C CB 8A 8D
 3B 24 8C 85 E8 41 20 61 7B 3F 89 26 D6 71 A7 42
 60 3D EB 2F C0 48 6B 69 80 DE 68 51 D6 09 A6 31
 1F 92 9E 7F 3B AC 8C 95 0A 78 F2 ED F4 BA D8 A0
 C4 B9 87 91 B9 55 89 5F 1E C5 77 DA 46 07 43 82
 54 13 F1 35 97 14 86 8D 58 52 31 64 00 1F 83 06
 4E A2 E5 8D 7E 85 0D 95 5F 35 79 60 5B 0D 42 A1
 25 B2 61 A0 7E 2F 3C 31 8D 71 6E B0 59 8D 67 2C
 36 58 70 70 80 94 93 56 81 BA 59 B0 01 9C 6F 20
 33 AD 7A BF 2B 39 9B 08 D0 DE 75 F5 89 25 C8 3A
 C0 64 DE CE E6 0C E5 4C C6 04 68 F1 B3 FD 77 71
 BE 96 5C 37 75 E8 7A 69 A2 63 98 02 96 72 CB F0
 79 CD 2B 33 32 C9 0E AB 64 3F 2C DC 4A 67 77 00
 C2 D3 69 70 B1 48 3F 68 60 F2 D8 8B E4 E2 00 59
 A0 86 86 88 55 DE 44 75 46 7E F7 C6 E6 B2 92 A8
 AE FC CA 82 F6 1E C8 51 79 E1 CB A1 4F 25 D7 BA
 42 FB 28 55 A7 95 C7 B3 47 23 8F 26 2A 20 9D 68
 F6 B8 81 F8 F8 08 3F 91 9C B7 67 0F 36 3F 3D 5E
 A1 1E 10 23 AB C2 B2 95 33 C0 84 96 DD 9F 5D 71
 C7 36 B6 3F DE 79 B4 09 FA 0A EC 37 1C 32 09 3C
 5F 18 56 6F 5D 03 F5 D6 4D 53 A7 FD A3 6B EE 9D
 60 AA A0 FA 6F FF 92 41 2A 97 A5 50 4B DF FC 1C
 14 F4 B3 21 3C 4E 00 E9 B4 98 C5 F5 D5 E0 0B AC
 71 53 0F A7 AE 60 E9 36 6D 9F 79 25 B9 0C 81 DE
 2A 6A C5 D8 E0 61 95 AF 0A 46 D2 DF 20 2F 29 A0
 98 DD 2C 8F 9F FF 9E 38 14 BF 91 CC 7E 0C 3C 55
 6C D3 0E EB C4 37 7D 8B 91 FE 94 18 FB 11 F8 88
 18 4E 75 0F F7 1A F3 22 42 18 3B 31 E8 A0 93 3F
 FD 07 DB 9F 4C F1 FC D1 A1 32 D5 94 B2 B8 DF 4B
 70 32 E2 0C F6 A2 36 63 A2 B7 61 9F 2A A2 2B 86
 E3 77 8B 10 6A 33 93 B5 BD 7F 55 7C A3 95 A3 A9
 59 B2 70 C4 17 52 23 25 E6 94 46 A4 F8 F3 A2 AF
 C0 5A 83 4B 06 BA 8D 62 F4 E7 F5 70 6F 59 B9 7C
 E6 C7 83 B7 40 D5 B9 AB DA 7C A2 1F C6 DE 7C F2
 4B 9A 69 CC DD 78 35 C4 C2 E6 56 CA 60 3D B0 1B
 5D 2B 6B 9D 8C BE 09 2D 27 7B 3E 59 D1 67 5F 3F
 26 BB A6 A2 5C 56 53 8E 97 D9 3E 30 AC D3 D0 D7
 DB AF CF A9 20 4A 62 9B 95 B8 32 94 E5 F8 AB 5B
 5C F6 54 2D 93 1B 9E EE E6 13 A9 6A 26 90 A1 A2
 F7 C5 58 CF 8D 19 7E DD 0B A3 93 0C 39 4C 60 DC
 00 B6 19 D5 4E A2 F3 34 F6 9E DE 3B 0F 86 3B 28
 CB E5 E5 1B 42 BF 10 7A 39 1C 02 25 A1 EA 00 8F
 57 57 6F 59 6D F6 02 38 C3 FE AB C6 27 12 62 DC
 A0 C7 79 29 38 29 56 9B 0B 04 28 33 2D 2D 2E B3
 28 04 88 C1 E6 97 FC 22 94 2C 07 D5 7D 97 13 AF
 63 05 C8 0E 18 6B 57 27 B2 1B 9B 28 7B 1D FB 1E
 FF CD CD 71 39 CA 9C 8B CB FF 2D 16 BB 07 6B 14
 EE 31 77 EE E8 C5 4B E7 DE AA 23 F0 03 74 9C 7E
 84 D5 9D DE 90 AA 7D 8C 63 3F 7A 55 31 EA F1 D1
 14 70 23 E9 D8 82 09 57 FD 55 CF D2 E7 DC 16 DA
 1A 8D 5C 5C B0 0A 7A 82 FD E3 18 BF 63 EE 5F 4B
 53 A5 87 90 F9 1B 87 CD AA CF A8 9D D6 73 34 A1
 78 3A AA 7A 24 81 8F D5 40 2B 4B 45 9E 64 CE 5D
 A7 66 18 8A BA A4 6E 06 7B EE F0 70 94 CA 2D 19
 04 72 D2 22 7D D4 AA CD 18 8D 0C E4 14 02 13 BB
 C8 93 4F 71 57 65 CA 97 21 86 EC F5 C7 0D E8 8E
 F0 D1 3D 42 D8 FE BD F0 12 E7 AC 5A 9E 13 B6 92
 B7 A8 C7 CE 74 69 12 D3 AA 2E F7 A1 DD 6E 28 89
 15 61 AB 91 CB 4B D3 44 3E FA 7D DC 2E 5E 6E 71
 E0 81 65 46 DF 01 C3 8A 2F 1E 4F 65 46 DD 11 20
 E7 41 45 93 4E 48 C9 E9 2E B2 48 88 C2 AD 0F A8
 61 61 5A 49 57 61 23 0C DD E6 CC DA FA 09 76 53
 91 75 EA 1D 7B 89 B7 FA E0 C2 70 7E 21 4E 51 C1
 D4 ED 14 13 8E 85 0E 97 C5 B2 27 BF 61 6D 26 94
 65 47 59 C4 35 80 B3 4F D1 4B CD A2 1A 8C 88 29
 56 25 35 2A B8 A1 1D 55 51 61 ED 4C 58 3D CC 9F
 FE 34 F3 B2 9A 81 0B ED B5 86 F9 F5 E2 C2 4E A8
 D1 17 46 2F 7A C8 12 FD 3E D5 AE 3E 80 18 82 26
 F3 7D 8F 59 42 0A 6B 58 B4 36 F6 AA 10 27 E4 56
 92 AC 80 9B 32 AC 2D A3 04 FD 8B 61 D7 BD 7B 59
 54 2F FD 66 8C FD C2 FB 2D CC 1A AD 29 6D 0E 5E
 71 F3 1F 93 6F 04 1F 72 88 60 A7 C8 2E C6 BF E8
 0A F7 2B 5A 8D 61 A5 AE 21 62 D6 B8 49 A7 6E E0
 B7 37 C8 0A BE 69 D9 CF E1 05 C6 56 4E C2 91 F3
 5F D7 E5 4B 02 A6 65 17 14 8D BE 48 FB DF 68 E9
 7B EC 28 66 F1 75 27 51 CB DA BB DF D6 3B 85 A3
 14 4B FD 90 46 70 ED BA 0D 90 30 77 D4 8E BA A7
 F0 D3 5F 05 42 9C 9F 58 87 2B 7B 7A 96 6D EC BC
 61 26 40 51 A8 7B 77 81 D4 42 5F 74 DB 0B 0C 40
 22 60 96 78 D4 55 83 50 2D 77 DD 69 41 56 D0 5E
 84 3F 6E C2 82 1F B8 C5 06 4C 98 19 91 7E 98 9D
 DF 3B 97 BE 18 2A A4 89 3A 3A 78 DF D7 15 A6 C2
 02 9B 87 D9 79 8D CF 34 9A 31 79 32 D9 16 18 67
 E6 77 67 AA 23 79 D3 7B 06 6E 16 49 23 05 D6 97
 AB B4 87 38 22 B7 D1 E9 C3 9B C6 E7 C4 6B 96 0B
 37 6A 65 E0 86 67 13 91 26 63 ED 85 14 CD CB 9C
 D0 D2 8C 8E 36 A4 91 B7 F9 E2 04 AD 08 25 59 20
 70 AD 08 79 8D 54 56 BE 9E 1C D1 10 C0 7B 3F 14
 0C A3 D9 1D 07 08 D2 54 BA C3 74 25 84 9F 93 33
 A3 A4 5D CF 5F 29 36 EE 6A 2D E1 F4 D5 18 42 A0
 BF D2 FC 0E FF B7 EA FC 70 21 B0 7D 0E 03 BA E6
 42 73 61 4E B0 D8 62 7D 30 C4 BA 41 12 FC 53 5F
 A5 77 49 41 31 98 13 C7 08 7C 7C B7 7F 4E CE FE
 37 28 AC 6C 39 DB B4 E6 30 5A CD D4 7D B8 B2 23
 37 15 BD F2 64 99 4C 93 F5 D3 D6 9E F7 CD 0C 0A
 B5 AB C7 DC EA 01 95 AB 62 E1 1E 41 27 C1 E7 63
 07 9D 19 21 AA E2 3D 63 F0 0B EB 0F 39 07 D8 77
 AA 12 C2 D1 0B 51 62 98 A3 3A 3F 32 F2 71 B5 CE
 FB 82 1E 42 C4 A0 7F EE 53 E0 7E C9 82 80 9D F4
 88 91 45 0B 54 B4 3F E9 52 FB 11 19 C2 00 2B 06
 25 FC D5 0C 48 72 20 2B 60 7B 16 05 A9 2E D3 53
 14 20 63 51 DA 63 4B A6 19 26 5E 1A 75 82 CF 2B
 C0 DD 88 9F 2E 27 B2 CE C1 39 45 67 2D 1D 8A 94
 01 65 38 05 4E 47 88 BE 64 AA 3C DF F5 50 96 65
 D1 02 61 CF 6E 58 10 30 BC F1 4B 6E 92 DB 70 EE
 30 CC 3B CA E9 98 BE C4 11 B9 D3 69 37 9C D8 6F
 3F 7E 34 E4 73 B6 CD 18 90 9E E3 8D 8A E3 7F 35
 26 82 CB 24 47 93 F7 A5 D8 62 4F 63 3B FC 85 6F
 7D 5F D2 CB 84 A6 CB 88 59 25 DD 8B C9 3E EC 94
 06 78 EB 3D 56 1F 59 5C 3D FE F2 89 18 DA 94 E3
 E7 43 F1 FE B7 28 F9 9A 84 C3 92 46 7F 4D 06 B2
 59 DC 2A 53 D8 11 8E 69 3D 7D 56 33 69 24 6A 2F
 8C C5 7C 97 86 E0 05 8A C8 D0 51 07 1E 47 DE A6
 B0 2C ED 9D 59 5E 76 7D 72 BE 93 7F EB 21 E0 25
 27 78 74 60 84 43 30 12 79 31 B8 B5 7D 91 C6 8A
 10 C7 91 DB A4 2E 7E 85 16 7B 05 DF 5E 30 A8 5B
 00 65 49 4D 14 04 F6 2D 58 12 B4 53 E7 71 E6 C3
 98 14 02 2F E8 2D 3B BF D8 58 BA 4D EB C5 A0 E4
 2C 65 0E B9 29 A3 C6 8F 88 02 48 A2 E1 73 0C 38
 04 E0 4D F0 50 79 4F 0E B3 F1 B9 C4 4F E3 24 6A
 DC B6 CA F0 C5 F4 F6 90 1B 5B 98 2A 2B A4 21 EC
 1A 8E 74 A4 82 A0 4D 73 E5 9A 3A FE 67 CA CB BB
 7D 5E 85 BA 8D 8A F7 1C 0F E9 F0 03 60 AE FA AC
 35 28 26 1F F4 90 07 C5 6D D6 E5 E9 5A 9C AE 37
 F2 E0 AC F8 37 2F 0B 78 06 21 AB 1C 62 1D D8 47
 F7 07 3B B2 F5 68 6B 9C 6F 38 41 26 9A 72 10 72
 AF C1 DD F7 1D 23 1D 33 75 64 26 E7 25 43 C2 51
 8A 23 50 9B CA 43 11 0B 30 52 55 55 E7 F4 6E 02
 B1 6E 42 0C D6 36 6E FF 1E 64 E5 AA B3 C3 A9 50
 52 44 A7 4A 48 62 D2 AD 49 2C CE CF 7E F5 DE DF
 41 91 CC D3 77 FF AB 94 B3 C2 0B 8C 54 A4 D4 53
 5A BF B4 FC 32 89 78 18 DD 85 55 03 3F 25 B4 24
 85 74 9F FB 95 C8 5C C4 99 EC 60 AB B1 8C 57 AF
 69 8D 08 24 A8 94 3F DD 80 69 08 D3 92 2E AB C0
 11 C1 48 8D 2A FD 5B 27 4C F7 DE 1F E5 29 65 C7
 41 54 A3 E6 03 8B 2D 11 A9 3C A9 40 B2 51 E8 AC
 29 2A 8D 16 91 D3 42 31 C4 A4 0A 39 FE 69 AA C9
 D3 50 A3 72 E2 37 DB 3C 97 9E 4D A2 2F 84 C4 0F
 01 7C CB ED 1E 51 F8 C9 FC 9D A1 3E 35 79 AA 5C
 0A 23 B4 06 86 28 AE 4E EE 6C FB D2 C9 AE 9F 8B
 04 88 CB 97 CF 21 E9 5D 5C EB C9 91 A8 D0 44 0D
 94 74 88 11 BD 82 C6 16 0D EA D1 2F A2 8A 20 C6
 79 3A 6E 24 59 9A 1D 51 31 34 B1 B0 F7 A6 34 C4
 49 31 EB 83 30 B0 AD A4 EE 1E 16 1D BF 28 14 EF
 A4 12 9E B7 6F 77 7B 77 A6 80 A1 1C E4 08 BC D5
 23 F2 12 DA 0C F6 EC 89 7A 02 0C 66 3C 47 4D B0
 6E DA F0 54 75 F3 98 16 82 83 3E 94 69 A6 30 DD
 8A C3 56 A6 18 5F A4 DD 59 58 24 9F 36 E6 E2 FD
 0E 25 E3 A8 C8 ED 5F FC 3E 1E 31 E6 86 66 6E A1
 B7 34 D4 C4 1D A7 A4 1D 17 D1 56 3F B4 18 6B 26
 C7 54 9C AF E9 49 19 9C 99 7E C3 7E DF F6 B3 AB
 49 AF 99 F5 79 0F 90 B0 E7 C3 92 32 DE D5 F3 60
 F8 97 59 50 50 C7 16 BD 78 C8 B5 D8 EF F4 88 CE
 13 41 7C CF 6E 74 58 B9 BE 69 B8 42 51 93 3A D4
 2B AA 3C B5 72 CF DA 89 9A A8 6B 0B 72 E0 50 E6
 AB 7D 3E C7 6A 7C CC DD 6A C2 61 4F 7C 8E 69 6F
 7B 15 CB 41 D1 9A F8 17 6A 73 83 04 70 E2 2E F2
 33 48 52 7E 2B F6 F9 46 C0 89 46 71 F4 5B C8 9B
 E2 7F BC D1 BF 65 7A 1B 1D 8D 07 8D F3 2B 4B 1F
 ED 26 1E 66 3C 0A 60 2E E3 28 E4 7B 40 AF 95 3D
 D6 7C F9 45 EC AC A2 21 9F CF 45 05 91 32 DA 7F
 28 4C 1A EB 2A F7 36 4F 83 60 81 83 E2 11 01 57
 1C C3 D3 97 84 E5 20 77 A9 DE DE 2C 78 45 93 95
 ED E2 9C 94 53 42 9A 64 5B 5B 50 72 8E EB C3 A4
 D2 7F 6F DB 09 F1 A5 7A 4C 80 56 D6 38 70 12 F6
 75 E8 BD D7 AB 8E 3F 86 47 A1 E0 B1 B6 74 8B 39
 70 8C AE 77 30 04 F7 97 27 24 05 63 18 AC 8E A7
 D5 9C 59 0C 30 64 89 F0 2C 76 7C C2 22 A6 DC 17
 A6 4A 3E 0B D1 C7 7C 44 DE 62 8D 04 16 A9 37 9C
 DA BA CD 5F 50 9B A8 1D 13 A4 F6 47 21 15 0C 44
 65 1D B9 D6 FB 12 5E A2 1F 04 1A FE 43 B1 17 91
 CC A2 C2 5B CA C7 DB 33 99 CC 3B 52 DA 50 67 8D
 21 43 FF 40 16 2A 19 BF BF 68 9D 92 22 45 CA A4
 EB 4D 3B D3 EF F2 DF A0 89 50 D7 9A 69 4D 7E BD
 05 BD 02 AA 07 77 25 21 7F 32 68 EF 10 4E 8A 2F
 A8 B3 12 B1 35 F0 C3 5B DB 27 C0 D0 DE 9A BC 22
 4E 9E 32 2C F8 7E 19 32 7F 9F 33 71 72 F6 5E 5D
 B7 AA 8F 8E 46 DE DA 26 F4 D0 5B DC D9 DA 4E CB
 FE 57 BF 57 FF 77 73 D4 46 18 7A 7E D7 0D 5D 7E
 C8 6E 63 74 B5 A6 F1 91 92 9E 3D 00 C1 EF DC E7
 4E 84 99 95 51 08 E5 C1 59 BA C8 FC 91 3E DC CF
 32 9A DB DA 0C 5D ED E9 19 79 2A 89 8C 65 7B FB
 A4 45 4A 85 B1 8A 12 3C B3 FF 89 33 82 8C DB FF
 D4 41 96 D6 2B B8 C3 39 79 54 EA E2 7F D1 76 01
 98 DC 75 D4 38 61 C0 00 CA 83 04 92 0B 40 AA D9
 EB 72 F4 73 B5 B9 43 98 B8 8B 65 BE 85 A3 5D 09
 70 71 ED F7 3E 2E 0B 9A 64 5A 6F D1 F2 7A 28 CC
 16 EC 7C 50 AE E8 E6 35 93 F3 F5 92 25 C8 65 2B
 D8 C0 42 93 83 50 59 4A 12 D1 17 E5 A4 42 19 D5
 A0 87 69 76 85 6E 4F 82 5A BE 59 78 08 ED 7E 72
 EF 07 8D 63 39 E0 2A 79 44 EA 74 A3 78 6F 5B D9
 F8 70 20 B3 78 20 E0 AB B2 FE BD CB 8E 9E 92 F4
 DA F4 B3 56 A5 23 A6 04 7C 86 64 E2 B1 BC 64 60
 30 AC E7 0A F9 96 24 03 69 B6 AD AA 0C 98 F1 D8
 1B 73 CD 04 D8 B1 CD 79 44 0E 1D 56 FB 4F 82 4A
 EE A0 B7 53 87 64 44 4D 81 5E AE AC CC A4 9F 93
 C1 88 45 01 57 D6 F6 90 DC 35 6D 24 96 C8 EF 07
 51 D3 6A 4A B1 CB F8 FB 30 A6 D8 1A 69 92 FD 6D
 73 31 FA 03 86 B2 8D 38 C6 04 1E 72 4F 72 63 0C
 2E 0D 64 7D E1 02 3A 80 BF 87 30 10 43 B3 15 3D
 3D A1 F4 EF 1F B1 97 90 14 0E 8D 80 E7 1C F6 AA
 1B 34 A1 E3 20 73 F3 9F 1C 61 5D 6D 75 53 88 D4
 00 5E E8 EE D7 3F 5A D2 9C 2F 4B 4B EC 6E 74 56
 7C 7C 51 CA 4D 2D C8 08 3D C7 7C 4E C4 60 47 15
 47 F0 D4 B6 59 7F D1 1B AB 9D 28 39 16 EF 1E 8D
 ED 3A 2B FD 57 36 4E 05 CD C0 90 AB 16 1C 3C D7
 F0 4A 4A 87 5F 58 9A 12 0A F7 D8 E9 12 2E C7 44
 50 4A D8 B6 6E 50 B6 97 FF 55 EC 1B 4D D3 4E 4A
 E1 EE E1 7D CF 44 F1 16 E7 5F A4 00 24 69 AD BD
 C6 E3 1B 91 29 7E 37 4A 0D 43 78 72 34 C7 D6 8A
 53 C0 FC 7D F6 E8 6C B9 E7 CB AC 5C 65 CE 99 47
 D3 DF D3 EE 55 CA C4 DC C0 5D 45 B8 83 C7 94 55
 E9 9C 2C 56 8B 09 DA EB 3B A3 D4 AF CC 1D 49 77
 DB B3 98 FD 0F E2 12 D1 9D 23 94 49 FD 9D 08 5A
 51 8D 7F EC 29 A3 11 E6 46 43 34 83 91 4C 69 68
 52 17 91 FC BD 02 64 4E 66 49 B7 11 86 65 5C 56
 1D 57 7B 4B CF 7D 9D DE D0 FC B1 A1 36 0D C8 93
 84 A0 B3 D6 DF 62 81 C1 5A 77 A2 ED 66 6E AB AE
 4E DD A3 22 32 82 28 90 9A 3D 9A E4 2D 7E 63 F6
 E8 5A 34 4C 9A E1 52 93 74 E4 84 6D 8A E0 DA 70
 2E 04 99 69 24 03 F8 86 F1 E2 D3 2B E1 3C A2 02
 C0 F0 8F AE C2 1D 77 97 1B 8F 79 45 90 75 9C CA
 DF 45 CA 73 95 65 09 34 0A 74 3E A5 21 8D D1 CA
 2A C4 B8 E2 EB 2C 81 C2 B3 7F 12 79 33 8A C4 D5
 F0 7A 5F C5 29 23 A7 82 45 3F 63 21 CE 92 78 9A
 8B 2B 7A B9 CE 17 CB 40 F1 0A 82 CB F1 11 9F EE
 DF 65 99 AB 3E 2E 86 8E A7 72 80 C7 D6 86 CA 03
 04 6C 35 A4 6E A1 8C 32 D7 4B F6 39 A6 28 15 F1
 D3 15 B7 EE 6B F2 A5 06 FA 45 91 7B A5 BF 2F 88
 9F A4 1D 0C AA 29 A6 C7 C8 DF 0B A0 E1 05 9B 33
 86 42 72 CF 61 D8 0C 2E 9F 81 EC 00 DC 06 F3 7A
 03 94 57 B8 26 78 D8 98 03 08 90 2D 50 55 AA 32
 BA 18 FE 4D 9A 51 A2 A5 FA 83 B9 93 E0 35 68 A0
 E8 07 3E CA AF 2A 52 26 DA 6D DB 3A D2 3F BB 89
 30 56 C6 D1 02 CE 9F 7A 8F B7 41 71 3B A1 89 8F
 85 BC A1 84 E5 C1 2E 4E 1B 9D B2 7C 16 EB 0A 9F
 93 51 C2 AC F3 D0 85 F9 16 ED 7F 68 78 56 34 B3
 D3 6E 62 BE AA 2C 37 12 1B 45 E2 84 70 3D 4A 59
 7F 27 7E 57 68 A0 EC B8 BB B1 CA 5C A0 F6 FD FE
 87 2C 6D B7 53 ED 97 86 AF 6D 01 E1 F1 10 0E B0
 12 5F 59 7C 89 9C 68 E2 E6 A7 A6 39 18 E3 E3 AB
 BB 21 2B C7 DA 2E DA 1B A0 BD 9F F2 12 A1 19 58
 42 DC C9 EA E5 96 B5 EE 0A 49 B6 17 26 F4 13 F9
 C2 15 C0 ED C6 AB 41 A2 77 0A 3D 1F 22 A8 AB 56
 0E 8B 7B EB 29 C3 71 98 CA B5 01 8C 74 67 5A 72
 73 23 93 15 18 48 CA AE 61 13 07 D8 D6 87 C4 44
 F5 BD DC 0A B0 24 E1 94 06 4D 68 A3 DF 5E B2 44
 91 98 C3 54 7E 97 F1 CE 20 B9 51 48 F6 7A 07 28
 24 F1 C9 3E 75 17 AD 14 43 62 8E C8 2C CF 12 0D
 D4 D6 DC 82 86 68 62 42 BF 28 B9 AD 32 9A B7 98
 65 32 A1 99 0E 36 11 25 DF 75 96 43 AB 0E 5E AE
 00 98 D4 C5 FE 07 3D 1F 7D 8B DE 3B 69 36 35 CA
 BB 2C DC CE 77 EE 65 FA 63 66 54 F6 0A 89 8E FD
 D1 60 36 3C 30 2E 56 4E 25 CA 32 58 C6 38 0C C7
 D3 CC E3 8A 25 BD BD 83 5B 6C 0B 6B 28 19 7B 55
 02 15 D0 22 AB 76 13 0D A8 9D CF 2E F0 73 14 75
 1D F9 C5 35 12 72 E4 45 5F 6A D1 E5 24 A6 38 F0
 44 0A 11 CF E6 3D F0 62 4C 59 EF 8A 86 D9 D4 AF
 C0 09 F8 1C B5 76 D1 89 C1 01 B5 D3 3B 88 B8 7B
 63 30 95 F4 69 38 FF 9E 57 76 04 44 D8 EF B1 8E
 CC 2B 09 F1 34 26 E8 4E F9 90 63 A4 B1 00 CC 62
 BA 21 FF 94 55 53 BE F7 1D 4F 7C F2 83 FC DE DA
 44 CF D5 12 0A 5F D4 60 74 D7 71 98 E7 EF 0B 79
 CF A4 ED D0 4F 50 9C 4F 02 BC ED 9E 67 73 A2 CD
 FB 1A FD 65 C5 77 6B 70 4C F7 76 DD 32 A0 35 14
 0D D0 02 B3 D9 7D 1D 70 94 89 5A DB 66 FE 96 4B
 C0 49 01 96 52 6F 8B 9F 3B 69 17 CD 49 6B 81 30
 E8 2B 9B 66 D2 B4 54 60 C4 BD 65 C8 8C D6 0A 61
 A7 9E 32 0C 30 47 0F 9F 3E A8 6B 15 5E 57 D7 EC
 73 1B 0F 0E 6C 92 36 B4 36 26 F9 BC A5 A9 5F 45
 25 DE 78 46 73 99 06 A3 65 BF F5 24 95 57 6C DF
 D2 E4 28 08 D2 A0 8F 73 53 18 CD 1B 8D 7F 5C 2B
 03 90 AF 6D 40 34 65 82 7F DB 5E 0B 95 05 CC EF
 46 54 5D DF EB 34 25 BA DD ED FD AC 82 99 84 F4
 71 19 79 73 F5 29 7C 92 DE 70 8B 36 3C 05 6B A0
 39 B6 A1 77 3D 91 3F D9 60 F6 4F 96 42 A0 A4 CE
 4E 27 01 1F 8A 87 FF CD 41 DF 60 02 9C 7E 96 48
 E1 4B 8D 34 65 CA E9 B3 7B D8 1D 36 E1 AF 32 1F
 97 C7 A0 E8 3F 89 AF 69 3F 45 E1 6B 66 1D 8A B3
 8B 44 32 CE 58 A7 71 0E 74 27 A4 7E 35 58 72 76
 2A E4 4C 6F E2 38 0D 03 A5 4A 06 4C BA 08 44 E0
 B7 A6 B9 9E 09 47 FE 0E 5E 2A A4 96 7C 09 1C AF
 A2 74 AA 17 83 D2 43 D3 3D 91 48 B4 B0 A5 3C 73
 27 24 07 E1 6A C6 B4 13 08 67 FE 69 B2 45 2C 68
 45 B9 3A 29 A0 59 87 89 57 A7 DC C3 0D 01 C5 9A
 2A AA 97 AF B3 AA DE BC 16 C7 F9 2E F1 F5 5F 2D
 BD 25 B3 EE E7 92 9E 19 23 C2 FB 39 2B 4D 3D 06
 E8 D6 CD C2 1B 68 2B A8 43 62 14 53 CA DB 0E 4B
 56 41 4E 66 85 34 27 DF 5B 31 A9 58 77 F1 5D A1
 72 8E 87 9D 2D A6 E0 76 C7 CF EB D8 37 D7 40 D6
 5A B5 BC 0B 6D 0E 1E 37 63 22 6E B9 76 60 70 2E
 71 AE 58 BA 1A 58 67 56 A2 18 DE E0 AF E1 EA 48
 8E D7 98 A7 6C 70 FB 40 79 AB 76 5E 60 8C 15 55
 D7 97 37 E3 B9 14 7A 3D 57 8B 07 B2 EA 92 C5 79
 68 1A 44 66 6F 67 41 E6 05 0D 6E C7 3C 06 56 A8
 4B 52 52 75 45 B8 81 56 E3 76 96 C6 00 27 26 BE
 14 09 93 10 A2 2D 4D 38 9B A7 2D 65 62 9C AE C2
 AF 98 B4 3C B6 0B 84 B6 8E F0 0E 26 8F 0B 60 DE
 BD E3 3D FA 5D 9B EC 46 64 D5 9B EC 5C 6E B5 3E
 96 BF 60 0A E8 74 91 6A 40 B6 21 9B BB 87 8A EB
 1E 24 65 D5 C8 BC 6A FC A2 65 5E 57 0F F4 05 44
 07 C7 B0 BB 51 CB 46 05 E2 08 DF F3 05 02 67 21
 FB 06 57 CB 65 FE 5C 03 56 E0 DC AB 60 95 82 6B
 68 CA A1 4C 0A 5C B3 7A 5A 35 D1 12 F6 3C 19 6F
 C1 74 3C 5F 71 68 D8 D4 51 75 E1 4B 8C 9B AC 0A
 F5 E0 62 AD C3 93 92 96 8B 0A D2 2F 35 0A 56 08
 67 FF 7F 6A A3 31 24 22 EF 14 4C DC 05 B5 8E 2B
 AF D2 68 75 85 2F 78 B2 54 EE F4 6D AE DD 97 42
 BB 46 0C 8C A0 43 FE 38 9C 25 02 52 4B CF 3D C8
 D1 6E C4 5E C3 9F CE 77 87 61 57 D5 70 85 40 F2
 53 1B 04 74 88 C1 C7 41 D9 A8 E8 C9 EA 9C 0F 63
 00 E3 BD B4 A9 8F B1 64 08 CD 34 E0 09 CF 88 F5
 40 6B 20 73 CB 35 6A 99 C7 2F 22 68 4C 8B AA 4B
 E8 A1 69 2E 15 81 A2 56 C6 CA 59 11 F9 85 4F 6B
 7C 18 36 5D 08 D3 60 09 0D 0A F9 C3 1A BC C6 1B
 D8 33 3B C2 AB E3 96 90 69 88 41 88 3F B6 74 C6
 BB 4A BC 87 7E 51 F6 85 86 E5 59 FE DC 07 6A 1A
 A3 72 50 A1 60 19 1C 9D 60 A7 B2 32 57 15 39 18
 2A 33 18 15 6D D1 6A 73 3F 51 B4 C4 EA 9B 92 99
 46 32 44 F8 7C 38 F4 C6 63 F3 00 04 8D 59 3E 92
 E9 11 4C 5F CC B6 F3 A9 02 C7 39 59 B6 9D E3 A4
 98 5A 09 B0 4C B2 33 63 46 B5 A3 7A C5 71 B5 3E
 45 B0 31 B3 29 78 81 48 B8 2B 05 9F E1 3F 2D 3A
 63 AD D0 69 56 04 85 21 47 65 9D 78 A1 B5 99 F3
 88 4C 72 13 65 2F 72 8F EB FB 21 29 04 AD F6 6E
 82 9A 13 78 6C D0 12 43 F5 76 3A 5C 90 E4 45 3D
 D3 14 38 02 E9 B0 9B 13 F0 C2 E7 C8 24 D3 50 85
 E0 38 5E F3 86 F9 88 17 41 5C C2 F9 E4 5B FA 1A
 E9 05 29 56 D7 31 43 78 E3 97 32 52 BA 80 4D 5D
 19 90 36 2E DE 53 1E 27 5A DE CD 0A A7 7A D5 03
 9D 42 89 71 0B 0B 69 43 EA 05 5C 7D 07 62 C1 FF
 C1 4E 2B 1A F8 80 40 79 4F 1B 6E 52 D8 06 63 8F
 DA AB 64 D9 5D EA A6 FB 69 90 BC 5B 46 D1 7B 3D
 50 85 E3 4C CA A7 1F DE 89 F5 B6 73 DB 89 E1 D4
 EC 44 32 0D 74 15 C0 B4 96 ED 8F 0C D3 9A E3 7F
 48 D7 4B B0 82 83 8B D1 FE C5 23 55 DB 0F 39 A7
 90 ED 52 5D D0 62 2D 3A 00 E4 34 89 94 B3 A3 40
 22 47 50 95 75 BB 5C 20 EC AD 4F 2C 08 27 CA D2
 F6 A7 34 C7 F0 4D 8A 48 42 BF 98 13 5F F8 1B B2
 D9 23 A4 49 29 B2 74 BB B3 48 50 72 D2 D7 1A E2
 6E DE 57 BA 19 3D EF 39 1F BC E9 F0 72 89 7A 2F
 20 FA F0 3D CA D2 A1 31 4C 02 0E 2B 37 D3 C1 AF
 BF C3 14 38 11 F5 7F 23 BC B1 D3 F8 5E 9C 9E 95
 98 BE 75 62 DE C7 CE FD 17 C4 6F D4 10 CE B6 B9
 F7 93 E5 73 E3 5D C5 6D 6A B3 03 71 F5 8E 1C 9F
 D6 B4 AE C2 DB 4B 11 62 C2 A1 84 CA 85 1F 03 76
 E5 1C 66 1E 52 EE 7F CF F3 A1 16 A3 5E DF F6 0C
 A1 92 D3 B9 F0 9E 4A E7 D9 00 BA 35 90 7D F4 BA
 AF CA 6C 33 B2 D3 A8 A0 F1 0F 21 EC E0 F1 C0 6E
 B4 1F DB 4F B0 36 EB 29 EA 91 D4 24 96 28 81 17
 C6 88 9E B9 DE 01 9C F2 60 74 8A BC 10 03 13 52
 1F C8 D2 E2 7F 04 0B 3C DE C5 43 03 DC 0B 69 38
 D0 A5 8D 05 F2 84 F3 C3 D1 9E 80 04 69 AD 6D 72
 8A 72 73 3D 88 24 80 59 27 D7 39 82 5D 10 2C 87
 55 40 32 10 9C B7 89 57 A9 04 68 FA 92 A1 D5 D3
 EA E7 DD 54 00 26 C2 49 78 DD 77 A6 4B 65 6F 2A
 95 80 F4 D3 E8 1D 83 B1 E3 2A F6 8C 14 A7 09 69
 66 8E A5 10 60 D0 E8 81 AB AC F0 2C 34 25 E3 C6
 6E 9E 6B 97 97 44 F4 D4 53 EF 48 58 92 C0 6D 48
 26 AE 13 CC C0 66 BB 90 C8 7D 6A 3F 3D E8 1C 15
 7E 79 6C 3D 42 4E A4 E9 4A 27 59 EB C8 86 93 90
 8D 18 0B E0 4A 8E D3 D2 7F B5 3F BE 90 71 22 54
 73 D2 FB 0F B9 31 98 96 23 2A 2C 55 CF 3D 98 D8
 44 00 4F B9 6C 6D E0 38 45 E7 DE BE FA 7B 3A D2
 FA 47 12 F2 C3 31 3B C1 E1 F0 42 F4 1E 5E F7 A9
 77 3A 68 C0 ED 1F 73 57 EA 93 F9 C8 B9 FD 63 A4
 41 26 6E CA A6 1C 54 A6 C2 D6 F2 7F ED BB A7 35
 18 93 00 54 30 04 C7 A0 E1 02 B6 CA BA 53 54 57
 95 FA 64 B2 C1 EB 49 32 62 52 27 41 55 E8 A6 94
 EF 25 89 E5 B4 5C 3F 96 9B 91 26 A4 BE 3C 20 C8
 0D 6E 57 65 ED 02 F1 74 56 81 9B 29 E0 51 53 FC
 6B D3 4A 9A 50 81 F8 82 B1 D0 C4 09 E5 28 D9 DA
 0C F8 2E AC CE 23 9F 5A 3E D0 F7 B1 0B DF 07 22
 73 6B C4 E0 1D 1B F0 02 A2 50 FD 25 18 9B B4 9C
 59 E5 4A A4 15 16 A6 F3 55 70 45 94 7F DB B1 7D
 CA C3 63 FD 24 80 06 8C 27 AC 41 7A 91 50 76 BD
 4D 5A 84 8F CA B4 DA B4 E9 2A CF 50 A8 B2 62 A5
 1E D3 71 1E 4B 83 E8 87 29 C1 FE 2C A9 1F AA 1D
 82 26 D0 12 70 E4 57 85 A5 11 42 64 7D 97 0C B5
 13 E0 77 4E 4B BD AC A0 98 F4 60 2B 93 33 5E 8F
 86 F4 24 18 57 78 9B DB A2 A6 04 8F 81 9A 9E 40
 94 71 C8 25 EA EF B0 FF 3C 02 D8 62 58 0F 1F 9D
 59 47 3F DE 97 B9 61 47 2C BA FA BB BD 79 28 C1
 E8 7C 2A D5 2C 93 44 99 4B 63 9C D6 4B 6C 6E A3
 E6 9F 1C A7 05 C8 77 5E E4 04 DD BC 83 17 5F 4A
 1E 93 C8 56 30 69 14 F5 E3 23 97 C7 BE 27 03 00
 82 FE 95 2E A4 46 7C C1 72 27 06 72 E2 A6 81 8D
 2C A8 89 F8 63 2C F5 CA 5E 49 63 4B 0E B7 0A B1
 BA 22 45 A1 55 61 3B D7 8A 85 EA 90 22 B8 1D F5
 6E 25 6B C5 10 9D 7F 7B 6B 87 89 7B 0C 82 3F 63
 0F DE 8F 63 FD 33 48 48 7D 9C 88 3E FE 5A 3F 5B
 9B 89 A2 C0 0C 68 EC 79 3A A8 78 02 B1 4F F7 3A
 F8 3C DF A8 5B 3E 52 F5 DD 65 7E 7A 27 F6 C5 6B
 3E A5 72 6C 71 C6 14 4D 89 12 12 5A B5 AB 18 C8
 74 BB B3 11 A4 77 F8 A5 CF B9 4F 3D 1D E0 D2 74
 BD 1F 6D AF 12 A7 EF 0F 3D EA D0 00 60 2A 4C 19
 DA 5A 46 CD FF 0B E5 A1 D4 B0 2A 57 CE 70 75 AB
 4E F6 EC 24 74 71 AB 97 17 02 04 0D 51 24 DD B6
 B4 48 39 20 0E 23 8C BE 4E AA E3 B0 DD 37 61 D7
 78 E3 68 3A BE 8C 17 9C 1B 96 85 37 F4 35 9B DD
 E8 3A A5 B0 7F 84 F1 A1 2A 43 A6 54 41 FD B3 F1
 60 46 6B 1F 05 CF 1A DB 11 15 82 49 78 8C AB AE
 97 98 C3 43 D3 D4 9D B9 67 5E 9F 3D A8 62 ED 43
 68 4D 9C 7C 1A 87 0D 3C 98 4D 77 27 8E 57 E5 E3
 A7 0D 5D 70 F0 BB 23 0A 98 68 42 88 AE F4 DC 4A
 AC 37 AE CF 31 52 A7 60 A5 D8 2C 6C B4 B0 01 C2
 31 00 0B C3 CE DE 67 E2 8D 6B 22 4D CA 97 FE 7B
 36 C9 06 58 56 56 28 C4 98 4E BB C7 E7 DF 15 CD
 45 58 49 6E 5D 6F 85 DE AB B9 1E DA 7D EA A5 E2
 73 EF 56 99 DD BE A0 CE 88 12 B6 7C 75 3E 03 18
 F2 3F 57 73 DE 6D 28 EA D3 A2 AF AA 92 51 35 5F
 A1 E2 DB F5 B4 37 69 0F 2F FC A1 14 8D 3A 06 FE
 64 84 C0 59 25 1C 9F 99 B2 3D FE 19 57 76 35 1B
 1B 61 11 EB 09 A3 A5 61 B0 23 77 36 94 1A 9F EF
 9B 89 1E B8 E4 10 5C 25 ED 76 0A 1E 56 C2 E1 49
 BB 6F 37 73 71 06 20 47 BD F1 F6 8A E2 3B A1 BE
 FB B2 52 B6 83 93 7F 5C 5E 4B 67 A3 26 60 47 83
 9C DE C7 10 61 BB 2F A6 09 0F 1B F1 95 D9 D7 B7
 D8 BE D3 14 B8 78 EC CE 9E E0 3E 2D 32 CE B9 9F
 03 84 54 49 80 ED F9 CD F5 9E D3 07 13 C0 B2 D2
 1C 84 66 58 A2 D0 55 2C C9 9A 7A 03 9E 8C 86 AC
 67 C2 4B 95 3E B1 17 76 07 D3 E8 B2 1E 77 CC 6C
 4C 96 69 F7 A3 C8 3E 6D 3D 4A 4E 81 E0 81 6C 9C
 44 1C 3D 2D 8C FB 89 97 DD AF DD 04 6B 6D 87 2F
 1F 3C D1 ED 20 80 77 A0 CE EF 1B F1 BA E7 56 B3
 BD 90 EB 34 ED E3 75 EF 67 B3 19 19 98 25 BC 60
 CA 1D 95 B5 80 77 D5 91 1C BE B2 ED D6 25 C9 33
 55 5A 90 80 E6 78 6D 88 65 4B 27 A0 09 B6 43 FE
 0E 23 6B 69 C0 5C BB BB 76 8C C0 D5 B5 AE DE AA
 40 77 B4 58 D7 D0 2C 32 64 12 92 E0 0A 15 12 94
 23 D5 B4 59 4C F0 EF F7 8A 6E FB 3A 73 2D BD 90
 39 47 52 60 CD E2 2D 2C AA 8A F8 1D 55 46 8B 92
 9D B1 8C 51 14 D3 8F AA 04 53 3E 67 68 80 C4 CD
 52 4E D5 BB FD 97 89 58 C7 CD 60 71 87 C7 F5 35
 F0 7C D5 6E 89 20 75 C5 4C 38 1E 22 E0 12 86 1D
 06 67 F4 75 96 FC 32 F4 8F 8E 48 83 70 5F 86 FA
 9B 30 1B 34 50 12 DA A1 C0 37 25 1F B0 AC 99 13
 6C 14 EF A0 3D 47 1F 24 64 E5 E1 63 28 C3 41 FC
 C8 EF E9 F7 34 88 3C 3D A0 7F 03 AF 07 89 B7 D2
 91 E0 61 A9 F1 10 E0 8E D1 C0 69 CA 88 7C 47 27
 AC 0E 49 C4 83 B8 C7 EA F6 EF E6 53 F5 BC F5 9D
 7E 01 0A 57 37 19 98 FE AF 63 5C F0 07 30 46 31
 AB C1 E3 6A 1E C5 54 02 65 C9 F6 0D 72 3E F7 F4
 54 98 6A F7 8E 7D 3B 0A 51 C6 19 18 CB D2 08 51
 8B BF 74 34 79 63 E1 4F 4F 4F F3 50 1B D0 A9 7B
 4A 87 8E 74 51 87 75 D7 B2 AA DC 49 E6 F7 9C 95
 34 6E FB 8D CB BC 55 C9 EB C7 5D 19 DF C9 97 7E
 2D 45 6A 6F 1B 6E E7 73 95 EA 56 E5 2E 85 F1 5D
 E5 A1 5C 54 2C 3B F3 70 D3 28 45 09 99 8B 2B 19
 18 49 4C E4 FE 70 3C 9B 46 68 E1 5C 51 DE B5 60
 55 53 78 A2 48 78 BD C8 41 FE AD 98 42 EF AF B3
 E9 09 D0 99 25 68 54 2B 84 07 19 98 5E F6 DB 67
 5C 96 5C 9D A9 56 FC E5 ED 37 24 72 91 A5 56 B9
 D8 FF 78 0C 47 C0 65 78 E8 E8 D4 05 A9 45 14 8C
 A7 69 E9 5A D6 56 7C 81 B0 38 8F 0E 29 E8 B0 DD
 C8 51 32 9D 20 4A 90 C3 AB C2 93 82 E7 C5 40 09
 98 61 8A 05 EB E2 9A 30 08 DF 15 4C 55 43 2E 9D
 F5 2D 52 C9 10 19 1B 63 52 C7 52 1E 0E A0 94 D2
 E2 46 46 20 D0 BA 4A 4C 12 E5 B7 3E F5 BF 54 E7
 77 01 2D 03 43 8D 48 C7 6D 83 5B 2C 07 D4 D0 CC
 A4 C4 34 D7 3E 7D AD A5 39 C3 00 E9 65 1E F0 1E
 DD 9C F1 5C 06 3E 3D 0B 31 B7 B5 6B 6E 25 97 B6
 2E 4F 90 F6 00 E9 04 76 F1 3B DB 85 4E F5 C5 2B
 51 D5 87 AD 03 89 10 C2 DC 2F A6 71 A6 A9 44 13
 F4 FF D8 FD 21 AC 40 F2 81 39 14 88 40 69 19 5C
 B9 69 9A CE A0 15 AA 91 1C C6 28 74 12 50 03 45
 2A E8 91 64 CA 24 BB FE CA CE C2 86 21 1A A4 58
 BF F4 EF 14 9F 7A D5 D6 DD D1 27 F2 E5 B9 B2 30
 15 97 D3 F3 AE 05 5E 3D 36 10 E1 7F 4E B7 52 24
 6B 88 55 70 63 AF E5 56 47 86 B0 59 DE 17 5F EC
 2C 2F 18 46 82 96 E8 CD 5F B3 E2 F0 98 5B BA 32
 6F AE 3E 52 EB 20 7C 33 76 8F 56 F1 0B E9 E4 D0
 1A A7 76 E6 A2 AF AE 6F 4E A2 7F 29 E3 D4 FB 0C
 32 23 EE 1A 62 0C F8 19 AC C3 6D 54 65 FA 6F 85
 44 70 95 D2 8E D7 C8 16 21 09 65 CD 71 CC 1A C7
 97 88 7E D3 71 91 9F B6 FD 2C B5 7D CF 85 CD A8
 09 7E CA 28 D9 55 2A 10 46 C6 6A 29 38 B0 FD EB
 3E 87 99 89 4B 25 3C 4D AC 3B 29 0E 30 8F 64 4E
 92 79 F4 BC 20 EF C4 45 5F 28 77 6E CA E5 C4 5D
 4F 09 E3 C3 58 33 27 8A 68 F8 0E 8F 9F 9A E5 D6
 A9 0C C3 5B 0F 31 C5 D1 7D 95 FB F3 95 88 16 8A
 90 02 FF 0D A2 E1 31 30 AA 0B C3 0D DF F6 05 78
 F7 51 E0 A2 ED C2 DA B4 8D A1 A4 AC 69 BB 41 D5
 8E 66 4C 98 69 3C 09 EA 76 20 5E E7 4B 37 B4 DC
 9D 86 3D 58 40 8C F0 CF 68 E2 56 7E 58 C3 41 0F
 7F 68 84 11 05 5D 3E A0 A4 54 3E A1 41 36 B4 A9
 9C 7E 07 72 46 09 DE F9 12 15 A0 90 C7 A1 B4 96
 6A A7 5A E3 00 04 86 78 69 26 1E 7D CD 38 16 B5
 32 9C BB C9 2A F4 D0 8C 76 29 33 F1 EC A6 16 0E
 79 DA F1 7B 3A 65 9A D0 08 89 00 4F 18 3D B5 D6
 69 53 35 5E AD A1 67 85 83 1D 4E DA F5 C4 8B 1F
 DF 35 7C C2 AA 2A C7 7D 86 BB F6 BE 8C 4B 09 86
 BC AD D4 69 7A E7 C5 50 4F 9B 52 E8 0F 5F CB 8D
 59 AE DB EB 54 48 25 EA E1 18 E4 0F 28 42 81 66
 C7 B6 E5 54 AE 41 B1 98 4C 3C EC AA BD 9B 0E A3
 EB 33 1B FE 22 94 47 EF C0 9D 39 71 BD E6 08 6F
 5A 00 DC 82 5A 12 4E 05 E1 46 0C 5D 23 63 01 0F
 29 86 24 1D B9 D3 59 C9 89 5F AF 65 68 6F C9 39
 DA CA AF F4 A5 A5 72 1D 16 C8 93 3A E2 B4 1F 29
 7B 1C 1C CE 28 FE 97 A0 14 42 DC 0B 51 D3 21 AD
 E9 56 38 A2 13 D3 BA E9 10 51 69 CB E5 25 0C C5
 6A 0B 9D BC 02 87 7F A9 51 43 EC 89 03 9C DD DB
 0C E3 72 D9 61 07 F6 C7 81 43 52 94 58 C3 F5 8D
 BB B6 86 AA 4D 85 7E 24 F6 71 A0 AB 6E DD 19 C7
 9C BC 0B 27 EE 2C 61 9D E9 62 85 08 B5 A3 3A DA
 BF 6F 6A 9A 37 40 3F C5 9B 4C C7 7F 1E 73 02 C2
 F4 FA 89 B5 24 81 27 91 66 4E C3 35 ED 1D 07 4A
 32 97 93 80 79 12 50 6C CF 55 4F 23 CE D2 67 20
 3C 83 E7 74 B3 8A 77 CA E6 B5 00 63 02 91 26 5E
 1D D0 4A FD 13 C7 86 4E DD E6 9D 6F DF EE 4D 90
 21 BC E0 EA 2A DD E5 21 F4 24 59 F7 7A B2 2A 6C
 19 3D 50 2B 2B AB 5F 6A 4C B6 FC 9C B1 C3 C0 43
 FA 27 B2 26 E3 F3 0D 3E 3D 9D E1 D8 E2 E5 E5 71
 6C CA 34 F7 23 B8 6C F5 5B E3 D3 C0 85 B8 BF 5F
 6F 91 31 F4 67 B9 78 B4 54 D7 36 31 36 0D D9 CE
 09 9E 57 9F D6 F4 AC CF 27 AE 91 98 60 58 97 0B
 8D 53 84 63 06 CF 31 4A CA 86 D1 32 74 85 72 C3
 21 A1 22 35 91 E2 36 EE 45 EE B7 04 F0 6D C9 FD
 79 30 A8 3B B4 48 53 68 6A B7 1D 28 DF 25 E9 B1
 1F 49 05 8F F6 5D A8 92 1F 8C 3B C1 E4 B8 B3 CB
 DD DC B4 DB 4B 1C 7A 22 46 E8 42 89 4C 4C 25 30
 A0 7B 15 46 15 EB B1 AC 03 49 B5 BE 48 B2 7E AE
 13 1A 5A 8B 66 CC E8 7A 10 97 90 F1 CD 9E 97 6E
 E9 52 C5 FE C4 59 99 45 8D 8D 01 C7 D5 56 D9 F5
 22 03 9C 0B 05 C6 3F AF E6 D0 ED 39 01 C3 91 BD
 6B 34 C3 6D 57 E9 00 6A 89 07 8B 80 5E 0D 48 3F
 B3 04 6E 68 9F DC 83 3B 8B C7 0E E4 2A 6B 2D AF
 36 94 63 E5 AE FC 21 77 11 8E F8 3F A2 E6 17 7F
 4B 4D E0 9A 5D 5F F7 D2 17 12 CD 1D A7 86 E0 2D
 9A 92 9F 9B 6D 31 AA C7 54 CB FA 70 8D 42 10 7D
 DB E6 60 6F 73 1C D6 5E BB 33 BD 44 29 A6 B1 7A
 99 AC 2A 35 A4 B5 AA 6E 76 68 C1 51 E9 E3 0F 6E
 34 29 9D 71 68 4C 50 35 95 CD 81 68 B6 07 BB 43
 29 FF CE 32 66 38 A4 94 1F 09 05 49 C8 A9 16 49
 E0 CB 5A AE 10 2B ED D2 BC F2 C7 C1 F0 75 F1 21
 3B 20 3E FF 62 1E 47 ED 1F F5 46 86 59 21 71 8C
 AA C3 9D 50 E4 2B E9 11 BA 51 EC 06 2C 8D 98 AD
 17 8D D5 3A 48 D6 A3 FB E6 AE F2 B1 96 20 C1 6B
 B3 27 54 08 29 66 6F 2B EE F9 26 D6 D9 07 61 03
 72 DD D5 45 C1 74 75 D0 C5 41 83 6D 84 26 CD EC
 23 44 2A DE 30 0E 79 EA 4B A1 E3 0E DE 21 68 76
 1D 60 7F 57 E0 C1 76 E2 F5 A5 12 4D 4B 1A 1B EF
 CA DA E7 FD 18 C1 E4 D9 A3 21 CF FF E1 E1 60 6E
 57 6E 6B 34 F8 E6 B8 4B CE F6 22 FE CB FE 16 66
 E1 E9 1B 8F 6A AE 17 70 B2 59 61 CD 02 59 85 7B
 D3 92 9D D3 ED C3 45 AE B3 2D 2A A4 BC 39 A9 9A
 65 5D 06 A8 52 2A 05 76 4E 5F 70 62 BD 78 5C 85
 75 BD 3D 9F B3 55 9B A9 AF 16 B6 9B 2A 6D 2E 05
 66 1F E9 2E F1 97 E1 C3 3C A6 F3 E5 CD F8 68 8E
 7E 9C 50 ED CE C6 C2 DB 5B 10 AD 70 48 47 A3 AD
 F5 58 21 32 DC DF A2 44 15 D4 68 0C D2 C3 A5 4A
 C1 A3 FE 14 8B 6E F8 58 B5 94 D1 20 5D 6D FA 73
 76 35 27 19 70 E1 8A 50 BA FF 79 D1 7E FC B6 3E
 05 E6 48 58 61 64 61 2C 89 C3 EB 5D F0 D3 0A 33
 11 65 2A 1F B8 26 02 CB 85 86 13 FB FA D7 F2 C5
 DC 53 BC B1 C4 9D A4 E9 D3 31 F2 DB A5 FC 4B 06
 56 B8 8B 95 4E D1 38 35 C0 10 A2 EA B1 A3 36 F0
 CE B0 FB 75 27 3E 43 E4 0B FB C5 EA F6 12 27 B1
 F9 8B 6B 2D FD 3C 34 7D CC 30 46 B3 0A A4 F8 7B
 D3 95 6B F7 E8 2B E6 2B 3B 01 67 C4 36 4F FA E4
 90 40 E0 85 32 3F F9 E6 DC 86 5B 4B D7 FA 06 DF
 4F D4 D0 45 9A 52 95 24 59 4B 98 9C 87 2F AA C0
 6A 7C BB 05 1D 71 5D 58 5C 2F DE 05 F3 F5 56 90
 CA 5A AC 82 DB A8 29 69 9E 00 72 7B FA 65 AD FA
 68 C6 FA B0 A1 60 42 4F 87 13 5E 61 75 10 62 5E
 6E 6D 45 4B F4 BC B1 00 5C C2 86 75 05 A8 C9 4B
 70 2A 55 95 24 06 73 BE 4D 3A 4E 65 E6 4F C5 E6
 E4 97 10 E3 9F 8C C3 7B A0 FF AD D2 D6 72 74 2A
 EC 68 1B 7E E9 63 AA 3A 12 8E B3 64 9D 63 CE 50
 6F 0A 6D 3A DF 81 79 4A 75 B1 D2 6D 86 5A 03 15
 FD F9 13 70 5C 6E 89 26 F0 7E 24 9C DF 79 1A 65
 F1 84 2F 69 3C A8 25 53 05 7D 9A AB EA 40 01 36
 D0 9D B4 2C C2 6A 08 09 81 B4 C3 C7 8E DD 55 C2
 FE 96 05 FA D5 88 55 AD 85 C1 9B 77 90 24 30 A1
 6B 19 6D 96 9B 30 29 83 D8 EC AB 46 B3 0E 5C 84
 88 06 ED 9D B8 57 AF FF 96 48 93 2C 5A 66 CF 49
 BA 8C E1 D3 5F 9D 08 D9 9D 55 EE 71 0F 88 BE A8
 92 CD 2A A9 71 DA C0 DA 51 5D CB E4 A3 FA C2 F0
 4F C1 17 E4 F0 85 6F 37 26 26 3C 96 C5 C5 C1 87
 5C 02 F5 5B 01 DE 07 C9 E7 FD 02 A2 54 47 95 CE
 97 2F 33 D1 6F 73 39 32 4C 2C E7 49 75 1A 16 45
 0C 37 F3 9C BF 2B 68 8B 1C 71 B6 FF 68 F9 56 E9
 05 99 30 8B 4B 68 5A 2C 14 FF 06 D9 C4 FA DC 27
 AB 67 0A 58 52 DF 81 4B A9 FB 86 AC 9E F3 70 B4
 50 A0 98 06 98 BA 95 EE B0 ED DE 02 9F 99 57 79
 E1 07 86 AB C6 1C CB 53 97 3E 52 EF 78 FA 5E 16
 66 79 F9 7B 20 22 D2 2C BF 5A 80 B3 1C B6 EC 1B
 91 0A 38 1C 65 0C DB FD 81 2B 22 49 ED 98 DF DA
 43 F4 17 C4 BD 1C 3F 8B D9 DB 90 6E 9A A8 91 EA
 37 62 58 9A 7F 60 AF BE D1 90 19 26 8E 3E 7E C4
 C7 2F 8D 37 6F 78 03 FA AB 19 5F B2 AF AF E2 9F
 A8 1D A5 EC 67 8A 75 4B 6E 7B 3F 8D 82 D2 23 81
 6D FA 5C 58 DA 9D 7B A6 EA D3 85 D5 35 74 1F 71
 FA 53 E1 85 82 4B 40 C1 2D B8 0B 9D 6C 5E 5E F2
 EA 01 E6 48 E3 8A F1 A5 20 0C 05 B5 94 D1 EA 55
 A2 13 C6 4F A4 E2 9E A0 3C A2 BB 7C B2 26 DC BF
 EB 87 F2 4F 23 01 B6 2D B8 7F 00 18 7E 55 65 3F
 B0 EA 06 F4 6B B3 84 E3 B2 2D AC 16 F4 0A 64 E7
 70 77 28 02 A0 84 38 0C 12 14 6C BE 1A 87 04 30
 B1 E8 6C BF 25 6B 54 1C 08 45 65 B3 3A 2E 0D 60
 1C 85 BC 1C FC 47 1A 1A 80 58 6D 49 1F 93 BD CB
 D4 55 72 85 69 17 F5 B4 16 1D DA AB C7 EA 20 23
 E3 E7 ED 74 18 8D 60 86 17 33 6D 3F 81 1C B9 88
 C4 C5 03 BA A2 BB 5E 14 88 8E 5E 53 11 DC A3 8A
 86 A5 D8 B9 64 61 43 94 94 B6 12 98 BB 1F 8C A6
 0B 0A 1F BA A0 85 21 1E 6C 61 4C 7C 8E EB A3 B7
 9F 81 86 9C D7 DD E0 9B 8C 02 98 45 A9 0D 42 33
 A4 57 05 01 6F D0 96 64 D1 24 F4 0A 82 A5 FB AB
 6B 02 E2 5E 5C 22 46 36 0D 09 48 39 25 CD 2C 1A
 DF DD 8F 41 95 DD 69 AB 02 05 32 6B A2 76 B1 CD
 4E A9 20 EB 78 F5 C0 9E 28 21 BA 6F B4 14 A7 33
 CB 73 CC 22 3F 2B 65 7A 78 BB 74 57 E0 57 52 0B
 70 59 2B 55 D5 23 32 3D 5C BC 93 7B CE 95 53 52
 F7 5A 73 09 40 23 6E 21 D4 9D 5C C6 D9 CA 3E F8
 C4 9F C3 E4 90 2D 8E 0F B8 03 B3 02 14 94 FA 9F
 10 CB 2A AD 30 75 E9 D8 81 B8 A8 58 A9 CA ED 55
 DC 0D 86 F1 8C 2A 00 E8 D5 9F B4 41 49 4C 29 C0
 3A 8E 06 F2 88 1F C5 0A 7A 79 B1 D0 E7 E7 4C 7F
 16 8A AD BD F9 F4 46 76 8D 65 3A FF CE 19 4A 4E
 B7 B3 F0 4E 1A E9 44 51 6D A8 7B 32 1B 79 BF 1D
 6F 60 F6 48 CC 87 7C 2F BB BE CB DA 13 8C DF 1D
 5B 49 C0 02 4E A5 CF 47 D1 8F 64 33 E6 89 86 5E
 17 8B 83 70 09 FE 0D B5 D3 06 C1 39 CD 6E 97 09
 1A CD 0F D7 87 6F 67 70 70 71 99 7F 2A 71 BD A0
 F6 28 F3 1E FA E4 3B 14 C3 EA 9D DE 39 34 87 8E
 B4 5F 15 F5 0E 30 C4 C5 23 95 AC 4A 4F 94 BC D7
 44 33 08 46 40 50 51 00 0B DA DB 6A A3 AE 01 C7
 D1 9B 0E F1 0C DF 91 2D 30 A7 3B E0 2D 0A 04 EC
 DB 20 70 48 63 61 6C E9 89 4E 82 63 A2 1B EB AD
 D6 94 6B CD A8 B0 50 74 DF 39 03 02 33 3D 04 AB
 D9 48 96 D5 F8 A7 4C 14 CD 13 8C B3 1B C5 95 29
 BA E0 5A 47 AA CF 67 17 39 93 6E 19 89 62 42 65
 B1 71 27 4D A9 98 51 44 C9 58 04 96 51 2F 90 97
 53 96 80 C6 22 07 82 97 34 83 6E 74 33 46 B7 61
 6C F0 59 92 37 09 0D E5 41 78 8D 6A 7D F1 0B A6
 C0 70 FE D5 22 5E 49 D3 78 AA 9D 3F 9A AD 33 D7
 83 36 F4 FF 09 ED 7F 16 61 1A 7A 4C 42 5B D3 3B
 D9 39 2F D0 CC 6A 56 3A 82 F6 42 23 F1 BF 86 6D
 F5 6D 51 B8 60 B3 1E BE 5E 89 1E 9E C1 43 F2 89
 E3 F2 5B DC AA 88 D7 84 1E B1 06 8A 97 F3 AD 2A
 51 5A 72 52 A0 5A 98 45 01 BA CF 7D AB BC E7 AF
 89 F3 DC 00 34 A1 DC 38 35 93 7B C5 20 3E 32 63
 0D B4 52 62 79 E8 F9 9D 00 B6 F2 99 FF D6 D2 35
 7D 18 12 3A C8 C9 C1 1B B5 DE E4 46 C0 4B 69 4D
 93 37 6F DB F7 47 14 F9 AA 91 C1 57 69 81 73 C6
 31 13 4D B2 F1 D7 68 C3 DA 02 53 A0 AB DE 3D 52
 18 54 70 A2 AD 9E 45 4A EC 15 96 E3 56 41 6C DC
 2D 98 73 05 76 BA AB 8F 2C 79 FA 62 8A 67 42 C9
 3E 18 E4 76 00 0B C9 ED 97 E1 B1 66 05 72 BF 70
 79 97 8D 79 03 A6 BA C6 39 5D AB 41 DE 0C E0 50
 A6 48 D8 3E F4 FC E2 B2 6D 4D 14 22 61 90 93 5E
 66 92 13 DF 03 41 36 07 1A 2C 5A C5 7A E7 C9 3D
 DC 7A 31 B1 2C 54 2E F7 83 58 59 46 BB 7E AC 56
 D9 31 77 61 68 A6 E5 27 B0 AE 60 72 43 F8 C9 37
 9C 5F 88 7D 49 DA 04 7C B0 EF E2 81 EB 8E DF 29
 41 7C 38 62 BB BC DE 36 00 59 E1 F4 90 90 95 6F
 E7 96 14 CD 6D 98 0A 07 DE AB 11 00 E7 A8 40 07
 3C 87 0F 20 84 C8 91 B9 84 BF D0 02 2A 70 5D 32
 C7 DF ED 03 A9 E0 64 11 67 09 5E 83 0B 11 E7 A2
 67 EC 3E A7 40 79 50 33 74 02 40 A3 5B 15 79 7C
 DC 19 DA 59 9B C1 7B 93 05 AE 97 E0 EE C9 A3 E7
 CD B9 51 04 5C D7 2E 83 4C 51 4F 18 9D 61 70 6A
 60 DD 8A 03 64 8B 76 36 AA 10 82 49 D1 20 DF 0D
 56 89 78 C6 9C EC BD 27 40 B7 3E 81 DE 3C 5B F2
 05 37 6B B7 5F 32 C4 16 82 40 75 B9 77 E2 BF FC
 65 18 4E 7B 68 86 6E 86 DD D0 69 1C 89 8E F9 5B
 99 64 56 D1 9C 41 F8 2D 14 60 4B E7 1D 13 8A E3
 AC 08 53 FD 29 F7 78 D5 5C 4D DC CD B5 9C 69 A5
 94 86 C7 C0 A9 F5 A1 2E 42 46 7F 0D 01 84 4B 16
 26 30 08 FA 62 6E 79 C5 73 17 D3 AA 3E 69 64 1E
 20 D1 A6 D9 18 D8 98 59 8E 3C B2 6A 3F 8F 3F 02
 8F 60 37 E5 68 57 48 D9 50 1B 2D 8A 46 C5 14 23
 65 11 05 32 9A CB E0 E0 BB 84 BA DE 29 94 2A 56
 63 87 EE 38 6F DD 20 B0 55 3B C0 2B B7 8D F5 B7
 1E F9 89 11 78 4E 0F 3C 1C 2F 9F AC 38 29 28 C6
 90 82 3D 08 8C F9 3B 07 0D B9 44 0E 84 1F 1D DE
 F1 40 2E 01 E6 BE 74 BF D6 5B 50 55 2B 3C F6 41
 C9 75 6C FF E3 93 0D 61 DC 7C 46 3B 95 6C 4B D7
 A8 AC F5 A1 C0 9B D3 6D 31 83 D2 02 F9 3C 93 53
 02 E0 68 53 19 D4 5B 8A 99 0B DE 86 89 78 29 AD
 6F 34 F1 59 9F C0 A1 47 0D BA D5 2B 5B 1C F7 E7
 CD 3A F7 F7 F7 EE EB DF E4 9E 5C 0C AA 1F 9F 94
 76 4C 3E 15 A4 50 46 38 B8 F4 AC A1 AD 8C AE 45
 66 2D 2E F1 0A EA 22 12 9F A4 34 2E 43 1C BB 5B
 AC 0C F6 5D C7 5A 9C EC BF D8 38 C4 D2 3B 78 6F
 1B 4C B7 35 47 91 51 7A E8 7F CF 68 24 4B 24 47
 D0 D9 82 A6 B1 82 58 BE 69 88 D4 DA E9 33 7E BC
 92 B1 78 78 68 21 C7 11 EB 18 F2 2E 8E 24 C4 95
 53 9E 42 3D C8 51 40 D4 04 B0 27 98 BD A1 92 EE
 16 A2 B1 AE A3 20 B6 7B C2 A0 29 F0 77 39 6D 96
 F9 F4 99 F2 D2 24 EB C7 B7 1D C2 82 DC B9 E2 E0
 3D 85 BF 56 2A D5 64 18 CB 67 D5 F4 B8 A3 51 81
 8B DA 71 50 16 7A 51 72 AE AF 38 08 3C F9 46 88
 4C FB E4 84 18 33 DC 26 5A EF 63 0E 8C C8 AC 3C
 BF 88 D7 50 B2 5C A6 56 42 66 09 44 1D CD FF 45
 CE 11 71 32 24 1E DB AD CA A4 16 9D 4D 68 16 67
 9D 58 91 B6 C2 37 AA FF B9 A7 6F 94 AA DA 3A B4
 B9 57 BC 98 B0 B8 84 D5 71 BE 00 01 54 B4 55 FD
 83 74 86 F0 9F C6 87 0D 4D FD 15 6E 52 EF B0 BD
 5A 11 65 05 6A 1A F6 AC E0 D5 02 86 EA 11 95 C9
 E6 F9 50 C6 72 50 54 7A 51 D9 B4 0B 2A D0 62 29
 FC CC 26 60 FF F2 F9 41 14 55 62 CA 77 65 76 CE
 33 7A C1 23 34 C2 97 9E 8F 89 BE 58 DA 60 F5 CE
 4D 22 F3 6F B4 62 EF D2 16 92 8A F3 BD 2A 41 A1
 E7 10 24 BE B8 40 C5 F4 76 2A 91 99 47 BB 41 95
 66 F5 92 81 94 20 F4 CC BA 80 AA FB 11 68 26 A1
 29 BF A7 B0 96 B6 D0 FC C4 59 0F 3F 0F 50 8A F9
 05 73 2A 73 56 48 87 3E 02 28 0B 36 5C A6 7B 29
 83 DB 98 71 B7 ED 7E 46 18 10 90 F6 7F EC E1 0A
 BF 2E E5 58 CF 6B 80 2F 99 B5 AC 81 49 75 45 FD
 DF 7F 69 DB 86 9A 87 36 E4 0B 4F B0 9E 79 F0 A9
 9C 72 14 C9 68 06 75 A3 C6 17 65 E4 42 C2 2E B6
 A6 90 5B 58 BE 58 2E 26 F0 7A F8 38 F2 33 99 90
 59 ED 67 96 9B FF 64 E3 06 F0 1C 28 E0 9F AC B9
 C5 48 EF 03 6F C5 49 93 25 7B AD 31 0A 3E 4F D8
 60 74 CB 72 9C 31 AE 96 A8 77 19 D1 D4 15 39 94
 52 3F B6 58 6F 77 25 B3 C0 11 79 A1 95 5A A2 C9
 A8 C2 90 D3 0A 89 31 B5 46 E5 0F D8 65 D1 AE B5
 96 2C AD B7 CE C3 E5 17 8F 9A 77 08 6B EC 0A 65
 E9 E5 BC 15 AC BB D3 2C DD FE B9 28 FE D0 83 60
 41 CE 02 49 EA 0E 4F 04 66 DA 61 66 37 2A EB FF
 AB 88 CA D8 97 DF CD 1B 29 06 09 8E A3 0C 4A 62
 7D 5B 1C CC D2 26 B9 F4 95 49 F1 F3 FC C3 C4 16
 4B C0 44 8D C2 A8 0C 29 4B 7B D6 BE 79 12 C0 D4
 5E E9 1A E1 31 1F AF 1B 0A 16 95 0F 13 92 CB 46
 91 E5 43 85 0F E2 17 40 D8 51 B1 8B 94 31 7D 98
 EC BD 39 36 4C 7B 0E 10 3D E8 73 50 10 72 18 2E
 FC 0D 53 C2 E4 6E 2A EE 09 41 3F CD 75 05 40 B7
 C1 84 34 B6 F0 C0 16 E5 5D 23 AE 25 24 7A C1 8F
 30 1B D5 17 4D 19 1A 8E E5 23 CE 34 A6 9E B7 23
 36 59 B1 A2 32 C7 6F 4C 9C BE 19 A8 30 90 A5 FA
 DF C9 17 0B 24 06 46 3E 26 1F 14 00 35 C8 6F 9A
 43 3F 5B 25 AF 56 D1 80 1D 9C D1 E5 A6 D5 95 E6
 58 97 36 4E F8 E5 CD 83 5D A8 E2 C1 60 93 CF 48
 C8 76 99 05 E7 DD 8D 2C DE 61 DC 1F 5B B4 72 7E
 8B 80 79 08 B5 8A A4 ED 9D 99 3C 86 C6 05 18 9F
 58 7E 04 54 B4 05 F3 F6 4C 3E 7A 70 16 82 C7 58
 43 95 9C EE 8A 05 A4 AD 40 6B 90 D3 78 E2 C3 99
 85 EA 35 53 4F A0 59 9F E5 F1 4E F2 A7 69 CD BF
 FF C0 B6 44 C0 9B 13 75 FF BE 76 DA C6 81 BF 32
 00 9E B8 DD 4C 92 45 70 73 EA 8A 7B E1 CD 3C 4F
 66 0D 54 94 34 99 30 1A 29 5F EE 2D 17 74 83 E6
 87 2D CB 5B B5 86 90 3B 4C 83 03 C5 CD DE 82 11
 E4 C2 98 63 F1 CB B1 35 B3 3D F2 4B E6 1A 50 1E
 9A D1 D0 13 46 76 78 2D 99 65 EB 22 FC 75 05 62
 9F 65 FD 1F CF 05 3D 50 13 F4 91 09 A8 45 2E 41
 99 38 CD C7 3A 42 6A 94 85 BB A9 90 F5 AB E2 AD
 D0 77 59 2B 61 9D 41 7A F6 83 B9 0F 64 D9 DE 48
 6E ED 01 24 76 45 41 49 CA FD F3 F8 DA 87 8E 5F
 F9 73 A1 F6 CA 85 51 14 67 3E 64 F4 6B AA C5 A0
 2E 7D 39 26 53 FD 2A D3 82 34 35 3A 13 9C 6C 10
 AC 39 24 E7 F6 0C D1 97 72 EE 2D F2 24 DF F1 59
 D1 A1 AF 18 F5 9F 81 8F BC 90 0C 08 FA 6F B9 56
 98 AC B9 ED FF 41 5B F2 F6 0B 62 C5 1E B1 0E 8F
 4E 31 F5 F4 E8 D4 4A 89 F5 6E 43 52 AF BD 00 50
 83 C0 5F 31 45 07 90 B0 CA F6 40 97 07 DB D7 D7
 49 2D 1C 96 E4 D8 FA 8F D5 3E 7B 7B CA 79 25 0E
 D4 9D D2 5D 66 93 FE 11 54 6B F7 10 63 BC AC 4D
 19 DD FA 12 37 B1 81 65 F4 39 D5 B4 43 2C 14 90
 B7 F7 B4 BD 50 CB 40 35 2C A4 57 DC DC A6 F2 D5
 1A 88 47 AE 1B E9 CC 8A C4 25 8E 62 CF 9E 2D 4A
 55 C1 9E 41 5F A5 F8 31 A0 BA BA 6C 60 C1 79 E3
 43 F8 E1 0D 67 B7 1C E4 23 46 63 6D BD C5 56 4D
 98 DE F7 CB 51 1F 84 75 F3 E0 1B 83 3B 84 3B 09
 35 7D 29 6F E5 96 26 F8 9D 1D D8 7D F7 F8 47 03
 F2 C5 55 11 72 43 79 91 C3 03 FE 92 B1 96 FD 79
 05 9F 5B 04 10 18 6B 8A A0 10 A9 98 6E F3 5F 6A
 88 30 25 58 E5 5B 5A 83 F7 6E 64 B0 47 5A BD 7C
 15 71 A6 8E 41 85 D2 14 36 B1 40 5C 99 4D 61 C6
 B6 91 4A 29 FE 2D 6E 14 52 30 6B 94 80 F8 C6 A1
 F8 16 EC C5 E5 EB 3E DC 01 DC 55 75 02 D6 58 DF
 B7 9B 3B 21 22 C3 C9 E5 FD 34 5E 10 4F 35 18 FC
 73 F7 D7 2E B5 56 96 E8 40 A7 43 01 D0 7E 46 35
 93 F4 91 D1 00 44 28 AF AE 31 AB BF 9C 61 31 EF
 A7 F4 B7 DF B8 54 A2 39 70 C5 C9 B2 A9 5F 22 49
 7A A4 F7 7E FB 2A B5 B8 AA E7 E3 3A 8A E7 6E 30
 79 4A 2F 50 50 F7 B8 A3 D4 0B 37 A2 17 F9 3C E4
 94 F5 86 83 28 6B 0F CC 62 84 42 22 BB C5 2D 54
 11 D3 25 D4 72 6B BB B5 2E C3 4A 20 6A 62 82 65
 96 7F 2D 0D 51 89 24 1C 85 68 1D 84 93 8D 96 E8
 F0 5C C0 E1 6A 69 87 DE 45 8D 32 F0 E5 21 37 C1
 62 D5 A0 A0 E1 89 B5 2B E0 32 F7 53 AE 04 0A AB
 81 2C 9D 8D B9 84 5D B3 C2 70 20 0E 1B C7 48 E3
 EF E0 CA E1 47 7D 34 4D 78 2C 25 98 1A 75 D2 34
 74 88 28 01 D3 78 BA 38 47 77 9C 77 BE 7A 73 C8
 30 F5 EE BF 75 C2 99 24 ED 3C 52 A1 5D 44 17 47
 82 77 C5 06 EF 00 C9 CE 49 B6 94 5C 80 03 BA 0E
 A4 D5 2E BC 29 04 2C 0B B0 17 46 B5 DE DD BF 1F
 A4 37 EE 87 13 C6 07 AF 88 63 B1 77 9B 69 FB 37
 06 56 F2 CF C7 11 6C B2 3F C4 28 38 2C D1 A7 8C
 04 95 2B 62 EF 7D 63 4B C2 E8 4B C8 08 4D 6D F4
 F8 5B 63 BD 51 B5 EF 58 6E BC 21 60 E6 29 E3 21
 5D 0C 8B D3 9E C3 11 6F 06 00 0D 9E D5 49 9F C4
 21 4C 2B 09 80 F2 7E 08 CD 46 AE 8A C9 95 79 16
 6D 79 E5 82 DB 5C 46 EF FA 82 CC 80 A7 C6 81 06
 AA E6 F0 03 E4 26 53 C7 DF B6 48 E4 F5 D5 11 D3
 53 1D 4B F0 65 8D 79 B1 F8 5D E7 84 F6 4F 74 15
 FF B4 9A F9 00 AB 84 0F 1C 5E F6 C6 71 AF 03 7B
 7F 4C FE F4 BC 26 6A C1 76 07 36 FC EB 27 76 12
 7F CB B8 58 28 99 04 9F 3E 5A 83 BC 84 A8 83 FD
 AB D3 87 13 52 67 9E A3 C0 B5 A4 AE 6C 95 67 AB
 03 7E C5 3C BA D5 44 89 D4 E0 AA AF 55 C1 B0 59
 E5 EC B8 FD 8F 5E 36 98 3D 94 07 06 94 99 FD 86
 1D FE BF AA 17 0D 2D 0A EA 69 81 6B EF 3A C6 1D
 D1 82 3F 34 A4 E5 D4 E3 F7 CF AA 30 B1 A2 02 F7
 69 64 16 DD E5 D2 11 E6 1F BA CE 60 AD 31 07 CB
 B3 74 39 F6 BF 18 57 A8 5B D5 55 DB 60 35 6B CA
 AB 04 DA CC C4 26 6D 55 18 D3 D4 9A C9 16 4C 70
 0D 35 DD 06 D6 34 31 07 71 EE 65 B7 6E 0C 81 C5
 0F 5A A6 67 AD B7 F9 60 9F 9A FD E4 A4 B7 AE 94
 A8 2D D6 47 93 36 E5 70 FB 56 48 17 2A A7 58 A1
 F9 47 E0 31 D2 25 04 CD 00 50 C0 D0 8D 4A A8 9C
 60 DC 73 BC FD 72 B4 52 61 CC 9A E4 7C 71 A2 ED
 7A 47 A3 DF B3 4F F7 B4 09 07 CD 0B 6B 15 F7 60
 23 6B BF CF 16 D6 07 DF ED 43 4F 80 C0 D8 21 CB
 C3 F3 28 C3 7F 89 94 B4 12 BA 27 6F 80 44 9F 2A
 F7 78 E7 C3 1A 13 1A F2 AF AC 70 F4 8D C9 BC D0
 BA FC 3A 92 52 4B ED B6 6B C9 0D FE 9E 45 44 40
 9A A2 02 C3 51 A4 C7 CE 17 11 8D FE 61 07 04 D1
 E4 D5 3E 28 E7 42 2E 75 DC 23 F3 80 D5 2F 63 5F
 A9 6E BC FB A9 34 EC 1B 05 C9 82 5B 0D 17 3D 2C
 25 0D 28 BE 1B FC 7F 10 ED 53 A6 A8 D0 5E 0E F4
 C8 37 6E C2 53 25 92 15 16 96 62 18 74 6A 34 7B
 DB 32 1E 07 3E 63 DF F1 2D B4 A4 EF 21 C0 C6 6C
 0B 0B 6A 8C FD 73 C7 47 55 27 FD 2E 6E C1 09 C3
 5F 15 AD B0 DB 7B D4 04 DD D5 21 FB A2 73 74 A6
 16 26 37 68 46 33 25 E7 9D 7B A9 E4 71 7B AB 95
 9D 3D 29 A5 C9 44 5C F4 18 7A 45 3D FE 9D 00 D6
 0A D1 FA DE D6 31 1E 97 69 B3 19 C1 C3 79 AE 92
 CA D9 B6 25 63 8A D1 6B 39 71 DF 52 50 20 04 9A
 16 3A 34 D8 B6 98 CC 4A 86 4B F8 EF 02 DE 32 AA
 7F E4 5A 98 18 DE F4 97 C1 B1 E0 0B B6 B3 30 81
 0F 5B 9A 31 82 27 99 02 A7 DC 85 0F 2A A6 C1 2A
 FA 94 5D ED 3C 93 F2 08 96 48 8A B0 AF 54 40 94
 B0 BD F8 F6 31 87 D1 61 A5 3E 55 72 0A A7 AD C1
 49 F8 B7 DA 79 FA 25 ED 51 73 37 87 A5 5D A9 9F
 72 3B 19 82 3D 12 05 05 47 CD E3 4D D6 37 41 E9
 F6 08 C4 60 5B 34 09 40 F4 6F 7D C7 CB D3 2F 94
 CE 97 64 55 9F 8C 61 E0 A8 21 CC 33 A6 1E 6A 1E
 FE 58 C7 20 32 E4 8E 04 B0 C0 C7 32 D6 7D 0B 1E
 A4 87 55 77 02 E6 61 E7 24 F0 89 5F 48 8C 93 85
 3E DF 05 7D 63 4C A9 41 1C 5C 2F BF 1F FE 2C 85
 5C 29 86 96 DC 4E 7C FE F3 40 A6 AC 5B 28 18 DE
 14 8D 31 35 1F A4 18 AC 61 1B 9F B3 99 6E 05 96
 D0 D4 52 2E 1A F8 EE E9 9F 55 3E 0D 20 D1 E4 D3
 19 F6 BE 9D A7 10 AC 2F EF CE 45 7E AC EB EF 1B
 33 32 03 B8 E7 DF 84 BC 53 CF F9 BB 4F 74 0E 63
 B0 21 57 37 61 33 26 01 68 1D C6 74 EB 3E 03 DC
 F0 4F F3 AB 15 4E 10 9F 22 C5 53 DA 2C 3F BD AA
 CB D6 79 90 29 5E AD E8 67 73 1F 23 E5 CC 41 DA
 93 64 19 01 7D 31 2A 52 3B C9 65 D1 4F CB 0D 34
 C1 A5 38 FA 79 88 7A 79 72 2F 1E C9 A0 0F 34 10
 4F 80 B8 5E 79 26 B6 1E C4 7B A6 C2 71 E5 B4 57
 66 39 61 A3 58 B7 AE A4 5D 5B CA FE 72 16 51 A4
 97 FD FF 3D 85 E9 A0 40 DF D0 E1 8F 19 C0 AB BC
 88 74 AD 9D 16 59 6C 5A 56 2F 1B 51 DC 6A 6F FF
 6F 63 F6 2D DA 9D 75 EB 55 F3 76 D9 78 6E 1E 25
 C3 B4 2E FA 45 78 4E 4E BA 69 84 AF BD 5E ED 4A
 BA AC AE 4A 73 6B 67 C8 D8 36 5D 68 B5 5F 42 FF
 5A D3 12 77 A7 5A 74 BB C6 BE 2E 65 56 8F 16 C9
 00 26 F9 76 9B 4C B7 6D 3B 01 34 F5 5C 06 C7 F7
 6C C9 2B B4 C3 D2 91 52 E9 AD EA B2 41 C6 09 1E
 E3 A6 85 FC 84 CC 48 55 34 45 18 C0 BC E2 B8 2B
 DA 33 B8 54 E2 1E CE 14 55 DC 05 BD 1D 1A 5C DA
 4D 90 BB 1E 40 FF 1C B7 F5 66 A0 27 C7 7F 4A DD
 E2 95 1C 64 12 34 54 95 90 A7 29 FD 25 B2 C0 F2
 EE 6E 04 D1 56 22 FB 16 51 4C 79 BB 2A 46 D9 0C
 8C 15 7E 6B 5F 14 48 70 ED FF BB B0 2D 4B DF E2
 CB 4D D1 BA 19 99 86 5D 5A 2C 43 DE 15 A8 9A 2C
 43 DB D4 2E DB 95 7E 83 EE 8A 3E 28 9C A8 54 50
 50 DB 21 93 FF 14 FD 78 8E 1F D0 B3 D2 F6 85 E8
 2F D9 9C BB 0F 55 71 50 28 4F B5 E4 9D 14 2B C9
 33 F8 0A 55 4E 3B 96 98 A5 C4 4F 93 82 D3 B5 AE
 EC 5C 7B D3 74 06 AD CA 6F 1A E8 9C 0F E5 3B 49
 FC 8E 9C 32 89 7B 92 DB CC AF 7C 3F 72 CE DC DF
 A4 B1 C7 89 C7 89 C1 20 31 BD 0B B7 44 FC 6A C4
 E8 FD C4 03 67 3B 9E 61 37 34 71 A5 03 29 7D AA
 F2 CC 53 34 A3 78 A4 B6 AC 38 0A AE 4A 40 A2 1A
 25 FA EB 93 05 72 83 26 8A A7 5E EB 6B C5 5A D1
 05 81 EF 67 7B 39 A1 04 AA 85 00 06 7E 87 F8 4F
 22 47 2B 3A 49 78 34 EF 80 AD 8A FF E5 B7 39 4D
 31 A0 19 9D F2 42 DD 5A 24 C0 09 A1 EF 08 CE 26
 5B 95 D7 86 BF 87 14 6F 21 1E E9 5B 0F 22 DF B9
 8D B0 86 FA A4 68 B0 19 63 27 63 24 3E 6D 27 0A
 1C 92 42 60 44 86 7B 3D C3 E6 11 AC 1A 84 6F 84
 5B 59 65 32 E8 C4 55 39 5F 27 F5 6C 14 92 7C 17
 95 6B D0 07 A0 70 95 49 9B 04 AE 21 C9 5C 4C 7D
 07 C0 38 95 F2 92 89 26 AE 18 E4 56 E3 C9 48 69
 FA 90 CD 65 90 F1 DE 33 B3 EB 6F 70 11 73 4D 76
 89 3F 84 26 59 F0 FD 8F 38 4F 89 E0 EE 58 87 44
 FB A1 70 45 4B 10 C8 3F 6D 36 85 DE C5 18 34 98
 0B A7 07 AC A9 9E D3 E3 3A 7A AA B5 0F 89 F9 E4
 77 8C B4 C3 56 2F B9 CA BA 9C 12 B5 C3 41 51 E9
 20 F5 02 8F 5D 07 AE 15 00 C3 87 20 17 21 40 07
 25 34 BE AA A3 6A 93 74 AA BE E8 8B AC 13 CF 1A
 D7 F8 37 0F F7 06 FB 89 B6 79 43 B2 7C 2C FB 72
 51 D1 52 B9 4B 2D C2 5F 6C FF 8A 0A 0D 86 1E A9
 A5 D2 DF D1 7E 4A F0 DC 70 2B 58 4C FB 59 23 2B
 3C 28 8E 6A 08 0B 60 35 16 E7 AE 27 FD 4A EB FA
 18 55 28 EA D0 4B 55 9C EC 25 7A A0 EC 4A 70 F5
 73 48 99 4B F0 1D 1D CD EA 97 C1 1A 74 AE 94 D8
 E0 5E C0 8F F2 A8 08 11 36 BD E3 A4 73 F7 7A BF
 25 CB C8 36 B1 5F 29 19 6B 79 07 BA D5 41 B9 F2
 7A 53 F6 8D 45 24 C5 7B 6F 77 68 CF CE DE 90 F1
 EA 7E 81 16 FD D8 EF 28 AC 0D EB 1A EF DF 04 47
 1C EA C2 56 3C C8 F6 13 B7 1D 9A 74 AF AD 6A 8E
 9B 6F 38 46 1C DA 2B B3 27 01 2D 72 C7 18 BC B5
 BA 1B 9D DA D6 3B E9 7A AA 8A D7 91 5E 40 39 FF
 61 CE F3 F5 C1 38 2E 08 F0 1A 9B BD C6 0C 20 8A
 DA 9B 32 FA E0 1C C8 D2 9D 13 56 93 D5 99 61 9D
 91 6F 30 B3 86 47 9E 36 1D C4 4A F4 12 75 F2 5A
 8A 68 EE B6 1F DD 6A 8B 11 17 31 7F 0E 26 E5 4B
 6E 08 D8 99 09 DB F0 8D 5F 1D 0C C1 B5 F1 4C 9B
 BC 8D F7 DD 80 99 5D DE A3 88 EC C4 CF CE 5F 71
 F6 86 61 9C 29 AB F8 4F 22 B6 0A D8 24 D4 F1 A9
 CB 38 AD 67 84 69 F2 A0 08 16 1D 14 C4 FC 47 37
 4E C4 8F C4 AD 4E 98 BB 80 62 ED 47 D7 41 49 3A
 13 8F 36 4E 54 06 AD D9 5F AF F5 54 14 BD 50 EB
 20 A9 35 05 69 61 4A 88 6E DF 8E 91 0C 1D 3B 1D
 04 BF 1C 80 39 E9 CA 4B 75 B9 F1 3B 18 4C 5B 9D
 15 1E 4C CA CE 22 5D 36 D1 12 C4 E3 39 41 A4 95
 16 1B D1 0C 92 EB B5 EB 71 E5 AE 96 F7 DA 03 11
 4A 83 52 A1 D7 C5 F8 6B 44 73 8C 22 7B 21 CD 97
 CB D4 94 C5 9E 26 8F 24 4B AB CC 19 E6 49 E1 DE
 D2 FB FE 74 2E 26 15 96 B4 9B E4 B4 F3 A4 BD 2D
 EA 8B A8 CC B9 9A 4C 2B 71 AA 84 D0 C9 15 CD 8B
 60 E6 1F A6 CA DD 19 15 28 C4 5A 36 8A 61 11 5B
 CC 8E 7E D9 EE 40 03 29 18 AC 51 EB 1B A9 81 2E
 4C E6 44 C1 8A 4E 12 EC 33 C7 AA 70 42 C2 DA FC
 18 5A 9C AE 50 13 C3 82 04 AB A7 05 5B 81 72 1F
 42 D9 E6 28 BB 37 83 3C 3E 16 94 9A 01 6C 4E F5
 3B 91 3D DD 65 ED 00 19 DD 4A 46 E8 BA C5 8C 84
 C2 C8 0C 36 4E 1F F7 EF 1F E9 AE BB CE 6E A3 01
 8B AB BE B7 0E 21 FC 78 94 7D D0 1A 08 A6 0F 76
 50 26 32 2C 7A 60 C3 3E FA 90 4E 31 DE 06 9F B7
 05 D2 FD 90 50 63 68 61 73 BD 42 AC 3B 2E 97 8B
 FB DF E7 40 16 D7 39 81 0A B4 A1 A3 C6 CC A8 A0
 E9 99 10 0B 3A 70 5C 06 31 AB 3B 87 E6 1D F1 D3
 05 A1 65 1D F9 57 44 00 2D BA A4 7A D8 DC 72 94
 19 25 9F A7 F3 E0 46 3F F7 91 65 26 5B 99 37 11
 9D 74 CC 32 23 43 BB 05 69 84 18 C1 4C 54 C9 19
 94 63 FE 7C E2 BD 34 B5 7A B7 C4 98 90 0C C6 3A
 A7 6C A4 B7 DA 7D 81 77 C0 1F E4 26 C9 FD 8A 47
 6F 3A 54 6C BA A3 28 D6 5F 57 21 AC E6 C7 C4 7A
 AF ED 90 BC BB D0 DA A2 D4 7C EC 5C 9C 37 0B 9B
 7F 1A 30 AA AE 3A 9A D0 A4 5F 9D F4 51 77 B6 93
 11 AF 9F B3 5A 4C 62 E5 BC B1 EB B5 BB 02 CF 3D
 9A B2 CC 66 C7 3B 5A 2A FF B5 65 E5 65 DF C0 69
 D2 13 E2 17 EB 83 39 89 14 C8 9D 95 E2 76 EA 60
 F0 0D 46 B5 89 14 98 B9 7C 79 C5 89 47 14 FD A7
 76 B0 02 C8 D4 45 D0 00 93 85 1B 4F A8 C6 35 3D
 99 6A E1 B7 EA 2C C7 76 1D C8 B6 50 A2 9A 4A 11
 3D 65 01 C6 2E DB C2 AB 34 88 CE AD 82 DB 67 08
 2B 89 A5 E7 EE 7A F6 65 29 50 E6 33 C8 B9 42 AD
 D2 5B EE D3 7F 86 81 EA 5D 52 CC 2F 63 9C 83 AA
 39 9A 2D 6A 64 D8 C4 8D 41 2F BE FF A5 BC 5C CC
 0A 0B 46 F6 A5 41 EE D5 AD A7 25 85 88 AE AF A1
 5C C3 0E 74 E5 B0 A3 9F 88 BD 04 5E 77 9A 10 8B
 1C 36 24 BC E8 44 CB 53 50 A9 6C 36 87 C6 1F 22
 CA 02 CE C5 C1 2F B4 6B 9C 21 E4 6E 1E 40 7B 67
 8A 26 AA 9D 50 07 D6 7A 41 58 6D 32 7F C1 A6 65
 4E A0 5D AC 10 39 3F DB 97 B7 4B 98 05 D8 58 3C
 5D 17 E6 99 B3 74 81 5A DC 12 44 C5 95 BE B8 97
 08 6E 72 8D 28 22 07 B2 03 C5 A0 AA 7C B2 78 8C
 81 0B F5 06 4B 90 F8 D4 08 2F 61 7D 24 ED E2 BF
 D6 28 92 72 A9 74 E4 4B 09 5F DB 3A 54 CF 4D A6
 14 BD 5F FE B4 54 C9 67 7D 6E A9 53 61 36 FA 0A
 8A 45 3B 6C ED A2 55 1B 96 72 AE 80 6C AC 54 FD
 9E DF 88 8C 10 6B 36 20 81 DB F0 51 31 24 7D DF
 AE 75 AE 7B 7E BD 19 E2 1A B5 D7 11 7B 1B 92 B6
 ED 78 5C ED DE B7 89 17 CD E6 64 6C 28 20 C4 7E
 5A 75 59 A7 01 B3 FE B6 C2 11 28 D5 AA 87 3E 6F
 8B 17 20 5F DA 10 11 1E 0B 5D F1 71 7C F6 86 0F
 05 70 A4 2E 2A C9 E0 AB 11 49 5F 64 6A 39 39 A6
 B2 EF 62 29 1D 54 4E E7 5B 10 51 A4 85 EC D2 42
 AD 69 AB 4C 72 55 8B 0F 14 6A 2C 0A 7C 42 7D 5A
 5A C7 F0 1E BD 6B 5C 13 EB D9 E0 B9 D7 B6 F9 A3
 A5 20 A8 F7 21 22 18 AA 39 7F 7E 0E E9 A1 7B E5
 F0 16 7B 74 0E 42 6D 5B 3F 89 CE BD EE 99 D1 B6
 8C 83 FC B6 D3 3E F2 D4 43 98 EC BD D1 60 A9 1E
 67 54 BE 03 0C 22 AF C9 80 33 5A 2C 81 7C 6F 4D
 2B BE F7 DF 4B 30 B4 B7 0D 67 BD 14 5E 36 6D 7D
 35 AE 04 AB 15 80 55 FC 8B 4D F7 23 72 01 BD 10
 29 8F 2F 33 48 D3 4B B7 66 9D F6 02 CB D2 7F DE
 85 1E DA 40 F8 5B 17 1E EA A0 33 9A 00 83 A0 21
 3F CB 63 80 9B 43 D3 F2 80 1D B9 9D 43 09 B5 C4
 F4 29 E3 2A DC 63 86 8D F2 EE 04 6C 11 69 02 43
 3B 92 DF 53 84 78 7A 92 72 64 54 55 AA BD F6 34
 7C 4D CD 6B 8C A4 C3 8A 50 DF 67 E4 8B D1 24 3C
 E0 75 78 42 82 4E 54 3D BA 8D F4 16 D5 BB 73 26
 2B AB 66 53 B2 13 42 62 99 98 EF 52 D3 A2 A1 B7
 98 EB 49 7C 05 37 48 3C F2 3D 61 DE 07 15 CA E1
 E4 EF 87 5D 32 A3 20 DF 3B 55 72 42 3D 14 5D FB
 AC C3 3D FA AA A8 D8 A1 CC C1 DA 97 78 AB 0A 37
 14 D4 C6 87 4C 5A E3 0E 0B 41 B1 66 A2 AC ED 89
 7D 23 FA C7 1B 94 13 E3 59 4F BB 52 C2 30 DA A8
 8A 2E 70 D8 05 B0 15 08 8B 69 3F 09 9E DE 87 47
 68 A3 C7 FF 4C 70 CB 6C DA 79 9B 4B 69 D5 05 18
 67 9A FD 1F 39 AA 34 EE D3 69 91 BC 65 58 FB 31
 5E 9F 10 00 84 DF 97 AD 23 D5 00 EC 69 7B 0C 8A
 14 19 EE 46 25 06 0D D7 94 04 6E 93 35 B8 22 F5
 06 2E 56 AF 63 8F F0 20 F0 A5 BB 0E BD FB 2B EF
 57 97 74 6C 2B 9B DD 95 01 89 12 06 69 61 44 B9
 86 89 B4 ED 1D CB 6C FA A6 5C E4 F7 F9 72 E4 BC
 BB BC 5A B0 7A 5B 1D 2A EB 49 F4 56 FE 47 4E 88
 4F BE B3 A2 4E FC 92 58 34 34 AA CD D1 3C 7E 33
 F1 CF EC 4D FD 07 18 59 AB 35 4E CB 92 39 23 64
 74 AF 72 04 39 D3 49 A6 7C C6 4B 8E AD 74 A6 50
 CC 64 EA 29 DB E8 9E B8 EF C4 2E 43 0F 2C 38 0C
 7B AF ED E1 D1 12 6A 4F 4A 09 8A F6 81 62 C9 4D
 DA A3 45 0D 8E A4 97 70 83 10 30 48 58 34 51 33
 60 C7 3A 0A 19 73 11 34 06 B3 CC 7B 87 C7 E6 5B
 3E 70 71 3B 5B 98 A7 F8 8D 4F C5 E2 CF 7B 1D CF
 A8 4D FC 64 3D 0B AB 1A AB 98 F1 A2 8B 89 24 FC
 EE 5D 1E AF 5E 96 B9 D2 F6 48 F3 5A 42 F0 59 F9
 DE 18 AF 84 F9 88 AC 76 72 64 52 6A 6F 19 D1 5C
 45 37 E2 CF 44 B7 83 07 0F DA 30 E1 AB 36 18 54
 A2 2F D8 BE 5D 84 9D B4 51 77 1B A2 E8 27 C5 FF
 F7 AC B9 74 B6 3A 78 8E 57 CC B7 7C 5A 7E 9A 73
 AA BC C3 8E 68 89 88 6F FE F2 1B 29 85 0E 30 8C
 40 DB DE 0E EF 6C F6 8D 0E 60 43 D9 67 73 68 BE
 19 FE 3C 94 EC D8 1F FC A4 C6 96 81 68 A9 93 66
 50 0F 7A DB 8F A0 4E 06 75 0B 4F AA 61 3D B1 70
 8A EC 12 E3 B1 EA 9D D8 56 14 94 22 CC 41 F6 69
 DE A7 74 EE 29 06 7F 44 CC 83 BF A2 58 20 FF E8
 20 15 1C 2E BD B8 78 89 59 11 C4 81 C7 3B B5 23
 A4 31 34 7A F6 7E D7 DB F3 FF 8D C6 61 5A FF 65
 27 8F 3D 36 AE C0 89 48 18 5D F9 A1 84 A9 AE 5B
 1B 63 01 36 A1 B0 B8 5B 3A 3F BE 49 89 F4 66 9D
 88 35 A7 89 99 84 4A 54 73 26 CE 30 B7 40 5E 5B
 6D 39 52 69 65 D5 22 7E 3A 73 D7 2A 46 2F D6 9D
 A2 1C 33 48 8D 06 CD 89 9B 51 F8 A2 D6 58 3F 3E
 1B 72 47 E0 5E 78 23 28 6D D1 0D A1 D9 18 70 93
 60 4B D4 45 0B 18 5E 50 18 5A 91 69 F3 F4 8A 28
 16 EE B3 16 B5 3C B4 89 51 76 88 26 E0 35 B9 C5
 10 BF 4B 29 C6 B5 7A A8 84 CB FF DA FB 23 15 BC
 D9 A6 F2 0E E5 9C 68 43 18 96 A0 1F EB A9 C3 AC
 11 C9 3C 33 5D A1 65 48 91 B8 E1 12 E0 6A 79 EE
 83 7E E1 97 BB 60 ED 7C EE AC 67 11 3A 58 83 E5
 FF 6A 74 D4 26 E7 9E 2E F5 55 B4 FA 99 1C 4F E6
 A6 90 A5 34 C2 CE 4B C4 F0 7D C0 68 B3 91 1E D2
 61 97 21 68 55 48 96 39 31 49 F0 FF 25 2D 41 E4
 6E AF 04 6A DB 5A 64 D8 A1 59 01 F9 1B E0 35 53
 00 EC F2 64 D1 E5 62 2A 68 80 A3 9B 9C 6C 8D 7C
 68 77 5D 95 E8 C9 A8 4C CF 4D 22 65 DA 04 17 43
 E3 60 67 1D 11 13 97 8D 5E 61 28 CA C3 E8 83 1E
 8C 57 47 1A 85 B2 23 47 6A 84 DE 65 5F E6 69 2B
 3D 86 56 26 3A 75 69 A6 AC 92 8E 15 A9 32 0B F5
 DF 8B 7C 09 CD D5 1F 3F A7 FA 3C E6 75 DB A6 42
 38 F6 A3 53 A5 CD 4E 11 81 56 7E F2 96 47 76 5A
 F5 6B 03 EA 10 1C 70 E4 C5 F0 63 51 35 5B FA 56
 ED A5 05 44 6A A0 A1 39 E0 3B EA D8 7E 9D DA 40
 25 E7 AA 19 5A BC D2 AE E6 13 F3 FE 0E 94 43 59
 D7 DF BB 87 5B 98 32 1F E8 52 19 60 AC 62 BF 19
 E8 1B 51 AF 03 48 2A 94 A5 4C 1D 23 DE 16 97 26
 D9 4E 82 82 53 89 72 2A 65 D8 35 69 A2 D2 01 8C
 A5 E7 FA 09 D5 ED 8D ED 66 38 3D 72 F1 CA 66 C9
 E1 67 E8 76 F0 CD F7 6C E3 6F 69 31 A7 93 74 A5
 3E 1E 27 D0 C7 C5 7F A3 EA C0 41 9F 60 5A 3E 93
 99 8F 1B 1E 49 AD A9 6C E0 43 FD 2C FE DA 5B 24
 9C FD E0 21 B3 E3 70 CD EF 73 51 0B FA C8 A7 7C
 D9 CC AD 3A AA 1B B0 75 C5 DF 11 C9 14 9D 69 08
 8D 4D EE 0C AF 9B 1D 4A CA DF CA 00 49 75 E6 F6
 18 65 F1 26 58 52 D4 29 2E A3 26 61 86 08 3E 7B
 AB 96 E3 38 21 C8 25 7E 53 23 4B CC A3 EB 34 AC
 21 39 7D 06 96 31 F1 25 9B EB AA B9 52 CA 9D B4
 0E DE 3E 48 DC 26 50 65 CC A5 7F 99 BE B8 69 B9
 C7 C1 5A 67 40 72 50 02 C4 1D 8E A7 19 C4 B1 64
 6D 95 4B B8 E0 58 5D DC CA DD 59 F3 9E 90 27 06
 B1 8B FB 1B 37 EC 75 E4 57 8E DD E9 11 32 20 D2
 D8 54 41 95 B1 F8 DE F4 5E D2 48 E7 DB 1D 03 F4
 4F 7E 99 87 7E 65 9B 55 EE DC 4B BC 26 4A 44 C3
 F7 DD 9D 4E C4 DE E0 7A 19 88 1B 8D 6E 61 3C 44
 A1 1C 4A CA 2D 9A D5 A7 7F 2F D1 12 FF 38 DF 0A
 74 DE C8 7D F6 D2 EE 78 BC 42 10 5A F2 98 F7 D2
 FD BE EF D4 77 A8 88 FA 91 12 E0 1F 1F 6B 11 2A
 B6 CD 87 06 F9 73 3B BB 5C AF DE 5D 83 19 77 6A
 4F 2D 28 D2 31 C2 87 10 E3 ED 4E 03 CD DE B5 4E
 E2 0D 2C 10 6E 03 8A C8 16 6B 40 93 AB ED 4E FE
 45 0D 90 E5 64 BD 35 32 F8 C9 86 89 6C E1 11 0A
 92 A9 C1 CF 30 D7 1A D9 9F E8 E3 A1 3A A2 18 69
 66 69 FF E7 5C ED 6F 69 77 28 BB 59 85 26 54 8A
 EF 40 3C E4 DC 2A 04 E3 52 13 5B 69 FB 8F 3B 94
 E8 88 68 1B D2 FC AA 4A 01 32 1B 5E 93 33 3E C2
 05 49 2E F2 23 9F 3D 38 86 9F 0B 7F 6E 25 A5 EF
 69 9A C5 68 00 51 95 EA D2 06 7D E5 07 0D BF C8
 E0 56 45 75 98 EA 4F 82 BC A5 67 2C 31 67 35 EB
 34 D6 20 15 10 AD 74 7C 09 61 87 5F FD 4F 5B 53
 5B 3D 2E 92 98 2C 73 B4 B1 EF 39 94 16 A9 E8 A4
 EB 52 01 B9 27 CA DB CE CD 64 B0 E5 BD D6 3A 3A
 44 34 8B 4D 28 7C CE 07 69 64 BA B9 FA F9 7B E5
 70 1B CA D1 AA CF F6 15 2B 14 02 D7 CA 18 1A 67
 4E 59 6E 18 24 0D 2C B9 B3 F9 A4 FD 59 6E 2A 07
 E1 CE B4 53 87 E3 C6 CB 53 6F 06 C8 D8 40 FE 06
 C3 F4 A7 D2 3B 98 CB B7 16 6A CB 48 2A 68 A9 AA
 50 99 D6 B6 A8 FA C7 78 E0 81 95 A8 84 4C 33 B5
 BB CA D8 E7 FF DF 90 50 A6 9B E9 20 D8 F8 2B 6C
 65 9E 17 85 5A 27 A4 CF 21 DD 32 47 FE F6 0E 33
 B3 47 C5 2D 00 51 80 42 FB 30 67 EE 95 96 3A BB
 26 D8 6E 1F 51 3B 84 B5 D0 38 06 49 98 6E 29 21
 7C 1C 1C 48 EF A4 D8 B6 FB F7 3E 6B 7F E0 E1 6B
 18 9B E7 E1 5B BE 7A 32 98 F1 7B 97 68 95 6E 26
 1A FA DA 55 18 F6 5D 91 E0 03 4D 50 36 AE 86 CF
 43 31 64 B6 C3 0D F1 C5 E5 EE 2A C3 E2 16 94 24
 27 4D B0 D5 24 C1 79 C4 54 1F A8 47 10 52 28 11
 FB 4C 81 E4 3F B7 0B 95 08 69 BB EF 64 E6 A3 E4
 39 E8 16 16 34 B0 EE 4B 99 EA 81 7B C5 BC 7A A4
 F8 18 AA AD BE FF 3E 07 D7 07 2A 60 3C D3 4E 9A
 2D 96 7A C9 C3 C7 EB A0 77 1A E8 FF D7 8B FF 28
 27 A1 A5 74 1C 1F C1 5B 3A CC 4A 78 6F A6 09 1A
 BC EB 0E 9C 17 79 83 5D 0C FF 37 CD 5B 8B 20 50
 1F F6 55 DF 83 B0 9F 2B 43 9D 22 DC 61 67 C1 5F
 70 10 51 B6 22 13 C3 A1 28 A5 B2 3A E5 26 5F 89
 24 BA 22 5B F2 BB C1 15 98 0F 13 2D EA 92 89 5B
 13 B1 47 76 3C 4E C3 03 30 51 56 CE 8C C3 CF 27
 D4 DB BB 21 73 7D F3 D4 C4 17 9D C3 5E 43 F7 7C
 82 7E 5B F1 1A 19 24 32 88 A2 8F 88 B5 8F DF A2
 16 B8 E5 47 0C 4F 23 9F E0 2B 22 7C DA AA 43 F9
 09 FD 78 2E 3D 86 99 FC D6 26 7E 32 19 25 A5 9D
 0F DD 5A C7 87 82 71 DE C5 27 A9 4D 42 20 A2 A8
 A5 12 56 A2 CE CC 98 C1 1D 64 0D F9 26 73 8B 4B
 A9 E1 75 FF 82 17 9F A1 4E 9C AB 46 40 AE 0D C4
 92 51 CD 05 CE 61 CB C2 90 13 8F 83 3A D3 30 72
 28 8E 10 60 AE 0D D4 DC AD 96 7F AB 2E DC 69 65
 A6 FE A8 96 C4 97 16 73 BB 34 D9 8D 75 CB 76 00
 AB 47 1A B4 6E 5C 14 41 1C 47 05 01 A7 CD AD 0D
 B5 99 53 55 15 D3 BD 64 C8 28 E9 7D 1A 56 EA 5D
 71 45 77 1A DB 8F 79 4B 53 97 A8 46 50 B2 62 AC
 F1 7C 2A 28 35 18 14 7E 47 69 02 45 49 B5 73 F4
 B2 13 0C 26 E4 00 E7 71 FE 71 48 DD BF B6 E3 72
 01 B3 74 21 55 74 C1 E0 CD A9 5A CA 3A FE DE 20
 5B 4E A9 6E 05 3E 76 A7 1C C0 56 DD EA D7 1B 1C
 24 F3 7F 91 3E E3 63 FC 14 4D 8D DD DB 82 4D 61
 62 04 62 FE FB 21 8D 37 FB 9B 47 E9 26 11 FD D7
 78 5A F9 D2 82 4B 53 99 E0 58 28 30 38 A7 63 18
 06 B7 A4 22 E5 6D A2 6A 38 E8 EC 1F 34 4C E6 68
 06 D2 84 1B FD CC 8A 5E BB 53 74 43 8F 30 D9 31
 0B 19 A7 5F AC 39 F8 8B C4 48 E8 09 12 4A EE 69
 FB C8 68 D9 A0 BF A6 52 9B 0B 80 E7 36 9C 40 7B
 47 21 DC 72 85 7A C6 F3 BE EC E7 76 DD 22 C3 F7
 20 D5 94 E8 02 DE 0B 8F A6 6C DF B5 C8 A1 D0 08
 E8 FE FF FF FD 8F 60 1B 23 21 B1 E0 74 7B 89 DD
 46 2D E6 3E 6E 10 2A 35 12 B5 95 11 9B 36 75 1A
 4E 32 F1 21 09 3A 70 4F 1A 11 0F F2 0A 5E C3 0E
 0E B8 DC 3E 8B 17 9B A5 4F 29 DC 4F AB E7 4B BA
 17 B4 1F 91 2E 43 41 0F 69 A9 0E 8A A6 05 5A 36
 29 C2 AB 73 A1 34 6A 23 E8 0E 53 29 22 E3 11 48
 DE B5 4A B4 C5 69 A2 3A 4B 15 EE 47 5E A8 B3 B9
 14 9D 57 8C B9 0B C8 65 17 32 36 5B 84 FF D9 69
 46 3A E2 86 B9 25 85 C7 B2 EB 2F 20 78 F0 B3 06
 21 2D 53 17 99 88 20 40 24 B7 07 A8 48 13 CC 06
 F0 56 C9 D9 D1 8A 84 AA CA C4 68 5F 4D 6D 29 EE
 C0 51 66 BA 03 B4 C3 2D E2 9C 8A 33 EB 56 72 43
 76 92 80 2D A4 E2 6F 31 17 E2 3E 9C E6 38 AD 68
 6C 9F 6F 9D E9 BB D7 71 40 6A FB 27 D4 CE 25 9E
 38 F5 28 5A AB 0C 81 45 CB 72 AA 8D 1F 43 45 96
 0F 17 E9 F5 61 5B A1 8F 11 30 08 24 6D 44 D8 9F
 82 E8 C1 62 DC B5 E1 72 36 B2 B1 1D 6C D9 64 C0
 DD B2 13 47 C6 7B 55 34 5D 23 10 5A F3 74 CE 5C
 C2 AD AC 3B EF B6 0D 66 41 4A B6 1F 7E CD FD E8
 77 8A 57 7D 45 94 FF E0 29 95 DB BC 42 D7 FF 38
 DA 37 1C 8A 5E B3 00 37 B0 49 98 18 54 1B 82 36
 9B B3 1B C7 9E 70 3A F0 FA 40 A2 15 5C C7 39 93
 DC 74 FB 54 F3 A3 E2 3E 8D 36 39 91 6E 4D 8B CE
 E8 A5 8A 34 9C 0C BD EE AD 0D 0D CA 8E D2 46 C8
 E4 16 25 5C D7 F7 48 B9 78 12 1B 5D 7F 60 15 30
 1A 5F 33 FB 5C A6 53 B6 F2 4E FD 23 F6 E1 9A 03
 40 22 D6 47 94 BE DA E7 F4 F7 80 D8 39 EC 12 A7
 51 72 96 20 EB 77 32 ED D8 26 32 C8 F3 30 5B 74
 D0 B9 A7 D1 0A FD 56 DC 43 16 22 58 F0 FB B5 0F
 21 43 48 31 04 90 D7 66 35 D8 27 E5 04 E2 6D 67
 EB 2F 60 47 C8 76 12 A0 25 E8 42 67 8C C5 E6 7B
 2E E2 6E 9B 50 C0 74 DF 7F 40 8C 68 80 BC 1E F4
 8B 91 A7 0E B3 7D 72 C2 60 0D 3B 18 9F 85 06 FD
 44 40 98 9F 5D 07 20 97 69 52 7B 1C 9A 3E 1C 57
 CF 77 9C F5 BD 9B 3D CC DB B8 8A 7D BD 98 E7 4C
 D3 58 5A F3 EC 24 9D E9 94 D8 3C 8E 0D AE 2F B5
 2A 7F 45 14 B9 34 4F 78 E2 D5 11 75 4F E0 C0 D9
 CF 68 45 50 81 DD 18 18 51 58 5B D0 4A 3D A3 BB
 4F 1F 22 40 05 5D 67 ED B8 36 EC 22 8B 10 1A 84
 40 B6 94 C7 19 44 38 77 28 A0 F2 1A 68 6B 91 CB
 0A D9 CB 19 CE F2 D6 E9 B8 4A 79 26 7B 32 FC C6
 77 86 E7 81 71 C0 53 37 B5 8B B0 32 C8 C1 8C 1D
 7A 46 1E 3D F4 B1 06 03 D4 5A 9B C3 FE 0C BB FC
 01 3B E1 D8 E1 AB 1B 4A A0 7A 6C E3 36 FA 83 D3
 AD 88 82 4C B8 33 87 EA E5 65 B6 A0 4A 5A 32 63
 C2 D7 8C 13 86 99 2D 12 DE ED 4D 2D 14 F1 BC EF
 1C 46 F0 2B DC 0E 57 0A AF 1B F6 50 20 C3 6C CB
 DE CA 01 B3 83 63 35 B2 B9 CC A9 37 91 06 68 85
 BF 12 4D F9 A9 26 8F F3 08 D8 17 F9 10 CC 49 0C
 8D 83 7B A1 2A A0 CD 11 99 E3 5B FD EA 7E D5 D2
 CC A8 FC 15 A7 EB 35 CF 61 8C EF 1C BF 7F F6 39
 41 80 52 A5 02 C2 94 13 A9 7B A4 12 DE 6C 0A B4
 49 D0 DC D2 C0 09 D0 0F 11 A7 F7 50 7F 2B 13 54
 4E D5 F4 AF F0 E8 51 A7 0E 70 0A A1 5E 2E 0B AD
 66 50 F8 72 54 11 C0 D9 2F C0 6B CA 77 52 31 14
 FF D2 78 C2 0A 02 7C 5E 35 42 54 C3 7F 75 B4 46
 63 EE AF 21 A7 2E EF F0 C4 3D 9E 2B C7 4C 4D 72
 EF D8 46 F7 16 C0 8B 00 12 64 58 40 C2 C8 DB 45
 EF 9A E2 66 AC 66 A6 07 D1 02 90 E0 1B 8B 61 92
 12 81 28 55 ED A6 44 C2 C6 F4 C9 0B 62 D4 7B 5D
 BE BF 35 30 04 EB 4E 0A EA 72 F9 03 9F 17 68 1C
 CB 44 B4 0B 6A 32 23 A0 DE 81 B2 E6 03 0C 6B F0
 FF A2 1B 4E 09 C9 11 AE 85 42 3A 37 7D 58 CF 39
 1E 67 1F 39 77 A9 24 9C 37 5F F4 DE BC 84 ED 31
 68 77 D8 DF 9E F8 FF E0 3C FB 94 D8 90 46 45 DF
 73 0D D4 2B 33 DC E7 37 F1 D6 9A CA 37 94 79 7A
 9D 91 DC 3F 50 3D 1F 44 9A 89 43 EC E7 61 95 1F
 E5 96 7B 8B BC F9 59 9B C8 27 2E CB E9 D0 06 10
 A8 DC A6 A9 1C 1D 8C 71 B1 8A 3D E1 B2 22 F8 EE
 9C 9B 58 B1 A2 5C 39 A6 D3 A3 0F BA 5A 66 AD AF
 85 B9 AC F2 8E 54 3F 24 67 60 C0 C3 6E F4 81 DE
 B1 19 F7 30 79 C7 14 E7 01 8A AC 49 83 F3 1B 3D
 83 99 FD 8B 92 A7 E7 0F F1 0C FE D8 E3 D4 FE 5B
 A9 66 29 A6 C7 3F AF B3 68 25 4F 97 B0 3B 02 E5
 DD 50 B2 3B BA E5 19 65 7B B9 3E 7E 8E 37 C4 AF
 38 4C BD 3B E0 4E AA 0E 07 AA 08 4E A9 98 A6 5A
 EB 1E F5 1A F0 E8 6B 2C 64 AF 2E F2 58 71 4C 65
 80 25 33 63 9F 82 EF A5 C2 B8 73 70 A4 DA 5A F3
 5B 2C 0C 4C 52 D1 C7 D3 FA E4 3D C7 7B 4A E8 79
 D9 7B E0 E9 0F 2F BA D5 E4 2B 42 CD B6 2B 4D C6
 6D 72 E1 63 FB 04 DC B3 68 5F B4 0F 9F 83 85 8E
 7B BE F9 D0 9C A5 15 04 7C 4D 80 38 34 66 28 E7
 C5 BD 67 85 46 DF EB B4 C3 4E 50 E7 21 4C 13 DA
 34 BD CF C2 23 CC 7D 04 64 53 CE 0C FF 19 8D 72
 17 6E B5 E3 EB 3B 6C 88 6A AD C2 A9 19 C7 D9 2D
 D2 53 97 C8 0D AE 7F 21 BB 8E 4B B1 49 07 0E DE
 19 1F D2 42 81 26 FE C8 29 A9 F5 43 89 D6 50 B2
 3B 3C 14 4D 4B 59 60 F6 21 82 5F 48 11 BB DB 3C
 0E 1A CC 40 BF 78 44 C6 B8 B2 47 2C 77 74 10 9E
 CC 6C C2 F4 A4 EA 73 33 DE F1 51 95 87 C2 0D B6
 90 30 F4 3B 0F 41 45 41 86 5E 23 A3 52 8B BA E0
 92 A9 70 50 F9 E1 00 CF 10 24 5A E7 6A DC 77 0A
 FA 38 DA CE D1 04 26 AD DB 79 E8 FB 0F 09 89 C4
 9F 8B 8F 3C 98 FB 6B D2 46 D6 1E 99 6E AB 59 E6
 15 6D 36 3F 6F 7D 06 AA 81 26 0A CA F5 2C 1F AE
 16 BA 50 BD 91 0E B1 96 46 C9 A7 4E 0B 6E 0B B8
 7F 87 4B 07 CC 1B 3A FF 36 89 FD 8F 63 A8 E2 ED
 87 F0 38 F4 EC F0 CD 22 5E 3A 29 2A 48 A7 21 07
 1B BA 74 9E 20 B9 F3 50 B1 AE E9 A1 21 32 7E 43
 2D A2 27 C6 0C 78 7F 04 CE B5 AF 38 DF 8E 50 F3
 3A C4 6C 68 F7 86 E7 18 73 1D 5B DA 1A C6 C8 92
 9F 36 2A D8 D6 78 26 1C DE C1 EF 6C C8 4F 0D D4
 83 79 6C A3 90 3C 7D 58 F7 E6 8A AE BE BB 6C 12
 A8 EE 88 B3 44 92 F6 D6 EB B4 C7 46 CC 74 FD 65
 34 3C 4A C1 5E 58 07 59 E9 C1 3A 22 B5 A6 7A 44
 0D BF 9B F0 7B 8D 89 D4 22 6B 9D 6D 10 C4 0B 23
 24 21 59 E1 5E 4F 43 5A F3 BA 7C F4 4A A2 AB 21
 0E 56 88 1D 5F 14 14 13 01 A4 88 0D 6C 20 9D 25
 43 70 EA 0F BA 94 94 BF 59 F2 43 A4 50 F3 A2 D0
 D5 74 FA F6 EC 87 26 C7 60 2A FF A2 F9 C9 AE 1A
 BE 17 D8 22 F8 F1 6B F8 A6 13 EA CA 7E EB 0C 6F
 65 F8 89 D7 10 02 0A 2E A7 B6 5F 50 37 CD FB 65
 0F 6D 6F 75 B7 08 9A 44 E1 57 FD 35 B6 B5 4F D4
 F7 CA 9C DB 45 6C 45 B7 92 82 C7 26 60 13 89 29
 C5 96 90 BF 15 8F D6 E3 3B 18 A2 22 78 EF 92 40
 C2 E6 7D D7 8D 2C C8 52 10 56 28 F4 77 48 C2 79
 58 45 99 BC 25 9D CF 99 B3 C2 06 01 F6 8B 2B 1F
 09 8F 30 94 0C 22 E2 7E F9 95 18 05 2F 33 E3 36
 2A 6E AA C8 06 F8 6A F6 9A 61 A3 66 57 FF F1 26
 45 48 94 2F AF 4F C1 28 31 54 13 B9 C3 88 88 17
 71 FD E3 78 88 A8 7A ED B4 74 9C 4C C6 B6 97 7F
 A2 4B 95 10 10 5E FD 0B BE 1C 54 C9 E2 9E F6 72
 C7 30 7E 12 86 39 21 AC 21 C4 86 CE F9 CD 44 6E
 EC EC FF C4 37 FA 99 18 EF 90 8A 7B B4 10 1E 91
 D5 73 34 5F 98 99 7A 2C 27 03 D7 EB 9E 68 0B D7
 42 70 ED E1 4A D1 B1 F1 F3 B4 B1 CA 30 6B CF 2E
 56 B3 AA 98 2D 86 37 D5 DB 2F 47 4F 72 A5 93 DF
 B1 2D 89 11 7D 87 40 C9 50 77 A4 0C D0 E6 88 94
 8E 0F 30 F7 EA 00 56 1F 29 67 54 71 38 9F 73 B7
 0E 60 1D 83 2C 82 5E 50 83 28 43 7E D7 ED 70 14
 40 F8 76 51 47 BE 10 68 68 BF D7 59 CA A0 8E 38
 7D 17 7C BC F2 1F B9 AA 6B 47 95 CA 6B DD 99 D1
 D5 42 29 91 BA 7C F7 36 76 B4 A6 4F 5C 57 25 31
 99 A3 5E 72 99 F0 97 5A A6 3D 78 BD AD C1 C8 5D
 DB A1 3C B4 BA 24 F0 04 2D 73 3C 4A 5E B2 A9 1C
 C4 3A B9 3C 4A ED 07 2B 21 98 E2 EE 00 6F 09 7C
 5F 38 01 F8 C5 A4 8B 7F 5D 99 8A 2D 91 0F 7C 41
 4B E0 4B D5 08 62 58 D1 B5 81 B3 89 F4 97 DB 9F
 44 3D D6 1C 4A 52 18 4C BA 22 03 43 F0 A7 E6 CC
 D2 AA 00 E6 8A D5 9C 45 4F 88 73 01 37 15 81 97
 10 86 F0 95 85 B2 5D CB DE 1F 23 72 66 07 25 01
 FD 33 09 4A 8B 78 FB 0E 5F 67 A7 1C 77 A6 E6 07
 63 F3 85 94 65 B9 CE 4B C7 E8 A3 63 0C BC 30 B3
 57 07 BB 06 B7 17 00 0A 72 95 02 08 9A 50 01 60
 91 50 1D 97 C2 38 82 E1 C7 1D 10 55 0F 5F A8 75
 6D 14 DD E4 E4 DD 68 3B 9B 00 9D 0B BA 55 25 57
 3E 7F 4E E8 E7 A4 C2 BB ED A4 22 47 04 0F DC 35
 CD 73 5D 2A 5B 62 8A 73 F8 0E E9 ED 55 98 0C 1F
 FD C6 55 7E 6A 33 98 99 B9 08 2B D6 24 08 92 79
 5B 51 8A 1E 72 19 C6 9B EC 50 28 91 A2 54 D8 A7
 05 76 2D E2 C2 60 1E BC 3B 07 B4 24 F8 D9 BC BB
 7E 5D CF 25 CA 56 87 FB 5E EA 1F 9D 6F B2 BC 8C
 23 6B 31 8C 1C BA FB B2 0B F5 EA 89 24 04 98 49
 D6 25 E4 E2 AA 48 DF E4 36 83 A5 22 54 ED 26 C3
 BD E7 85 0A 62 2A A6 39 91 53 C6 11 EA 54 80 B6
 5F 49 54 5C F5 1A 5E 8A A3 A4 B9 18 B0 52 65 FB
 E2 25 B1 D5 FD B7 D9 62 EC BF 60 57 C9 17 6B 90
 5A 05 8A 48 AB 7D B8 52 F2 65 58 AD CA 92 11 05
 E8 7D 75 C8 11 A9 95 07 AB 03 88 16 A9 7F 31 24
 0A E2 A0 86 89 30 72 C1 91 28 68 F3 27 2C 3F 6C
 78 9A 22 9A 84 33 A3 72 C3 7F 9A 3B 72 09 7B A4
 8A FD 1B 5F 7E E8 EB 98 29 6B 8E 2C DC 20 EF 78
 98 E6 97 65 27 67 1D BD 15 18 83 01 3E 08 3D 0E
 32 BC 44 42 45 6A 09 AF 85 E5 E3 B2 80 78 F0 BC
 AA D5 93 3B 4C B4 BE 50 CA 66 F5 CA B5 60 D6 09
 F7 0B C4 E7 C4 16 3B 87 93 2D 27 19 AE 49 B2 2E
 92 CE 02 C0 65 F4 DF DE 3E 38 47 8B 1D 91 1E C5
 5D 6A ED 18 31 8A F9 A4 60 D0 E9 34 E2 76 CD AC
 0A FF 9F B2 4F C1 68 20 44 93 7B 78 8E A5 77 2A
 9A 51 2D 82 E9 65 68 0A 7A E9 77 91 31 CA 5D A7
 DD C0 A7 31 20 7F 81 85 FA 0D 9B 0F 18 45 25 B9
 7C 53 2C 37 60 6E 50 39 63 90 15 80 E9 B2 0E 8D
 10 AB 93 DA 66 BD 53 B6 4B 40 40 22 68 E3 E9 36
 18 F1 45 04 41 44 3E ED 05 9A 75 EB 1E 0C 5C 53
 8C DA CE 7A 40 28 6F 98 5B 8D 9B D3 9B CD B7 0E
 94 A4 C1 E6 C1 9F 7F BD 15 FB 9D 58 00 67 A8 9B
 2A 77 92 A3 EC 88 71 5A 8F DD C9 0F 9B 0B 8C 2C
 8B 17 22 A4 1C C0 13 EE EE 91 11 A5 8E 83 86 8B
 9E AA 40 20 DE DF BD A3 43 41 75 A2 C6 96 9D 83
 6C 23 4D 46 7A 21 EE 46 64 3B 3D A9 AC B9 2A D3
 81 97 AD EA A2 F5 79 DB 60 20 C0 41 8D 4D 10 75
 89 4D 1A B1 0A 49 BB 1A 8E 1D 0A 31 7F 07 E1 18
 F0 63 C7 F4 E3 40 12 6E 09 E6 E4 19 67 57 3A 14
 0B 82 FB 84 CC D1 A7 DE 55 87 9E 1E BA 04 86 E6
 1C 39 7F F9 64 74 84 FF 94 E9 E9 60 8C 49 84 AA
 8C FA 97 C2 59 5A D3 8F F4 3D 95 F3 54 1A 6F 33
 94 17 4E 5A F4 B2 D9 BB A4 6B 54 5E FB 28 CC 19
 D0 65 BA 63 9A AE 32 53 4A E1 E7 03 4A 55 18 D0
 1D 77 25 21 2C 64 B7 CE F2 C9 A3 0C D0 4D 6E 8C
 47 44 66 F6 6A E3 4D 2E 17 3A 52 8F 79 73 E9 AF
 1E F7 7A BC C0 37 A4 98 A2 5C 18 25 AB 8F FA 27
 EC 51 33 1C F1 D2 43 59 DD 87 90 C7 72 9D 00 5C
 76 6D 21 E3 41 1D B2 15 E7 ED 07 58 D1 66 06 54
 13 12 A3 4C 4A F1 B5 57 1C 12 1A 94 99 B5 94 F2
 6C E3 C7 13 99 87 B5 E8 B3 82 9C 14 64 E1 CB 8A
 FE 53 8F 1B 45 9D 65 2A 2A 00 ED C1 9F FE 7E 65
 6C 11 71 12 A7 4C DD 79 19 76 0F 07 7F EE B7 42
 81 62 0F 23 80 C3 F2 A7 9A 44 38 F8 21 BC F0 2B
 59 A5 14 CF EB 82 D0 86 C5 DE C9 D5 52 EF E4 E7
 07 89 00 34 6A 91 B4 30 80 4D 81 24 7D 06 CB 00
 22 1C 30 13 F7 DF 30 8E 21 65 25 6E 95 6B A3 BF
 CB E3 38 03 31 90 AC D2 6F F0 9B 77 FB 61 30 22
 55 5B 3A C1 44 E8 4B B5 B5 1D A1 F5 3D 31 FD 3A
 1A 68 B6 98 91 40 4E C1 EF 27 BA 36 04 75 D6 EC
 35 C2 32 03 D3 2D 3D E7 E2 B2 D2 A9 7A 6D 1B 08
 6C 91 75 7A F0 69 4C 26 9A 86 AC 64 9A B0 D1 36
 16 E4 FE 5D 8E 79 69 30 5C 9D D0 02 FD B6 B5 37
 40 C8 D2 59 14 1F CD 8F 51 66 8F 58 C0 7D E8 33
 B6 AF 13 C1 BB 1A 1B 4F 28 9F 7C BD B6 F1 99 93
 7F 88 4E D3 9B 0E E2 60 76 76 15 10 F7 3D 11 D0
 78 A3 7A 76 6F FA 06 2D E8 BE 40 E1 E5 A9 3D 6F
 7B 1A B0 E5 F1 90 F5 51 C3 92 5C 15 4C D3 16 38
 E2 F1 28 CE 58 01 84 87 9C 88 C3 0A 8D 0F F8 9A
 D3 C3 D5 F7 48 4E 8F CC A2 90 B3 B0 3E AD 36 DD
 64 3C 27 75 DB F5 CD 1B 5D 4B FE A5 5A EA 26 92
 2B DE 2E C7 B1 EC 1C 94 01 42 42 39 1E E4 E0 4C
 5F FC C8 71 FE 18 C5 05 5D A9 D2 2E A1 C1 08 34
 7B D3 78 22 A1 28 99 EA FC C4 57 CC 10 35 87 09
 C6 A8 F5 58 9C E1 D8 3D 9F BB B6 8D 5E BD 01 A1
 7C 56 2A 26 FB 0F 43 6E C8 F2 FC 31 15 DF 87 8C
 CF 8C 30 92 90 3E 14 91 ED 46 23 CB B3 E2 05 2B
 3C 84 26 EE 4A E7 AE 53 05 41 C7 15 B3 0E 0A D2
 1D A7 2C 73 22 06 C2 6F FB CF A4 EA AA 8E 51 D6
 DE 53 14 13 D8 FF E0 C4 F0 E0 93 96 D0 8C E6 00
 81 0F E1 76 D1 2A BF 0E 01 81 FA 2F 92 94 B0 07
 4B 8A 1D A3 7A 86 B9 7E 55 44 86 0F 3A 5E CC EF
 D7 48 5F 20 3D DB 0A 90 FF F9 B5 FE E8 C3 F8 34
 47 32 4C CA 84 33 BC E1 EC 0F 9D 9B 3E F7 62 14
 C6 B5 93 EB 20 B3 CD 99 EA 05 1D DB 69 3B 32 D9
 20 CB 1C 56 2E CD A6 7A 76 ED B4 0D AB 92 30 07
 38 EE 92 E4 69 89 02 A2 36 19 CA 9B CC 11 D2 BF
 F9 EC A7 7B D9 AF D7 69 C5 7F FE 98 95 16 75 93
 71 38 85 4A F8 D0 31 59 5A 75 DC 55 E6 DB 8D D0
 EA A7 F9 2B 2D 52 FA 1B AE 82 DC 16 84 9C 84 0E
 E5 D5 D7 95 44 F4 54 9D 15 75 6A 54 BA C7 15 00
 D1 64 C0 8B 1E 76 03 04 F8 51 77 1B 65 88 2D 30
 3F 4D 54 67 18 82 55 FB 2D B7 3C F7 F6 0F C4 4F
 7A 6E 73 BE 08 33 61 8C 9D 3D 0A DE 9D F1 84 64
 E8 B2 79 AB 27 EF 72 92 F7 23 40 FA 9B E6 ED 94
 C6 3B 5C 0D 3B 2D FB B3 3C E6 E8 99 FF 57 95 11
 64 47 E8 7F 6B EA 72 46 A1 9A 1B 7D CD FB 17 F8
 37 01 6B 73 F7 FA A0 91 BB A0 D3 97 51 DD 6B AA
 09 74 8C 6A 93 57 41 A8 13 0B 9B C3 5C 53 EA 04
 FB D3 36 5F 66 BF A7 E7 11 D5 FC 5F 66 27 04 1E
 41 40 4D D0 2C 2A 47 83 CF C2 D9 17 B1 6D 8C F2
 AD 26 68 66 1D 78 1D 0E D7 4D 16 83 25 BE 4E F5
 30 95 05 8D 05 CA F4 D7 D1 F0 A1 B7 2A 3D 48 65
 3C C3 FD AC 79 8E E2 6E 29 04 9E 48 E3 E3 40 67
 32 84 0A 58 F5 10 9F 15 2F CC 7A 84 03 A4 31 8A
 43 22 75 50 66 A2 D6 7B BF 29 27 13 E0 BA 17 C6
 27 2B 4F 6D 06 B8 5A 09 49 F2 CC BC 5E A9 E9 B9
 B6 27 F6 26 38 F2 76 F7 C7 8F F4 7D A1 A8 27 FA
 61 AF 06 C4 2B 3B 1B 20 06 BF 59 D4 F4 0D 66 A6
 DB F2 8B 23 B0 2F A3 4F 89 EC 16 CE C7 E0 1A 88
 1E 5C B9 41 7B 57 8A 86 30 4A 25 53 A3 96 00 D3
 B3 35 46 FA 30 5B 23 68 14 1D 16 40 1F 47 50 9C
 50 14 9E 3E 50 3C 55 1B 3A C9 B1 EC CC 2A 59 00
 CB 45 E0 CF D4 77 BC AE CC C2 3A F1 11 24 88 17
 15 A0 6D 68 C6 20 B8 79 8F 5A ED A4 E8 62 C7 99
 C3 A1 00 E8 EE 3C D9 9A 16 2F 62 30 87 BC 29 78
 F8 9E 72 C9 71 32 B0 35 F3 C7 1B 80 BC 1D 3D 88
 DE B8 5D 7A 88 29 07 EA 66 D2 B5 C1 A9 B9 42 42
 5C 9A 1B 45 D3 4A 3D 95 BE F0 90 39 8A 47 E4 F5
 47 3E 51 58 61 AA 62 6E 8C DA 35 FD 09 19 5B 09
 88 93 12 CD 86 B4 16 FA B1 A9 BD A3 05 D1 AC 46
 21 C6 E4 98 77 14 3A DF 3C 5E 6F 36 79 ED 3C 13
 BA 7D 38 CB E0 8C A0 E6 59 C3 45 F1 15 9F 8E B0
 51 12 8E F2 1F 3B 21 C4 FE 9E C2 2A 4A ED 9F 23
 CF 50 6D 37 B4 F5 09 CC 2B 04 4A E4 01 BB B3 26
 94 CD F8 DA EB 7D 1C C6 C6 AC BE CD 49 0B F7 BB
 BA DB 7A 3F 41 2E 1A 10 C5 E1 47 72 2C 51 F4 5F
 73 8C 7E 0A D6 49 F0 45 7A 92 77 96 FC 5A C0 3D
 21 3F 6D 66 BE FC EC 6B 69 97 88 33 8B 42 87 8A
 A0 34 21 1D 09 FC 24 8F 76 26 F4 3E F1 A9 AD D6
 2C E3 29 C0 F5 B7 84 91 4C 47 40 2A F8 86 55 02
 0D BC 97 89 4F 7F 8F AC 13 04 F1 0C 41 C9 DF AB
 35 A5 00 E7 08 89 30 46 88 5D 76 20 7E B6 76 98
 7E E4 54 0E 21 A5 D7 3A 98 10 03 A6 D1 33 EA 4D
 2F 88 81 04 2E 99 1F 2D 2D 8F DF 63 1C 8C D1 19
 64 14 5E 7D 6C CD 0E 60 76 58 AC 58 AE 84 78 C6
 FC E9 C9 50 79 F8 4E 8B 6B E7 46 EB CB 95 BA 25
 CE E9 EF 97 B2 78 59 71 A0 75 82 59 1E 3D FD C1
 8C 1E A0 51 76 A3 B4 C0 7A D2 66 59 CB EE B4 86
 4B 7A B6 E9 B7 F8 1C 22 12 41 DA CB EC E6 4A A0
 A6 6D CD D1 ED D2 27 EE DB B8 FC FE 7F DE 59 62
 83 B4 9F C0 76 F5 53 A8 7E 01 66 28 56 7A EF 31
 39 95 FC 9A 1B 25 FE 6D 8B A8 93 A6 DA C4 EE 86
 42 12 86 5D CC 34 B7 D1 C8 95 59 F4 34 6D 40 B9
 FD C8 23 0F 63 4B F7 A8 C7 80 8B A3 5D 88 62 90
 C3 A6 27 33 F7 4E D4 AC 4D 5B 05 D0 FA 05 54 58
 AA 9B FF A5 94 CC CA 19 9B D6 4B A2 81 4C 76 05
 3C 98 54 57 2D 24 FF 7C 06 A3 C7 E0 AA 75 F8 5D
 46 99 77 4A 55 4D C1 1B 4B 8F CD 40 55 09 62 BA
 B4 8E B7 CE 98 BA 4C 6B B6 1C DC A4 32 BC EB 07
 74 50 05 E6 7A A6 CC 5E 80 FE CF 97 FB 4B EE CB
 33 73 0F 8B 1D 6A 30 84 AE 52 04 A9 B9 54 4C BF
 54 1E B3 AB C1 00 49 8A A3 4D BC 99 E9 5C 33 9A
 DD 3B EB 86 40 C9 EB 26 5C E5 E5 28 ED 3B 1B 61
 FD 1B 2D 40 2E 94 A9 3B C6 F1 14 6C D4 EC FF E1
 91 CB 8A 05 A4 45 33 58 B4 8E 9F D6 47 C5 5A 09
 59 10 E9 44 8F 2B 70 DC B1 FD 5E 08 F9 EE 52 2E
 40 CB B9 AC C4 D7 8B 7F 18 85 4E 95 7B 73 72 05
 8D 5A 51 B5 C1 CA 78 9A 3B 96 12 AE 86 49 6D 24
 DF C4 B1 61 FF 81 14 A7 13 91 E8 50 61 0A 48 2A
 E2 5D 77 FA 82 61 7D F4 DC 75 CF 5A 8D 27 D2 76
 C5 00 F4 02 66 2A 27 C3 35 FD 95 72 17 BB 9C 89
 DC 10 C7 4D 82 46 53 E7 68 05 86 16 58 01 82 3E
 05 79 B2 0A A3 62 81 A1 A9 E0 05 73 0C 77 7F D2
 82 7C 81 69 D8 B0 AA B5 2D 6F 30 8B 8B 09 45 C4
 8B 53 B8 F5 8C 50 56 B8 DE E0 F6 F4 39 22 D7 E8
 C4 52 0F 9C 01 27 0E 0B 93 2A 9E EC 8F 79 E5 C8
 92 C1 C1 34 29 B6 CC CF 86 3D 4D 4B C2 BC 82 74
 F3 8D 1E 08 8E CE 0B 43 9E C7 23 02 26 91 50 3E
 3A 0B B3 50 2D 58 40 64 AB FC 36 46 58 F2 4E 3D
 29 9B 56 7C A0 27 F8 B4 AA C6 D2 AB 80 80 C7 E9
 D7 73 8D 9D FE 9C A6 DA 86 EA 7F 14 FF 94 DF D8
 42 D6 89 81 CD B1 1D C8 1E 20 26 56 78 6E 1F AE
 50 67 3E 71 B6 11 87 29 78 22 24 1D 33 20 2B 74
 13 3E 16 35 56 E8 B2 11 DD 96 AF 1C B0 21 AD 7F
 CE B7 56 00 57 3F 5F 05 CC 68 EF D4 1B D7 5E 56
 EA 86 49 88 9D 16 DC 03 66 E0 C0 AD 13 B1 C4 F1
 B1 86 E8 E5 2C 89 BB 6F 07 B9 70 9A FA 70 E5 C6
 09 AA FA 45 7D E7 A2 C7 32 30 2F 14 0F F7 09 EA
 0C 65 15 A7 F0 A7 3B E4 D9 C3 B3 72 44 95 70 58
 C4 BF 07 58 D8 13 54 0F 1E 42 41 C6 6A 99 BE 76
 54 7A 28 7D F1 9E A1 03 65 0C FD 7E 56 E3 32 A4
 28 B7 A5 0E B1 93 EB 71 93 F8 C1 C2 0E 51 35 40
 24 93 A8 70 20 6D C0 D4 43 F0 66 5E B1 67 26 60
 61 EA 48 4B 9C B9 68 58 EC 05 75 E0 EC 28 5C EA
 61 72 BB 24 30 4E 05 EC 99 EC 84 11 3C 5A 9A BE
 A2 9F 0B FD 0E AD 0E 7A 13 89 F6 C9 5D 6A DA EB
 98 7E FF B9 66 3F 42 D2 87 84 48 42 40 45 D9 F6
 82 47 8D C4 5C E6 25 CA 58 F8 2C 80 9F 37 40 15
 58 CD 3B 4F 07 46 CA 45 20 BE 64 BC DF 44 63 95
 7A 94 A1 13 E5 80 E7 F2 B0 8E E6 EB D9 72 D7 27
 BC A7 E8 4A FC F2 6D B1 42 C6 38 92 DE 48 A9 BE
 AF A6 52 EA 2E E9 35 D5 7A D9 47 5D 6A 1E 60 AE
 BB C9 4E 5E 62 1D 4D 53 46 6C EA 25 C6 A2 1B 59
 33 91 35 39 E6 00 85 09 C5 CD 0F 74 58 ED E5 C0
 29 D6 D3 9D F4 F7 7C 91 A3 8E 5B 2C 1A 76 C7 E0
 D8 33 1B B7 30 58 4D 1F 6B 5B B3 C3 57 09 B8 5A
 A4 AB 23 C8 F6 15 BE 98 B7 3A B9 BA 9E 6C 77 94
 0C E0 A2 9C B6 B3 96 72 17 9D 8D 35 BE F6 B8 BC
 37 88 FE 08 DB 0D A3 4F C4 FE C0 91 B8 52 7C BF
 B5 A6 E1 7E 2D 54 2A 44 EC 3E 7E 64 AA 18 2D BF
 B7 FC DE C1 B2 76 28 6A 44 FC 7C BE 2E 6C D9 97
 F0 5C 12 C8 04 6A 4D 55 AB 8F E1 20 72 31 C7 43
 D7 9D F9 8A A1 D2 90 90 E7 DA 03 38 40 C6 D4 4B
 88 D5 D8 22 63 F5 2F EC 6A 19 02 DB 17 34 27 89
 7A A4 B9 A8 23 D7 8F 2E 9E 83 BE 40 35 54 E0 7B
 76 DD 8E 2C 84 57 1D 5C FC 39 AD D0 3E F1 44 91
 05 27 73 C0 50 D9 D7 1C 36 32 1B AD 72 07 72 09
 BA FC 6E 56 A8 D8 13 65 AC 9E FF 92 24 E1 F8 32
 8C A6 4F 73 01 B6 5D DD BA 41 EB BD FE ED 78 2B
 3C 97 59 AB 32 D6 46 D7 3B A8 5A 52 1A 27 61 4D
 04 2C 9F 33 FC DE 0B EA 36 C6 9A 01 DD 56 4C 92
 AA 6F 25 77 B8 39 C1 B4 8A 0B 8B 4D 96 19 F9 35
 64 EA 71 DE 6A D1 51 01 B8 C6 00 13 FE FF 4E 5B
 61 14 F1 37 08 27 09 96 1A 8E 68 E2 5E 64 12 15
 49 51 1B 12 D1 91 0A 1B 9C 1D 46 7F 4A B2 CF E3
 2E 65 12 AC 00 AA E3 7A B7 19 8D CF E5 93 C2 E2
 B3 EC 57 F2 BA 20 70 28 CF 77 DA 25 EB 9C E2 EA
 9C 5A FD B6 AD 0D 53 A8 4B FA 6D 51 D3 D2 B7 11
 E9 6E 89 B0 F2 BC 8A 34 C8 97 E0 40 B8 BC 8B 5C
 6C 5C EC 43 65 06 84 D4 E5 DC 91 D3 12 E0 5F C5
 7F 79 CA 7B 33 9F 0A 83 C9 03 4E 39 A9 46 51 1E
 6F 03 BB 10 DA 51 1C 92 0F F7 BC 41 CB C4 F2 89
 17 CC 1E C9 FC F9 DB 98 06 D7 12 12 0E 8A 7F C5
 A8 A6 82 92 03 E1 64 7B 74 68 70 6D 9F A2 44 C0
 70 AF 87 B8 61 F2 CB 57 84 1D 60 75 87 B3 90 C3
 FC BC DB FE AD 28 38 6D 88 19 B3 87 FB 98 89 0C
 60 BD 11 53 02 BD 01 D5 0D 26 9F A2 DA 33 CA 29
 95 0D EC 24 DE 8D 60 09 EA 94 19 77 7E 72 57 CA
 A4 83 72 30 10 D9 B6 5B D1 9A 2B F4 75 C1 21 84
 A4 6B 84 A8 EB 70 E3 0F 8F E1 11 24 93 50 1E 32
 80 32 42 A6 98 B5 D6 27 2F 06 B6 C2 36 85 08 7D
 C1 37 DD FA 3A A4 AA C9 2E 8B 90 AB 70 58 C8 92
 F7 96 C6 F5 FD 8E C9 F5 CA 8E 07 56 20 D9 FC BD
 A5 5F 06 60 5C 14 4E 31 28 EE 57 70 FF 6C 9F 5B
 AD A8 BC C8 BD E0 F4 F0 57 FC 9A 4F E4 54 6F BA
 FD 88 BC 93 9B 18 5F 10 EB A4 E9 BD 14 98 E1 C6
 74 17 66 56 20 15 37 C5 B1 6D 77 C2 E1 AF C2 DD
 57 6E DB D7 F8 F4 16 35 22 31 18 1D A8 3F 13 80
 36 78 2A D4 1B BE 69 CF 40 2F 1F A0 A6 2F 80 B1
 7A F6 E8 C5 31 C1 01 2F 24 39 B9 91 CE EA D9 D1
 DA C4 89 D5 0B 91 84 31 89 4F 82 08 1A 7E EC 1A
 7D F7 62 23 C1 C9 34 FE D3 FD 73 AE 4C 93 0B 1C
 4E C3 B3 D7 C0 70 A7 A3 31 09 1B D0 46 71 89 6D
 47 4A F1 C0 6F F8 5F 69 C2 7B C6 07 34 81 CF D1
 D9 B3 BC 7D DB 27 8D 89 29 5A 2B 21 7B C8 CC D4
 F9 8F D3 8A 90 90 FE 2A CA 58 46 3F 29 69 67 AD
 3D 24 CF E5 A6 9F 0D 18 72 A7 E2 26 8F 72 7C A5
 57 97 B4 2D C7 F9 03 4B 08 9A 00 3E 02 D5 55 D3
 63 C0 16 08 A8 22 E4 01 75 80 C8 88 E5 20 00 9C
 13 72 EE 75 3F 15 5B 18 57 EF A5 CF 6B 6A 21 CE
 E6 65 66 67 AC 10 10 0F 8E 7D 04 18 16 3A 29 2E
 2B C7 E1 C0 5C CD 7B AE 50 73 3D FA 5C 79 0D B7
 80 58 E5 3A 1C 2A 27 66 2D 10 A4 80 40 0D 20 FD
 58 8B 42 A2 2F 8F 7C E8 63 E2 75 EC 23 64 71 C6
 4A 70 2C A4 99 7C D8 6B FB 7B 12 22 77 38 45 17
 BC E3 45 0D CE 48 FA CD B5 AD C7 54 7C 2C 8F E7
 86 FB 17 85 06 49 F8 AA 4E FD 93 94 66 0D F6 8A
 57 75 3C 70 03 EF F1 1D 6E E6 03 65 46 39 BE 5C
 49 BD CC 80 E9 E8 22 EC 9B BF 24 43 B8 A2 C6 76
 C1 96 EA 60 9D 45 B1 83 4A A8 36 D0 CB 3F 32 E7
 D2 45 B0 81 E4 C7 68 9E AB BD 09 87 C8 AE 30 02
 3E 86 1C AE 0D 39 9A CF 07 33 37 41 FB 3D 7D 9A
 3F F0 AB BB 9D FD ED 36 2E 32 BE 3A C3 AF 8F F2
 68 CF 61 E8 14 9B FB AA A1 78 AD B8 BE 54 7A D5
 5B 58 07 03 A2 DD 17 BA BC 8D 55 FC 5C 90 0A 06
 EF 9B 56 C5 09 0D 9E AB 31 96 42 03 19 7D 9E 51
 56 80 20 BB A1 00 87 C8 F3 38 EC 25 98 4D 9C 1D
 13 70 04 06 98 31 CC A9 95 0D E8 AB 34 74 6D D8
 B7 4F CF 6C D4 8F DA FC 5D 11 0F 88 97 BB FE 0D
 EE AB C4 C3 19 2C 34 7A B3 32 77 93 F5 8F 27 C1
 7B 57 94 74 A4 EA 37 9D EA BD 4E EA 20 30 65 2D
 B3 06 FA A5 02 6E 8B 02 58 77 C9 12 6D 35 61 07
 3A F3 12 9A 0C 2A 7C 2A F1 40 87 D4 97 65 44 E2
 89 74 22 7E FE AA 2C F1 22 23 95 C9 0A D4 58 B7
 D1 A1 36 9C 50 51 45 DD 14 97 5A 0C D1 F4 7E 86
 F2 30 48 6A DD 09 3C B2 1E D8 C6 9F E1 99 16 6B
 53 19 32 5F 2F 5E 93 48 BF 9E 69 AA 5F 73 34 F4
 76 14 04 99 2C 61 CB 92 87 83 30 C9 A7 4D ED 3E
 9F 94 07 1B 92 2E 2A E4 71 C3 95 27 20 A0 C2 D3
 F1 F7 66 C9 F0 23 C5 77 3E A9 6D 37 99 09 18 FF
 BB AC 86 A2 4A DA FF 01 39 5B 4D F4 94 EF B5 0D
 77 AC 6A E9 41 2B 51 C0 D5 D2 1D B7 1E 15 C7 1C
 92 3D 76 4B E7 66 D8 6B 03 FE 27 8D 78 B6 FB B0
 7F 5C 92 35 69 14 5D B3 43 B4 A5 BE 9E 33 0D C4
 C9 3B E9 DA 4F 12 BE A2 C1 A3 A8 2D D4 00 FE A7
 15 92 97 C6 13 0D 2D 36 A3 0D C2 D5 EA 7F 2A CC
 44 A2 96 24 BD A8 6B 03 49 25 72 3D EE 6E 44 B7
 9F 56 5A A9 89 3A 3D 39 3A 61 52 1D 3F 52 97 8A
 98 CC A3 F6 BE 10 E6 CB 34 F3 EC AB DC A2 46 CE
 78 68 70 FE 76 C6 E5 3F 37 58 07 B2 84 F6 97 78
 13 BD 46 60 28 3C 9E C4 6B BE 18 65 75 16 C4 6A
 2A 21 C4 9C AF CD 50 F7 F3 9E 40 9C 6E 46 D6 B6
 6A B5 DF 41 6B 2B C6 C8 3D B4 0C DB A1 B2 ED C4
 79 42 E7 55 AE C5 31 A5 DE 82 70 F5 8A 9F 7D 77
 9D DE 86 29 9D 42 D4 75 9C 39 A7 06 50 5A FD EB
 08 CE 74 C9 D9 CC 5A F4 BB 73 18 AE C1 AC 7A B9
 4D 30 4B 34 22 0E 8A 96 C5 8F C6 4E E6 ED E1 07
 AA 2A BE 15 09 0D 20 DB 1B 69 8C 1D 8A 58 A7 AC
 A1 A8 38 37 CA 9B 17 D3 0F 9D 40 6E D0 21 CB 26
 E5 ED D2 65 D8 BC 98 A5 64 DF 37 B9 BA 4E F2 5D
 B6 A4 44 6F 96 D7 7B 7D 93 6E 0E BD EC F4 CE 53
 80 11 B2 E3 67 15 8A D7 A2 84 51 49 44 2C FC D7
 CB 85 74 BF A8 9E 75 6D 6F 9B 30 D3 3C 11 F0 66
 64 3D FB A0 93 30 BD A8 26 4E BF C6 E7 FC 45 3E
 EB 3D 2C 4C FA 41 72 C2 96 8C D0 B5 35 A8 14 A8
 34 7E 60 75 F0 1A 91 99 4A 2E 2C 78 EB 44 27 6E
 F6 C1 8D 9D 6E 6C 08 A3 4B 6B 6E 8C 93 A7 D5 1A
 6A 7F 3F 5A E0 82 BB 7E F2 CE E7 9A 04 F8 7E 7A
 E2 D9 B8 04 AE 2C 3E 6D 1B 08 0D A2 71 94 38 4B
 1B EC A5 78 58 6B 76 1A 1E 4A 25 F8 33 CE 62 D6
 9C 6A 68 98 C6 D8 40 AD 23 DC AA 30 EF A0 EE CA
 B7 6C 29 58 8F 0C B1 1E DF EE 6D AE 69 3C 24 6C
 B0 44 25 F6 FE B1 E5 E7 10 2E 2E B8 31 68 13 5A
 C5 C7 84 AE 5E 80 A3 9C BF 5B 6D 50 6B 2A 4E 9D
 E8 F5 40 B3 D2 BE 95 3B FC 58 7F D5 CC 20 61 23
 18 53 88 7F CC F1 EB D7 A7 14 87 97 12 96 28 98
 20 68 0C 6D DA AC 3F 8B E6 D4 F4 BC 12 61 7F 32
 15 2E EB 46 E1 D6 33 25 10 0A F5 AB 7B 34 CC DD
 A9 E7 9F 8D F7 9A 25 7A 42 EB 60 22 86 9E 8F F7
 13 95 67 D6 E5 E9 61 23 BB 96 89 0F 4F 62 D7 74
 97 DE A9 07 E2 E4 D9 62 7C EC 02 31 92 BB CC FC
 DB 21 48 67 77 5A DB 7C 7E 7A 39 DA 02 DA 04 77
 40 34 95 EE 13 FA 61 E7 79 93 4F 10 FA E9 94 B2
 32 09 C9 13 B7 81 B8 DC AF 9A 06 36 81 5B 58 29
 95 AF D8 17 37 C4 FB 1B 3D C0 0B 59 98 43 50 04
 18 C8 A9 FF CA CB 9A 27 E0 C4 BC D9 89 76 34 52
 EA E6 A2 41 47 3F 73 A2 E5 68 1F A0 64 43 D6 AC
 13 C3 AE 2C CB 75 9A E8 EF 54 04 8D 5D A0 E5 31
 B0 4A 58 B9 39 4E 85 90 BA AE C8 71 34 56 CC 7F
 69 CB 43 F6 46 69 14 E7 58 EA E5 D9 DF 30 CE 77
 D3 B5 CE 2E 7E 67 61 47 09 45 63 A4 2F 1D 3C 42
 F6 3E 23 C4 FF 81 DC 79 81 7E 92 55 33 EF 47 A4
 A8 0F 59 9C FA 0F 65 AA 32 11 9C D1 2B C3 DC 6B
 96 7A 0F 92 A2 41 28 4D B7 A1 F9 D8 2D 59 89 94
 CA B4 72 7C EA 1B 3A 51 69 43 0D D2 A8 23 A1 D3
 3D 76 B3 25 B3 6D 45 4F AD 82 01 B9 F0 96 A8 80
 79 46 4B 32 F1 0C F8 6F 6C 20 BF 6D E7 D8 A3 12
 26 5D 71 D5 96 E5 FA 76 3F 92 EB 69 CD 9C 0F B1
 97 84 28 0C 20 F3 7F E0 EA DB 20 44 DE A8 0A ED
 C6 77 B7 B1 0A 9C 3E E9 3A 35 01 D5 08 5C F9 29
 C4 9C FD CB 96 F2 92 50 A3 7B C3 5E AC E5 AB CB
 34 6F 50 38 3E B7 34 45 62 13 4C A1 B8 CC D9 E2
 5D 26 C4 10 BE 44 EE 16 AF 46 E5 74 2C 6D 7C 2B
 B8 43 5E 49 CC 67 1F 48 47 86 60 A8 80 AF 5E 43
 CE 07 A4 89 2E D1 9D F4 94 B6 C3 6D 84 62 D8 F0
 D6 72 9F 0D A6 6A 9F AA B6 91 FC 15 A3 45 A0 A4
 72 FD F2 F3 03 31 13 CF B1 24 6D 13 C0 5C A1 2B
 88 64 C5 2F FB D0 82 60 81 A1 A1 1A CA D8 CF 9F
 9E ED FF FD C5 02 ED F7 DB C8 5D 79 F6 4E BA 11
 17 15 52 D3 BF 5F A9 57 D9 E2 67 26 92 45 F4 E7
 56 D4 2B 09 7F 5B 55 1B 77 C4 93 6C 64 46 FC BF
 8D 30 9D B8 A7 9C 23 CD 88 3B 9B 25 B5 3D C2 74
 F5 06 96 02 7F 71 66 35 7A F1 45 C0 49 DD 46 F0
 32 19 67 4E 73 08 4D F0 CB E1 98 D6 D7 07 E0 F0
 B8 AF D5 DF 09 6E 36 2C 14 32 BC 96 32 F5 75 38
 1C C3 F6 1A C1 13 B6 46 9D D4 55 4C 5E B8 4C D5
 50 6C A3 30 E9 EC 87 32 3A 91 33 86 4D A0 00 24
 7B B8 67 C7 23 D7 27 EA FB FD 40 03 D9 73 CE 17
 F9 B0 10 0E 71 B0 1D B3 DE BF E9 9F 4C AC CC 6F
 15 1C 63 63 30 4C D1 09 58 4C 5A 06 40 96 69 9D
 04 FB DA 52 68 67 63 4A 9A A6 7B 65 8B E9 CA 5B
 44 E7 34 A8 0D C3 43 48 11 A4 84 30 34 0B A1 AE
 84 C5 68 76 7D D2 BE 01 75 CA 8B 49 B2 0B 8C 8A
 63 8C 0D 1B 98 E4 D6 37 67 03 24 90 4C 54 70 8B
 DA 94 A9 35 96 6D C6 E3 A3 1B 17 0A B8 CE E7 6E
 58 D8 90 2D 3C 2D 32 B5 9F 94 12 08 41 E3 C6 4B
 86 25 B0 F8 16 3C 56 22 76 1E 53 FD 91 DA 87 2A
 CD 46 5F B2 4A 4E AB 6F 64 72 82 7A 5D D4 C1 86
 F4 22 D8 A4 BB BE 59 87 DC D9 8B 0D F0 F0 A5 F3
 22 B7 13 16 51 9F FE 93 C4 E5 93 56 83 3A AB 60
 B2 E5 85 5C BB D1 44 1C 78 EE 60 13 5F 7C 32 11
 81 5F 52 7D 58 45 50 97 12 C4 7E B0 F0 75 86 21
 29 34 2D B0 EC 90 AB 0F A2 19 28 4C 82 40 17 BD
 A3 EE 88 A2 ED 3A B3 73 E2 D9 7C F3 DD 16 95 1B
 C4 F3 B7 4A 2A 9E 3A 90 3E C7 68 FF 4A B5 4E FD
 E9 F5 F3 46 53 12 6D 87 99 F1 6A BF 28 0D BC D2
 06 A9 23 B4 3C B7 98 A7 4F 05 64 D2 BB 55 79 0C
 69 11 75 92 D3 1A 7E 80 E5 E1 BF 40 71 BE 9D 8B
 E6 2A 2F D0 B7 6F 25 77 61 BD BD 8A C4 A1 C4 3C
 9D BE E6 DA 24 DA 8E CE C9 00 2D 1F DB 85 AA F5
 38 9E 47 96 8A FB 32 06 6C B4 B0 3A 03 E6 B4 6E
 99 5E 72 5D 73 7E 92 6C 7A DC D0 94 98 4D B4 46
 44 CD ED E8 EC 0E 5C 64 F3 05 1E D0 A9 F5 46 BB
 07 31 59 57 84 35 0E A2 17 44 08 96 FA 49 40 26
 C2 13 57 AA 81 AA 12 67 63 18 F4 D0 0E A0 4F 54
 2A 05 0B B9 3A 55 0B D4 E2 AC C3 0C 7F 73 0A 4E
 FC 00 06 56 9F D4 B3 43 72 4A 29 D7 DD 00 35 9A
 B0 82 1A 2D 67 7E 53 FE 59 61 87 73 85 41 BB D8
 53 3D D8 26 F5 73 98 A3 92 E6 AA E8 3F AE 3B A0
 C6 B2 14 10 45 DE 0B 27 B3 4D 73 AF 88 F5 A9 BB
 84 89 CD E9 D0 D3 31 E6 B1 CB AB 15 13 13 F5 EA
 FA 37 21 3C AC 60 61 A2 89 2B FD 07 8E 27 5D 67
 43 9E BB 58 12 74 09 B8 1E 61 65 57 86 0A A7 4A
 52 9E 87 A0 8B 35 AF 41 77 0B B1 0B A8 96 04 4C
 C0 1A 06 E4 85 89 4E 2C 27 DD 07 F1 2B FB 93 AF
 66 25 BE 4E F4 1B BA 24 66 86 FA CB 44 F9 B6 40
 69 AB 46 9E D0 B2 FD CE A5 78 52 97 1C E9 E0 B8
 97 4B A2 B8 34 B7 90 9F B3 99 2D 63 E6 1F 77 A6
 F3 92 DA 64 EF 30 5C 53 43 AB 7C 1D 78 B5 83 03
 C2 0C 65 D6 67 21 B6 7E 90 12 E1 62 F0 DD 2C F0
 3D FC 1F 92 59 D9 EA C5 CD 33 97 47 54 56 C5 68
 2E 85 00 03 CC BE 12 29 CD 7A F6 D6 CF FE 02 B0
 27 9E 3F E0 E6 19 7D 27 B5 ED FE DD 7A 5B 4B F6
 B7 72 25 78 DF 3E 30 A5 DD 4D E3 07 B7 38 7D 15
 68 CA EA 79 C5 39 A0 DE 8F 38 95 62 86 33 0C 98
 7C 9F 20 33 44 3C 22 77 C0 F9 BB 67 D9 FE 40 37
 FE C3 FE C4 B1 E9 0B 56 74 8F 69 A0 37 22 62 C4
 E9 5D E6 15 FF 58 1A 64 F7 03 19 AE 84 1A 00 7E
 85 88 DE C1 07 72 F6 1C 35 92 8E 20 D0 AF 32 0C
 ED 3C 50 FA 54 46 80 BD E7 51 42 40 9B E5 FC 2E
 8B F5 F1 15 9D 1D 59 C8 21 AD 77 4E EB 0A 60 85
 0E 9F 0B 88 B1 26 88 B1 17 B3 46 EF DB 2D E1 CC
 5F 13 5C 4C BE A0 50 FF 8A 62 34 94 3E 4C 22 08
 90 28 85 26 D7 C7 DA 19 1E 38 0C 3D 65 76 A0 44
 80 09 4C 49 9D 95 22 CE 1D 32 E1 6A B9 07 50 11
 C4 6D FA C0 C9 F1 F5 59 88 F7 90 3A 66 96 C5 69
 A4 70 B0 05 41 97 12 C4 02 E9 44 8B 5E 27 BB D3
 88 66 A8 58 DA 53 62 9E 71 FA 35 F4 DE D7 20 58
 79 3A 4A 7F D0 5B 9C 11 4F 6E BA 28 24 97 DF D0
 9B 7D 8A AA EE DC 16 6B B8 B6 D8 D6 87 1B DE 8A
 1C FC 4B 5F 5E 5A CC D5 09 0E FE D7 5B 76 40 81
 88 15 E6 96 40 F2 C9 68 52 F6 6B EA C2 42 84 9C
 39 0E BD 9A 63 66 6F A2 EA A9 94 94 A9 FB 13 6D
 68 E1 77 A6 B5 A4 94 27 D6 37 0E 16 C9 11 8D 5F
 CE 89 44 A4 AE DF A0 F5 44 87 B9 B9 37 D0 B1 6F
 E0 59 39 EC 9B CE 00 CE AD 1B 1A EB 17 0F 8A A5
 DE D0 B0 02 AA 80 2F 91 06 8C D0 92 D5 EF 0B 73
 05 F0 7F AD D7 2F 24 6C FD 2E 2A 10 93 34 CC A0
 AC C0 11 24 C5 AA DD 5A 01 ED F1 33 24 F4 BE 01
 11 B1 42 58 4E D5 E0 31 23 B5 19 6A 7F F2 F6 68
 01 25 C7 8D 8E 98 9D 0A C7 92 68 84 AF D9 2A 29
 47 53 0B 0F AA AF 13 88 E0 A0 90 1A 41 9D 65 7C
 01 37 02 08 78 BB 10 87 4A 36 8B D3 C0 5B D1 3E
 E8 8B 74 BF F2 AD 12 EF 81 2E E5 5E E9 41 6D B7
 EC C6 E5 22 3B 69 D7 FD 2C 82 B5 85 10 84 4D E0
 1F DF 4C A9 B2 70 86 03 93 4D 8B D4 AE 3F DF 90
 93 87 98 B2 5A 7D BF 5D 8F 52 65 27 48 EF 74 25
 F6 54 74 37 8F 7E 5A 2E A1 67 19 2D E4 6F 50 09
 B6 D7 9C FF 7A 60 4E B8 4E 7C B7 25 8A DD 0C EE
 B7 C7 10 0F AB F0 91 6B C9 A6 25 C6 4E 5F 5D E9
 5F A8 F1 3C CE 6A DD 4B B6 AA DB E9 6B E3 2A EF
 C5 4C C4 25 44 BA C6 E6 64 DA DF DE 05 39 DF CB
 F6 6A 66 65 C0 F4 CF 87 42 81 25 F8 CA E4 D1 FB
 CB 16 DB 30 30 90 17 F2 6A CC F8 69 69 E0 25 56
 58 3C F1 27 89 61 EB 0A C3 99 C0 2E 63 C8 72 E0
 4A D4 C4 C5 B7 7F 0C 37 CA 30 7E 61 0A E9 50 15
 B0 E0 17 06 CC 8D 2D 85 1B 03 E7 54 A1 B7 CB BF
 BF 50 BB 62 AA 1C F7 C7 1C 59 40 F3 79 DF C7 3F
 17 A1 51 05 74 7A 27 F7 CC D5 9B 10 29 56 1F B4
 A6 E5 E4 A8 F0 A5 89 6B E4 43 8B 80 3E 4E AF 61
 0E 71 B5 18 9A B0 C3 8C FC 21 00 5C 87 05 68 5B
 5C D6 90 FF 62 D7 40 A0 84 08 AB B1 24 0A 73 BC
 2E 0C 1B 6B 21 F4 69 0F B1 4C EC B2 CA C6 CF 62
 2C 5D 5F 73 81 56 56 1A 80 60 4D 2F 5D D7 F3 D9
 6D 0F E7 B0 92 FE 6A 63 1D 13 E0 15 5D BB 9C 36
 88 9C A1 C4 DC 79 F4 BF 69 E4 D4 A2 1E A3 5B 73
 44 20 5B E3 B5 A8 2A A9 62 F6 E0 A7 02 C9 2B A3
 6B 2D 1B AF 2B 22 41 F6 D6 12 75 0D 49 7B A4 8D
 20 DE B9 12 67 EF BA CC B4 77 80 59 DA C5 C1 10
 55 FC E5 38 F8 99 46 2A 15 36 06 A4 34 7B F2 17
 5A 70 6B 35 4F A6 95 D1 06 AA 3A 6C A5 E8 5F D1
 5B 2F 88 A0 35 48 6D D3 D4 8A AA EA A0 91 C8 C6
 2F 0F 9E 6C 13 5E 80 92 7D B2 98 AF 3A 5C CF 07
 AC 15 BF 37 25 15 BD DC 3C EF 84 D5 EA 1D 25 C0
 9E FC 73 90 D7 E8 B4 DF 58 66 8B 09 D1 FF B7 A5
 54 13 99 A9 0B 50 07 D5 0D 05 C2 ED 0B 00 32 F3
 EE 0D 3B 69 09 91 AD 4A E8 95 5F 23 C4 10 F5 F8
 3F 06 B4 46 B9 E9 8F D9 35 8F 69 93 8B E4 EA 76
 2A FC 02 0D 72 38 9F 4C 37 93 B7 3C F1 AC F5 7D
 3D 5C 54 9B C2 51 B6 A5 64 51 CD 02 BD 36 88 9B
 22 09 AC 02 D9 DC AE 7F DC 3F 00 0A FE 67 1E C7
 35 B9 68 E8 C6 31 39 1C 3B 0F 9F 57 42 3C 12 5E
 45 0F E3 73 49 62 46 32 E2 1C 5C 4C B2 1E F4 31
 94 FF FB 26 9A 90 D0 DF 2C B2 33 2A 7A F2 4E E1
 EB DF D6 D3 0F A6 DA 16 1E 67 3E DE E4 99 94 00
 36 C8 69 0A 7C 75 70 B5 6A 4C 2E 3C DE 1E 09 5E
 83 17 29 D4 D5 A0 78 BA 54 54 A2 4F 12 28 FC 8B
 D5 B0 5F 10 3C DA 1F 57 B9 8D 92 60 57 F1 44 08
 DE 24 78 EE D8 CC 86 97 8C DA 05 FA 30 D7 0A 1E
 70 86 3D 93 E3 C5 74 6D 77 44 81 69 3A F2 98 A8
 6F 82 44 4B 3C AA CA 76 D8 4D 29 21 70 E1 96 5C
 EB 06 76 2D D4 58 21 B0 64 55 E5 FC 9B 96 72 95
 9A D2 CE 92 3C B5 7E DE 2A 35 42 10 A8 D3 EB EA
 2B 89 CA 09 19 4B BC 96 02 42 31 D8 4A 69 78 68
 9B 22 84 AE 6E B2 32 70 44 AF 32 38 88 B8 10 97
 83 83 7F 34 6E 03 13 70 36 70 BC 88 F6 D6 CE 97
 AF 7E 59 4D 88 05 3B 72 3D 96 92 27 D2 C0 DD 17
 1C C4 0F 62 B0 70 72 DD BF 79 24 A7 A3 C2 12 29
 A4 DA 47 33 37 36 E3 C3 08 93 1D BE 12 B3 21 6F
 0C 9C C8 91 27 AA ED 02 38 0D 39 26 3D D8 67 26
 CF B6 E3 34 8E D4 E1 4D 2D 78 53 17 E5 9A 6B AA
 28 64 44 DA 62 6C 4B AC 51 9D 04 5E 41 4A 46 74
 14 6A 31 F9 2A 26 6A 89 A9 76 13 11 C9 D7 34 42
 14 67 2A 1B 46 D1 70 03 B9 58 50 EE 39 9A 08 68
 41 06 77 FE 7B CD D0 19 C3 3B 1A 7F A7 EF D7 5B
 38 B5 60 12 9B A1 95 54 EF 58 CF 91 EE D2 42 F8
 7C AD 94 C2 0C 6A B5 C6 35 A4 63 A2 E8 1C CF 14
 11 C1 F7 C9 DA 1A 81 4A 40 F7 16 B9 25 EE 68 AA
 75 FE 57 5A 74 32 BC 7C 3D 42 1E 1B ED A1 33 53
 C9 16 A4 59 26 DD 76 BC 11 27 A1 A5 F5 B3 FE 50
 12 23 B0 2E A8 39 37 42 1C 0A C3 7F E3 53 0B 51
 A2 43 61 00 4B 06 F0 C8 57 BB D4 E2 F9 30 6D 98
 21 1F 08 23 19 E7 2B 7F 6E 98 DF A3 39 6F B5 30
 99 C3 AB EC AF E9 12 1E D3 E8 59 16 2D 19 D9 80
 AF 8D 94 EF 26 AC 1C 3C 40 33 F5 6E DF 5E 21 28
 8B AD 5B 7F 60 1D E8 B3 6F 58 66 D5 DF 6F 68 BE
 56 7E 5B 1C 57 7A 7A DE 60 46 93 CD 5D 02 C5 12
 39 DD E1 01 09 97 A7 7E 58 7C 8E 40 45 B2 89 9B
 46 67 09 0D 54 E6 CA AA 6C EE C8 70 41 37 34 69
 EE 78 85 FE 51 2D 8B 08 DE 5A 8A FF 70 CE D0 51
 20 59 08 1A F9 36 89 EC 94 71 4A B5 A3 5C A2 FB
 AA BE 5C A1 A0 32 70 D3 4C 67 45 D9 B3 D5 6D 91
 FE B0 EC 9B BA 75 C4 2B F5 16 37 E2 EB 0A CE 5B
 A7 7D E1 0A A2 FA 5C 27 03 E7 3D 29 37 78 01 25
 2A CD 63 06 2A 82 A5 BC 7A A3 C3 EC C7 11 92 45
 16 08 56 7B 49 09 0F 1F FA D2 68 7B 35 A2 C1 3F
 4F B3 A3 52 1B 51 A6 B9 3F 1B 2E 93 E0 59 F9 B5
 DA 72 FE BA D0 F5 F3 44 74 8B E9 00 B6 BD 3D B3
 7F 3C 7F 0D D7 BB D5 10 4A 50 0D C0 00 EE 30 86
 47 D3 1C F7 AF 92 F2 6F 8F BC D1 86 E9 AB 8A FE
 AA 8F 23 51 BB 65 D1 61 CD B0 59 DD A4 EE 6D 2C
 5D 03 13 E0 A2 AE 02 40 31 5E FB 77 F8 C1 4B 3C
 B9 AB B2 D3 61 C0 CD 7D AF EC 66 FD 1A FC E0 4D
 39 23 5C 50 51 BD 66 02 D1 ED 75 8A B7 A2 BF 2E
 7F A6 8D 28 7F 75 BF 20 43 88 88 90 71 25 78 6A
 ED DD 92 45 A5 25 8B 75 7F 59 98 33 77 4D 4C 84
 0D D2 27 A2 1B ED D7 DA 35 24 37 21 C4 20 66 98
 D4 90 FE 57 7D 65 D1 BC 32 62 38 B8 88 8C 5E 2C
 8E F8 DE 38 90 DE 30 3D 09 A8 27 8C D4 5E FA 8C
 CC 6A FA 03 48 EB 20 E8 C1 F5 F6 15 69 FC 76 0D
 FD 1A 52 4D 72 CD FD B0 8D 5D E8 37 89 61 1D B6
 C0 29 C6 6D 82 68 E4 B5 67 7C 7C 0A BD DB B5 82
 8C 50 42 33 3E 9B 84 5F A7 3A EE BE 65 BD F0 4B
 93 56 DA F4 27 8C 53 90 E5 A8 23 89 4F E7 E6 AB
 36 09 AE D2 69 90 15 BC 40 C7 00 45 37 0D 94 ED
 74 78 9E A6 7A 66 B2 FF 81 B7 DB 94 CE 28 30 E2
 81 25 E6 49 91 B1 FD 2E 02 CF 57 01 C2 0B 25 8E
 06 DB F0 C8 22 4F F4 C7 04 20 D6 18 FA 38 5C 63
 E3 71 C3 08 91 28 BB DE 6C CA 92 A6 1D DD AA 0B
 F0 AF F7 F0 05 9F F7 C5 F9 E3 56 EC 10 49 7F 3E
 CA BB 37 10 D8 CD B2 74 C2 3A 36 10 15 67 78 18
 D6 CE 3B 79 78 3B EF 3B 69 A1 8F 6D 1B B8 0A 9F
 30 B6 F3 54 43 5B ED 3B 42 0F 39 7E D7 64 16 AC
 B0 AD 20 82 77 36 F4 23 31 12 D7 0C 84 06 D1 E8
 11 71 9E A9 5F C4 BB 9C FA 0B A1 A4 78 8B 49 28
 10 B2 19 0D 87 79 47 16 E2 0E 2F 21 C5 AB 5A 57
 FF 90 76 3A 6D 12 BA 00 42 27 66 52 33 7C 50 12
 38 4E B0 5F BB C2 3E A4 B2 A0 3E A8 6C 58 8B FE
 9F 36 F2 A5 64 61 3B 6D 54 5B F9 CB 26 38 FC 5E
 D9 FA 26 E5 76 D8 90 63 1E 3B FA D0 A5 F1 27 F8
 98 6A 69 AA 11 F8 40 62 E5 C1 7F D5 61 31 2F C1
 66 A8 15 55 7A 2F EC D2 2F 60 24 84 77 72 90 09
 26 57 7F 9B 9C 74 83 13 F8 49 40 27 42 B4 16 84
 C8 FB DF 4D 6B 21 56 73 85 E4 B3 A1 42 B6 A6 67
 47 BB 95 05 3F D7 24 12 12 89 AF 08 87 E6 6E D5
 CA 11 19 A7 97 7A D3 4E DC 9C 36 DE 4C 64 2D 83
 79 EF 8B A7 11 08 98 9C D3 A2 24 4C D4 00 82 E9
 AF 8F 26 FB 69 46 85 B7 D2 A2 AA FF 8B FE 3C 66
 38 EE EB 39 3A 5B 9F 52 28 D8 6C 5F 7A B0 D5 6F
 F3 CC 55 20 17 9E 90 FD EF EB 9A D9 BF 74 74 07
 B9 6B 7B FB 96 8D 64 BD 2E DF 9F EA 87 2A A6 18
 01 3E E7 3F C0 66 96 BC F9 2C 1D AF CB 50 A8 4B
 A9 15 1A 2E 4F C3 FF A7 53 AA 0D 0C F5 04 95 F1
 E7 A0 6A E3 5C 92 3E F2 FA FE EF B0 01 2F C8 92
 05 E6 BA E7 5A 03 72 29 EC 93 78 E9 D8 D9 01 24
 DC 46 3A 05 74 1E 61 B1 74 28 CB 4A EE 94 76 1F
 4D 6E 12 76 53 B3 AE E6 99 A5 B2 95 D1 88 B6 29
 D3 52 42 AE AB FC 9B F8 B3 E9 DB FF 96 4C 69 E3
 3A 4A 81 A6 73 62 F5 AF 5F D8 CD 68 0D 52 89 F4
 0A E2 E9 57 E7 34 6B AA D8 44 D6 93 51 1E 82 F7
 85 E0 14 59 A0 56 91 A7 25 00 06 78 D4 40 BA 64
 82 D4 4F B0 B9 FF 58 CF 4B C0 48 E1 63 4F F0 3C
 CA 4B 8B DC 2C D1 2F 35 77 93 DA 17 50 A5 F0 24
 C1 21 D5 26 55 2A DC 37 44 A4 D9 5B FD E5 FD D8
 67 D7 CF C5 29 3E 71 B6 83 B8 84 86 A8 C1 B4 AE
 84 01 4A CC 5E B3 A6 F2 CE 68 76 B7 25 F9 F6 E6
 32 AB 69 EE A1 99 25 7D 3B 8D CE FB 24 6A 33 85
 9B A2 BD CC 3A 81 4E 8E D1 57 A3 DC 96 47 30 64
 74 39 7E 27 96 32 74 BA A7 E6 9C F8 5A 74 0B CB
 8A CF 39 23 EA 1B 08 8D A8 14 D2 8B F5 BE D8 E3
 F8 8F 98 27 69 11 7C FA 1C BC 69 99 B6 2A 3A 04
 A2 29 4A 0C BB 5D B6 BA 87 5D B9 FE 60 7F B4 2C
 D4 B0 14 FF 90 DB 82 BC B5 EA 81 5F 90 35 F1 2A
 A5 48 B7 C6 63 56 62 4E 1F DD 4F 4A B6 16 A6 EA
 AB 96 5F 94 6A 51 CB F7 64 D7 3F 96 E8 99 97 F7
 A1 26 DD D3 2B 47 CB CC AC 62 27 32 92 43 DA ED
 E6 2F CE 7A 7B 53 01 CA 5B 40 8A 08 6D 67 FA 83
 0D E2 E2 83 72 21 1C 35 C2 52 45 71 E7 5E 67 D8
 C7 36 D4 79 BD 44 D7 69 7C BB 9A 3F F7 1A 98 CA
 B5 42 37 01 18 E1 A1 27 57 84 7B A7 21 F6 64 7E
 9C 3F CD D2 D1 00 17 E4 95 E9 27 0B 00 4E 2B 45
 95 3E 90 CD F7 70 B0 7C 97 9A 6C 80 AF B5 2B 6A
 8D 19 A8 BB A7 D3 49 04 15 76 C0 C7 1D 89 4A B7
 7E B5 4F 35 F9 94 9E 2F B5 66 4F 3A 45 51 1C D3
 3F 3D 25 E5 4A DE 31 89 3A AA 7D 18 05 61 15 C5
 73 DB 59 FF F0 06 C0 D1 AA 6D C9 2B 71 28 AE D3
 37 39 8E A8 55 05 A6 3E C9 47 A4 C8 F7 24 C7 34
 D1 34 9C 4B 03 F3 5E 73 A8 18 A5 E4 FA EE 5A 6E
 62 3E CF A3 BA F2 AE 62 C5 28 BC 51 7E 9B FE BA
 68 64 E1 A7 E9 8C 3E 04 8C DA 3E AF EE B2 C2 D8
 86 8F F1 DD 33 24 70 42 F0 3A 27 31 F7 39 05 73
 2D 5B D8 B2 09 A2 8E B1 FB 67 91 69 88 19 D7 2F
 44 AF 55 2C 37 66 C1 4D EA 7D E3 D1 59 60 F9 60
 39 FC 39 BC AC C1 7D 30 1D BB 9F BE 0D 42 ED 28
 98 CE 8E 93 99 C1 E5 E2 80 2C 0F F3 C1 9F 28 2D
 D4 EA 19 58 55 B3 25 89 C4 D4 7E D2 12 A3 60 70
 D0 1E 42 C2 04 E4 34 39 12 38 28 D7 0C B7 9E D9
 E6 5D 4D 31 94 6B 0D 3B 3B C6 53 41 53 96 79 A3
 C9 74 6E 83 45 62 75 B2 4C 8E E6 B9 09 8D B7 9D
 9C DE 6C 54 05 A7 60 9E 78 93 96 F0 FE 61 02 B0
 27 0C 8C 03 E8 55 AC 00 D4 81 83 C5 05 A6 23 75
 E2 DD A8 97 F2 2F 8A B4 75 85 37 B2 6B CD 73 73
 D6 5E 67 EC 56 DD 5D 36 AD 38 A3 5E BB A4 41 6E
 4F 76 95 04 0B A0 82 E0 9B EB 9F 6E DA 87 AD 90
 E6 45 C0 E3 7A 9C 0B E0 48 9E C4 C9 5C C0 4B 00
 96 C0 44 8D E8 D4 E5 65 15 4C B7 C1 B0 DF 9B 67
 2A D2 63 0F C1 33 50 8A 88 0D 5F CC D8 68 4A 2B
 9E 70 EA 69 4A 55 34 02 E1 59 C9 66 6A 8E 39 74
 9B E6 BC 56 28 2F 65 42 8A 82 D5 2D 53 7A F3 94
 B5 48 40 5C 7F D2 77 67 1E 51 FA FD 3A 45 AD 8A
 E2 BB 1B AA 29 B2 34 F0 D3 49 BA 8F 4B A9 16 5B
 35 B8 C6 91 66 7C 04 7E F8 E5 73 0F 90 7B 98 7F
 04 F0 89 78 CE CA 92 4F A6 79 C2 C6 AD 7F 1D 17
 8D 4D 8E 77 68 59 6A 4F 88 19 2F 77 DA 90 F8 8E
 14 D3 F1 FF B3 23 9D C5 8D 25 B7 24 2A 30 6D 49
 A6 D7 BB 02 A1 59 CC CA 57 25 47 74 E5 E5 70 98
 B0 4C 87 0E D3 BC 22 21 92 FD 2E F7 8B 7A ED 21
 2D BB E8 71 81 CA 21 6D 5C 6C A3 8C 4D 3D 47 03
 82 98 FF 85 2C 55 E5 61 C1 B8 A5 2D C4 AA F5 2A
 7D 16 63 98 C6 C3 5B C6 A7 6E 3A 5C CE B2 1A EE
 16 7C 06 F1 A5 5E 12 32 C8 89 83 0B F6 1A C9 01
 77 13 EF 6B 53 8B 79 C5 4B 89 F0 19 C9 0E 89 84
 89 40 B6 40 56 67 5F A9 2C 2A 46 E4 7D 5E D4 0F
 17 2B B5 7A 34 79 CB 2A 09 41 09 A4 85 99 10 9F
 42 0E 14 98 66 17 6B DB 46 D9 04 EC 83 54 CF 06
 CB DB 3B 11 C8 EB 39 9A DE 99 95 52 8C EA B5 78
 EC 61 8B 1A CC 77 03 26 0B 73 D8 C4 61 68 84 20
 93 42 7A 44 17 25 0B FD 5C 80 CF 59 84 19 52 28
 1B 06 B4 9D 9D 43 AA E5 95 AA D8 8A 0E 38 D9 8D
 E5 BB 9D AB 5C 3B 64 40 25 BB 77 2C C1 C5 F4 33
 2D 1A A8 53 CF 8E 2E 77 40 26 D0 92 CB E6 38 98
 33 94 7D 41 2A F9 FE 23 F4 D8 5C 16 7D C1 8C EA
 E4 8C 06 A9 A4 C2 D2 14 2B 90 79 B4 31 74 CA EA
 12 A2 B8 55 BF 0E 47 C2 3A 12 D4 D8 BC E6 19 2F
 D0 D9 91 65 06 38 6F 54 D9 FB 56 12 EA B9 43 C8
 48 FA 17 C7 24 DF B4 8B 29 FE AB AD 65 23 DE DD
 85 E2 1A 19 48 99 75 E5 74 87 45 C3 21 89 DF 1D
 B0 19 51 46 29 4F B4 67 5D C6 59 F1 08 29 3C CF
 B6 7C 56 DF A7 30 7B 11 FD 6F 05 E1 EF A6 57 22
 91 B8 EF A6 9D D5 E1 22 96 E9 70 FC BD F1 F5 51
 E0 8B A2 DF 28 2A 96 61 E1 04 77 56 DA BD D0 A4
 0C DA 0D 6D E3 B6 03 C0 67 6F 24 DC 4E 5E 89 53
 92 BC D6 CC 28 F7 24 64 7C 6A D4 2F 28 A1 FE 45
 2C 3F 51 E7 D3 F2 BC CA 25 41 4D E2 02 01 C6 BB
 C3 3A 3F 95 EE 5F DF FC 04 27 56 B1 89 95 46 6C
 77 F0 B3 D9 29 70 26 82 FB 60 F4 BE E7 94 1D D3
 1B 3A 80 53 99 61 66 28 6D BE 47 8B BC B4 3D AD
 96 0C C6 79 B6 A8 27 39 7A 3E 86 F2 0B 24 96 88
 BF 8A 9E ED B3 40 FB 74 5D E0 58 1B 3C A2 49 29
 7D DB 27 63 26 C9 47 EE 6F 8C 29 AF CA C3 3D F6
 F8 96 E3 7F AE 35 50 2D A1 78 03 1C 6E 1D 61 7D
 3F 17 49 A1 29 77 72 F8 B6 B0 1B 5A 00 17 BA 34
 CE 6A 8D 27 D1 CF CC BB 34 67 F5 85 E4 8A 53 DB
 04 23 91 0F B4 D1 BC 64 7B 3B B1 2E A4 66 88 DE
 93 7C EF 3F B4 48 D4 49 A0 85 9E 01 F2 FA B1 D6
 43 EA DF FF 96 B1 C2 C2 80 DF 88 06 BB B0 94 4D
 D5 CB 28 66 2C 4E 93 52 6E AF B9 EF 24 8F FC D9
 2F 62 E7 A0 E0 6E EE 7C 52 CF 55 68 D7 25 FC 63
 9E 78 7B 6D 13 FB A7 36 CA 8B A1 B5 93 DD 39 30
 01 1C 16 DD 5D B8 0A 14 BC B9 21 C6 DE D8 C2 62
 62 AC 7C CA EE 2B F0 4B 43 BC 06 AF 8A C9 DB FA
 20 AE 48 DB 32 B4 BA D6 5B 0C 9F 4B 55 EB D1 3B
 30 19 DA CE AD 71 42 A3 34 A4 1C DA E3 05 1F 4C
 14 A2 12 A1 7B 9F 4E AE E7 71 27 7B 6D 6A D5 E2
 D1 35 E1 DD 2F 6C AA F7 5D 29 9A A2 09 B0 75 CB
 E5 99 3A C5 27 51 25 C7 5E 60 D1 6C 53 A0 80 F2
 C3 2D 44 BA 50 0C 16 B6 5A 5C A2 22 A4 9B 24 29
 D9 21 26 D6 8E 16 8B B1 EE 75 81 E4 C6 9C 9B 75
 80 19 8F 55 AB CC E5 05 4A AA 0A 12 F1 D8 1A 39
 03 90 19 07 C7 53 AD 29 11 FF 86 14 73 D7 08 D4
 04 1E A8 F2 9D 7C D8 06 71 9B C0 C0 1A 65 0A E2
 67 6B 9D B0 14 D2 F8 0B 6B F7 6B E5 4C 8F E6 86
 EF F9 0F F4 62 5E 22 9A 81 F1 0D BD FE 65 C5 8C
 EA B1 20 22 67 B5 62 FE FB 32 C9 D4 D8 11 F3 94
 A9 3C 47 01 84 B8 B0 73 56 37 7B CA FB 83 F8 A8
 AC 7D 0A 4B 7C A0 39 F5 02 DA 0B 94 DC A2 F5 8B
 A3 1D D9 BB 3E 38 43 CC 8C FD 9D 2E 8C D9 C2 84
 D0 08 F2 7E 8F D8 E7 3B 28 A1 4D 4F 33 BB 86 E5
 AB 01 CB D3 AF 13 0D 3F 99 67 72 DA 72 68 3D 8A
 85 49 EB A4 D9 39 EE 66 7C 2D 5E E5 33 A3 5B C2
 DF 98 12 74 FB 05 9A 9C 31 2C C2 4D F2 C7 70 07
 1A 9E 3F 07 FC D6 4F 68 9E AF 81 B5 3D 46 E8 EF
 70 97 97 34 85 C1 59 FA F6 DC D4 F7 A6 0F 7B E2
 FF 25 BE AF 66 AF 4A E1 D1 B6 C1 7B D6 5E 62 42
 FC 90 11 03 4E A5 D6 B2 32 08 D3 33 C8 5D A7 5C
 A2 0E FD 1A 0B 57 A0 9A 28 37 B5 5B D0 2B BF 2E
 EF 62 22 FC 8F 5E 02 CE E4 16 34 AB 4E 43 D0 53
 C6 3B 2B 0C 15 64 AF 50 79 B4 7E D7 6E 3C AD BE
 13 0F 97 08 C1 24 B8 6A 4B 4A 84 0D 78 A4 72 B0
 4E 56 4F 7B C0 E3 00 EF 92 8B EC 6B 64 8F CC E9
 1B 5F 22 D3 34 B2 60 F8 8C 75 52 D5 DF C3 6E EE
 42 9E 52 CC 2F E4 AA 2F E5 64 25 BB 9B D6 B1 95
 49 81 49 91 25 E9 81 F0 92 C5 8A 9B 73 A7 EC 1E
 AC 0C 37 49 78 C8 F6 12 18 67 D1 D4 7C 61 A1 C2
 BE 36 22 52 0F E5 30 E7 36 2B 9E C1 FF 28 20 0B
 FD 2B A8 DF 1A 07 E4 57 E7 B1 A2 9A 4F 06 74 38
 64 19 4D 45 C5 07 40 D7 CE 8A C1 BE 60 A9 05 71
 17 39 D3 D9 43 F3 2C 2F CF DD 6C CF 73 A8 6D A7
 C5 7A DD C7 92 4C D7 C7 50 47 3D 2E F7 1C D9 10
 AA 21 62 1A A2 77 3C 29 C5 C6 BA 6D B9 88 B7 89
 F7 89 81 73 56 FA 4A 4D 14 7F 96 BA 0B AE 9A 93
 2F D9 07 56 54 C1 51 57 C0 75 DE 1E 5E 54 99 68
 7B 8B F7 38 09 17 BA 49 DB 23 62 04 B6 F9 12 4F
 E0 DE CB 98 8D 48 0B 52 00 88 F0 E3 5A 5D 3D 79
 A8 5E 41 58 BA 67 E6 86 12 77 C5 6C B1 62 7F DD
 FE 1F 75 53 63 AE FF 8E 01 08 1B DF F9 CE 5F 35
 EB FC 7E 06 22 3E 24 FF 12 79 FB E5 B4 4F 2C 4D
 6F C4 2E E2 55 63 C3 82 BC D5 3E EC DE DB 49 C5
 A5 8C B5 F7 E7 04 35 42 94 74 57 72 DF F9 D7 FF
 B0 16 EA 69 D1 A3 A5 35 F4 0C 66 14 99 16 94 7F
 0E C0 4B A4 81 DD C0 61 F3 3C 3B 02 9A 26 5D 28
 61 D3 19 AF A0 FF 45 CD F3 3E CB 7C 95 CC 06 3E
 AD 07 01 8C 40 9A E9 1D E7 2F 55 71 9D B4 35 2A
 E6 5C 92 31 AD EF C1 2C BF E4 1D 39 0B 21 52 9E
 FA 3F A3 04 D4 B4 39 14 64 51 AD 6E BD 35 9E 7A
 31 AF 24 3A 8E 3C 78 47 B3 B9 84 C5 9A 15 99 EB
 5B 77 F0 98 F5 41 3A 7E D8 9D 10 62 07 03 7B C2
 26 A1 65 FD BE 3C 65 D3 4D DB 9D A1 F7 1C A9 6B
 AB 83 5F 8B 69 C6 43 C6 39 E0 0F 49 EF E7 3D DA
 79 90 30 CC 56 12 B0 6B 09 B1 65 33 4D 82 89 9D
 C8 2D 59 9C 65 E7 F8 64 36 CB 26 EF 9F 09 6A F6
 DD A9 8C B1 4C 27 E3 26 4C 4B C7 7B 3E C6 CE 34
 10 6E C0 5F D9 C0 85 31 76 FE C1 BE 7B ED AD 7C
 59 BF 8B 9B 8E E4 8E 2B 51 04 93 BE 39 B4 EE B7
 AA 71 37 41 C8 99 F0 22 74 BD 5F 04 43 B2 AD 24
 98 9D A6 E8 82 E4 75 8A 9B D5 AB E8 03 A3 B6 68
 80 66 D1 96 60 AF FC 2C EF AF 9A E0 13 71 CD 31
 70 6C 95 3C 1F 6F 7B 43 5C 25 79 B6 9C 46 F4 17
 07 93 CB E3 6F 8B 37 0A 29 5B FE 69 EE 7A A5 B3
 6E 41 AE 3F E2 E0 64 76 82 B8 47 05 54 87 FB 11
 56 9A DA 76 DD 27 F0 8E D6 E9 24 A5 22 09 D5 8F
 AD CE F5 9B 22 6A 1C C4 BB E7 1C 87 42 DD 43 2D
 F1 C6 0C CA 78 1E 45 FB 21 06 58 78 0E 13 8A 4A
 D3 4B 4A 78 D5 B5 E4 5F 3A F2 C3 1A F8 C2 52 59
 31 A3 41 06 60 F8 D9 80 B3 8A AF 6C A4 C7 9D 45
 BB 86 AA 6F DE 92 D8 1A AD 7E EA 2F DE EC 1A 2A
 9A 46 F0 3C 92 FA 19 8F BC E6 12 D0 DB D6 22 6E
 3E 71 9B FE E3 4F DE 06 42 10 22 D5 BB 6E A0 C1
 A0 F6 E5 75 D7 62 47 58 22 E3 E5 67 14 5A 9F 69
 13 BE E4 C5 6F 84 71 81 4A C3 D4 AE 34 16 18 D5
 AC F4 A9 6E 38 88 71 C8 8B 92 2C 24 D5 99 72 F6
 8B 0A 07 CD 83 89 0F 65 AE 29 06 4B 00 1E DF 80
 30 03 28 34 F3 AA E9 42 23 6E 05 3E 0F 4F 25 C0
 0A 5A BE 71 38 BC 77 4C BB F6 76 75 F2 35 97 A3
 4D 2A 4F 54 2D F8 21 B2 5E 22 66 50 A0 F4 01 21
 02 8A 35 A5 84 BC 82 15 9A BF 27 0B 4B FF C5 AA
 98 52 95 75 F8 DC C1 0E 86 EE 9E 26 CC 08 3C 96
 00 9A 6D A3 5A 8E E9 2F 8A 5A F9 B0 34 8C E1 32
 F5 5F BA 17 8B 76 4F 5D 6C C3 2E 34 63 C0 E8 7F
 C8 4B EE E9 3D 2F A4 21 F2 3B 07 31 4D 04 B1 87
 16 1A F9 39 93 05 95 48 E5 82 59 68 E7 9C A4 7A
 B9 CF E0 F4 A1 A7 E8 18 98 B6 79 9D 51 6F 0A 53
 CA 8C A9 8D 70 82 4B 76 43 E2 5C 84 02 29 C6 B7
 8D AB 69 4E 3C B9 A9 5E F8 8E 7F EC 39 D5 07 68
 04 55 C6 9E E9 1F 74 60 6D 62 CC 3E D6 71 4C BC
 89 81 2A D1 83 57 53 81 8C 05 0B 2C A5 94 F6 EE
 D9 05 3A 57 B4 0F EE DA 9A 64 8C 49 23 C4 08 36
 0D 45 0E 7C D8 BB B6 F9 0C A6 EC 73 29 DC E9 51
 18 5B 67 9B 2E DF D2 CA F4 0F 55 4F 3A C5 F0 42
 EA C4 1D 55 3F BF AC E3 F0 C8 D4 9E F1 A7 C0 2B
 BF 0C AA 02 82 BF 8C 3D 65 E9 71 93 A9 F4 E4 5A
 92 05 84 FD 3E 1C 4A 9F 2B F4 17 41 34 C9 BD 42
 F7 95 01 43 26 1D 92 21 27 AC 87 59 D4 11 C3 FC
 82 DB 99 91 98 6D DE 8C 8E 3E 7D E1 49 C5 0C 8B
 66 9F 51 54 C2 3C 26 7D 6D A8 64 02 0E 33 AE 54
 F3 26 65 22 EC 67 2D 1F AE 5F EB 24 B0 75 3D 07
 58 DA 6E 0F 96 F8 3F E9 B9 1E 9F DE 28 58 C7 EB
 EF 61 39 8E F5 79 A7 6B 5A E0 64 3F 87 E4 C5 F9
 CF A5 38 E8 A1 1C 43 3C F2 8F 5A A2 25 EE 55 0D
 EC 5B 04 57 DD AA E5 C2 BF 07 95 41 0E 6B 97 0A
 86 F2 A5 08 A5 DF A8 7B D5 88 C4 F7 D0 41 92 A7
 B6 83 4D 6C B6 01 BD 0C 53 30 E4 9A F7 71 A2 57
 5E 3D 50 EF 3B 65 33 37 FD 9C 6E 58 5C 99 F6 52
 ED D5 74 32 B6 65 75 13 28 D8 34 C5 C0 80 02 13
 EA A9 F3 6D A6 6E 0C 16 B2 AC 50 8F 35 F5 2C 2F
 81 99 92 F2 D1 97 BF 41 4B 27 A7 1C DF 2E CD 33
 44 B3 54 36 E4 8D 79 39 BD 72 2D 56 EE 62 C7 6D
 E5 18 EA F0 8C 85 8A 75 41 2B 2C F4 92 3E E9 5B
 DA E2 D4 E4 5A 55 E5 62 BB 86 AE 6E CC 1D 9E CA
 ED 20 A0 07 B7 7D 5D 63 3F 85 6A E5 83 DC 04 68
 B7 37 D8 47 09 DE BA 19 6E E2 81 D6 D8 32 52 C7
 30 4F FC 24 E3 46 12 2E F8 11 C4 ED 2F D5 B9 69
 36 21 1C 01 3C C3 DE 13 E5 78 94 F5 7E 8D FD E3
 47 05 05 32 0B CB 5D 7F 77 67 0D 38 2E AA 35 1C
 92 9F B3 B5 42 E7 A4 F4 8F 35 32 6D EF EE AE 87
 49 05 DB 95 C6 A0 C4 F0 0E 17 2F B7 2C A2 F7 E7
 C1 27 E4 F0 B2 E2 5B C6 58 C1 A0 FB 2A 81 8F E7
 49 B0 61 DD DE D7 56 BE C2 D3 F7 F3 67 42 9A 22
 E9 1B 1D 5C 2A 41 FB 54 12 FF E0 77 DB 5D FE 09
 09 F1 45 74 F1 05 D9 9E 76 40 3F 8F 9B E6 50 FE
 8A 70 A8 51 7D 46 94 D8 70 94 34 51 6A 93 DD 0B
 37 05 DB FF 84 DC 36 32 0D 3B 6F 57 AE 4B 6D E0
 55 B7 5D E9 5F B2 F5 B4 8F D3 E5 5F 8C 9A C0 6B
 B8 20 F9 91 42 F0 7A C7 32 90 0A 2F 3E 41 25 E9
 88 AE 63 DE 2B 0E 1B 96 9A 7B 92 D2 0C 80 55 B1
 D8 D8 DD 35 E9 BA A6 86 34 49 0B 45 CF 0D 53 F1
 D1 BF 8F 59 AF C5 75 8A FD 10 43 62 D3 35 D5 55
 8B 24 EF 7E 8E 80 63 34 D8 4A C9 F4 47 8F 34 71
 D3 3E BD E8 97 2E 69 81 82 01 B2 13 30 60 2F 77
 EB 35 AE 73 55 3B BB D3 91 02 91 B9 52 F5 62 13
 4F 78 3B C0 DA 96 45 FB 62 66 B3 E7 E3 8F F3 23
 F5 94 41 73 4E 43 4F D1 5D 5A D6 1D 2F D6 C9 40
 33 98 40 57 4B AD 86 7C E2 7D B0 60 C3 0C 64 E3
 F2 69 8C 53 3A D7 99 FD B8 AE E4 C8 AA A3 78 30
 48 91 DF CA 99 5E 21 75 F4 E7 90 53 63 7D 5E 3A
 6F EA 8D CC BF 9B 06 D2 48 A2 38 8E E9 D0 60 4F
 B7 68 53 C8 0E 52 FC 26 3D 1E F0 B1 97 F6 0D 6D
 8E DD 07 27 CE CA 1A 7A 59 2A E6 C6 15 F3 3D CD
 EA C4 B8 B1 12 D3 BC 42 B7 DE C5 A7 B3 8E 1D E0
 04 5B 3C FD 40 09 0A D8 AD 65 EA B3 6D 96 02 26
 BF 22 0F EF 53 32 BA 1C 2A 0F 1E 29 7D 2F E1 80
 73 9D FB C7 2F 28 4E 11 45 97 4A C9 8F 2D 22 BE
 8C 7C F8 26 25 44 14 88 66 61 3E 30 B0 39 13 A9
 7E 3C 01 72 F0 6A C3 9F AC 9A 33 DD 75 6C 45 A7
 D3 AF 84 E1 01 17 BC 8A BC FD 65 F6 2B 9F 18 CC
 C0 33 20 8C 46 D0 08 92 90 E0 56 ED 73 88 ED 11
 59 70 C7 75 7A 3D 16 DA A5 89 1E 1E 6B 0E 08 A9
 1E 82 F6 32 BF AB 0B D7 F7 39 E9 7A 1A 73 06 6D
 E6 2E 3B 37 B4 0E 72 7B 8F 50 CC F7 05 F1 74 3D
 D8 28 2A 38 47 FA 92 D8 08 E8 44 5E 3C 3E 55 D8
 81 B7 D3 BD 5D 73 A3 0C DE 45 54 BC CC 5E ED B9
 B1 34 A5 EC CD 1D F4 EC 43 F3 BB DB 08 3A 35 B2
 D0 18 04 58 F8 D7 B9 E5 8B C0 3D ED 80 AE D8 CA
 7A 90 D6 48 8D F8 8C 48 D4 DE 48 A6 6C 43 C9 58
 1A 4E B9 A9 F1 C7 20 24 AD F1 DF 1E 4E DE E4 F9
 88 D2 E6 6D BC E8 6D 30 BD E8 22 05 8F 21 9E EB
 30 A8 A1 29 2D C8 2E 7E 83 CE 06 F7 9E BE 8D 70
 DE 64 03 F4 73 BE C1 80 32 72 98 1C F1 C2 12 61
 F0 62 D9 41 AF 35 DF 1F F4 E3 07 55 D9 96 07 0F
 78 29 34 23 56 86 59 1E 23 72 99 C9 DE 40 EB 28
 53 6E B2 CC 7D 76 38 CD 20 40 9A 02 B6 2E 30 F0
 C0 32 90 E0 1B 5B 6C F1 7E FF 8F AD F3 99 E7 55
 E0 66 A9 D7 38 8D D6 6B EA E6 A4 40 48 A7 0C 3F
 45 64 CE EF 7D 75 BF 3F 30 B3 3F 9F 7F 16 A5 36
 31 88 7C BA 0C 15 3E 1F A4 F6 19 78 81 91 3F 79
 FD F2 2B 44 93 6B 4A 1B 13 82 90 5F 32 F5 AC 4C
 22 13 D1 FA 1C FF A5 E7 AB 96 3B A3 8E 77 58 05
 4D CC 49 DB 30 9E 70 C5 E7 6D 86 E7 32 B2 DF 00
 76 40 06 ED 93 63 55 67 0B 8C A2 D7 C7 F3 96 0C
 DC 67 34 00 F8 54 58 C0 C8 B0 11 30 0D 16 28 53
 A8 F7 54 DC 4F 90 73 53 73 99 AA 05 0C 22 84 24
 D0 B1 20 14 80 46 A2 12 0A 91 AD 41 42 E8 45 9F
 D3 F2 1D E5 35 C3 2A 77 CC 8D 39 45 07 9E 64 0A
 BA 40 C5 F4 F8 FF 77 35 2E FA 0A 77 4B 3A 88 B0
 4D 60 43 AF 8E 75 61 F3 28 AD 5E 10 F7 3E 8A B8
 E9 37 71 A5 1F 65 40 B5 A0 AC 8A 2F 03 70 31 96
 09 A5 F9 E1 C5 63 90 5C 8E DF 02 EE 61 3F 8A F2
 F4 B4 E7 9D 3E 0C 86 E5 B7 86 BC 13 B3 F1 D1 9D
 0A 3D 8D 3D BD A6 02 B6 75 61 B1 05 16 B8 9C E1
 DD 9A B7 BC 80 D3 AA 32 78 A8 AC 62 B4 59 A4 71
 18 CF 97 25 9F 57 37 56 E6 47 6C C7 34 A4 9F 1B
 59 63 32 EC 7F 93 48 2D 8C 89 BC E1 39 17 03 35
 78 53 92 5F 23 DB DB 0A 8D 3D 3F EF B9 F4 12 9E
 B7 7D 1C 3A 74 37 AC 78 A0 3E CA FE 6C B7 E9 65
 CE F4 EB 3D 49 AC 38 18 A7 E0 12 21 3C 7E 3C E6
 9B 10 EE 08 32 C7 B3 2D ED 33 A7 98 8D 86 12 5E
 BA 16 18 E7 74 0F 56 1A 96 70 68 0F E1 95 47 10
 6C 28 5F 0E A3 7B 7B B6 D0 90 ED 66 E0 3F 4D 6B
 C7 2D 2C C2 B0 CF 63 AD D5 A5 8C 88 DC 22 2F 1E
 6E 9B E8 1F C9 CB B1 52 56 26 FD 92 8F AA FB EF
 54 9A B7 6B 36 F4 4D 6F CA D0 97 31 54 D0 48 79
 05 F3 9D 66 5D 19 B2 61 72 AA AF F7 D4 3C 8F 24
 69 C1 8A FC D6 5E 6B 85 3B 65 CC 5E 13 87 44 5A
 7B D5 2A A0 71 8D D4 5A 1A 89 0C E6 4F EF AB E4
 C7 48 06 65 AE BC D7 65 7B CC 03 AD 28 56 85 F0
 D4 B1 3C EA D7 6B DF 8A 0D 1B 23 5F 32 34 ED E6
 B4 A5 7D 86 8E A9 D7 B4 54 53 B7 D9 5B C1 34 D8
 E4 D5 CA C0 20 72 56 A1 0F E1 19 DE F2 A8 77 6E
 51 F6 32 A9 15 FC BE 2D EB 5B EF 39 61 FB 67 1C
 69 95 FA 98 71 19 92 22 46 FE 47 BA 0D 36 1D 77
 29 9F 62 21 1E AD F4 59 13 60 C4 CE 3B 59 61 DF
 91 06 3D C2 24 0B 6D 74 DA EA 90 8D 8F 0C AE 15
 85 35 3F AD F9 E9 22 77 30 20 0B 06 A1 0C D7 3F
 55 16 8A D0 6A FB 43 9C 65 A0 A6 87 90 A3 A3 CF
 63 7B 52 AC D7 8B 06 31 29 18 D0 5B CC 4F 85 81
 E9 E1 26 24 5C 1A AB 1D F1 22 1E AD CB B7 57 E3
 6F 75 98 59 4A 46 BF 0C C8 FC 1D 83 E3 1D 0B EC
 FD 2A 91 C7 FF 27 A8 95 0F 67 7E 8E 10 2B 66 1D
 4D D9 E7 53 D6 2B 3C 97 40 21 40 D9 3A 3F 39 F3
 17 2C 20 69 94 21 F6 52 D0 7D 72 5B 80 41 49 F9
 92 9F F7 A0 BA BA EB 05 47 EF 10 E9 A4 29 FC E4
 42 6F 34 09 10 4F 09 BC DF 6C 64 94 90 CD 18 E8
 32 EF C5 11 A4 C3 73 EE E8 E4 FD 69 14 B8 95 5C
 92 5C 26 DE 24 EE 43 78 C3 9C 85 75 BC 37 5B 34
 39 FE 10 10 C1 1E E3 1B BD E9 3E 5F A4 9E 7C 4D
 08 EA B0 1E 54 74 80 03 B5 EF B1 71 F6 0C D5 B8
 93 4E 8F DF AD A8 BB 8E F7 30 10 01 E9 30 78 B1
 D0 A3 E1 FD 4D 1A 5D 5A 67 65 71 80 98 A0 C7 67
 08 A7 DC 55 9C 6D BC 5C BE B5 E8 95 21 39 9D C8
 18 2B C8 BD FF 03 14 D8 D0 1E 88 68 E7 A5 C3 4F
 D8 42 17 8B E5 DF E1 FF 8C 0B BB DE 2D 40 D0 D4
 C1 D3 95 4A C4 B1 A9 D4 36 52 F6 8B F7 51 EE 53
 98 01 13 7D 47 84 6E FE A2 B4 2E 5B E1 12 AF 41
 4D D3 52 47 90 59 DF E7 BF 5D 58 9D D3 45 12 F3
 42 4E C8 DB AF DC A9 45 6C DB 01 0A 26 D1 73 78
 41 29 BD 08 EE 2C F8 83 14 D6 91 7F A8 00 0B DC
 9B A3 0C F1 91 30 1B 15 F5 C1 94 10 30 13 33 F4
 9C D3 00 9D 3A BB A7 9C D5 D0 E1 E5 08 77 AB 37
 E7 2C 51 1B 6C 9A CE 3A C0 62 FA A9 87 A2 F6 65
 21 BF 52 35 75 19 6C CD 33 5E 20 AF 96 60 71 9C
 EE 6E 46 E2 7F 53 B3 A4 86 18 B0 65 E5 FD 33 3B
 DA 55 10 69 03 99 DC 35 F9 54 D1 3B 79 9E F2 7F
 B0 E0 0E F2 C4 3A 2F 24 BE FD 51 27 2B 46 9C B5
 93 43 59 1A 2A A5 E7 E1 02 3E 77 B6 2D 42 01 45
 CC 0F 38 0F A6 46 36 E5 9C 25 6D 4C 39 95 AC 71
 21 CD 3D B3 48 7F 79 0B A0 02 50 FF D5 72 DC 13
 5E 41 0F B6 00 70 70 C0 5E 02 AC 4B 38 B8 D8 E5
 2B A0 39 8B B5 C4 F3 A5 69 51 C5 BB 57 B7 EB EC
 A4 1A 98 03 11 6A DC DB 4C 81 32 9D 8B 50 57 A9
 11 35 B5 84 89 E6 CE 95 59 D4 DB 57 46 1C DA D9
 95 FB 5A 01 83 9C 6C 88 21 2F D4 DE BF 92 2C 59
 36 AF E3 A4 C1 21 A9 DB 60 17 08 46 9D 6E 4E 2A
 A1 70 CE ED 2B 09 21 37 FD AB EB A4 9D B1 AB 25
 9E 28 F2 44 D6 29 DF CD DC 41 7D C8 93 F6 37 60
 18 F4 E9 11 03 42 AB A7 E5 1E 1E 97 A0 08 DA AA
 09 3D 9E B1 21 E5 9D AC 87 14 C0 36 ED 7F DD D9
 42 4D C5 C2 C7 5D 16 F0 F4 22 E9 63 79 43 65 32
 E1 14 8C E9 D1 BD 0E 0F AF 3D 5F B9 18 0F AE F4
 C5 3B BB 74 EA 45 21 76 ED 82 02 66 40 38 A7 D0
 57 83 4C C0 8B FE 77 FF F2 CB D1 44 8F EB F4 8E
 D0 73 8F 09 8C BA 58 06 FF 99 6B B7 07 DF 50 7F
 F4 3A C5 50 E2 EA 81 5B 31 56 D6 A4 01 90 D1 17
 8A AD F6 7D D1 CC 6E D4 DE 95 AB 0D 0A 62 3F DE
 89 64 49 C0 1D 63 DF 66 4D 5E 59 CD 61 1E 20 FE
 AA 8A F5 3A 2F 70 A6 09 37 A4 5D F5 A8 74 B7 81
 05 3D D1 A0 27 89 65 67 6F 41 FF 73 31 C2 46 27
 43 AC 10 96 93 D1 4A 96 88 1D 4A 12 C4 C6 E1 F9
 3D 9B 9C 8B 58 7C 1F 6F 33 97 85 FF B6 05 41 05
 8B A4 F1 EF CF 6B CA 3E 12 7C A2 3B F3 B9 AF 4C
 90 AB 7F F1 C7 9F A0 D7 03 77 BE F4 2E 69 2A 68
 A0 51 29 78 63 2C D5 74 7B C0 93 C3 D3 0B 35 5D
 5E A0 65 47 8B 7D 1A 6B ED B6 CD E1 11 85 D0 DC
 F2 2B E7 12 EE A3 AD 46 54 80 D8 F9 09 C4 85 FA
 4E 63 7F 67 61 AD FB 67 99 37 4A B6 C3 F2 12 20
 CC 73 EE 73 1E EB 27 4C 54 C6 1B 96 44 7A 78 25
 D8 67 8B 6F D4 3A 2A 66 91 97 62 29 28 3F 94 29
 44 8A 76 18 34 49 87 DF 6C 2F 96 CB D1 59 8E CB
 2C 66 66 74 28 19 CB 21 1B 0B BD A9 7E C3 DC 65
 7F 8A FB DD C5 AD FA 57 B6 54 73 18 C1 27 2E 6B
 7A F3 9A 90 5D F9 25 A9 11 77 36 B1 CF 6A FE AE
 BF 91 86 56 28 F0 32 C7 C5 B7 89 80 B3 A9 79 7C
 80 23 E8 96 DC E6 B2 07 01 89 9C E3 FA 04 F2 A0
 CA FC C9 DD 63 DB FD 27 42 96 85 82 32 14 A0 69
 32 3B C5 98 4F CA 3C 6B D8 50 7A 84 F2 8B 84 F3
 EF FC 8D DA 8D 4E A4 AB B7 0C 8D 25 68 1F 6B A3
 8F 16 D3 75 49 16 90 1D BC 23 66 52 09 2D 85 0C
 99 F4 C9 DD 30 4C 3E A4 E7 60 1B BB 81 ED 88 4F
 83 57 D6 F2 9F ED AB B1 AE F3 D9 F5 CD 38 3C C1
 25 33 C7 5C 5A 2A FB E2 5C 48 F0 6C 8B AE 41 27
 50 DB C9 8B 2C 14 FF D1 0D 39 14 48 B0 9A 8B 5A
 2A F5 36 44 62 AD 1F 1B 1A 1E 32 81 28 75 D0 97
 4E E0 79 77 3F 2E 71 18 4C B0 9F 2E 38 F6 92 D0
 67 CC D9 26 65 32 FF 63 4C D5 BC BA 27 5E 4D 00
 EB C6 5E A5 03 46 4F 2B 5B 36 52 5C F8 6D 4E FE
 4C 5E 4B 23 F5 F7 11 5B 56 38 F8 21 01 01 7A E2
 FC 7A FD C0 07 5D 22 BB C0 2D 6B 29 C0 C2 1C CF
 27 4B 16 B0 0D 87 97 2F E4 5A 65 61 9D ED C1 20
 48 AF 78 63 02 0D C7 B3 DC 1B B4 FC 85 E9 40 1D
 E6 F3 49 E5 07 77 AC 3D 46 09 17 46 8E EA 4F 7D
 0D E9 92 B1 67 CC DB E7 00 33 E5 1F 70 34 F9 86
 A6 78 92 8E 9E 4F 92 EF 10 DA 05 15 68 51 1A 56
 BB 28 D6 93 06 8C 9B 05 D9 44 9F 1E 3E CC 70 9D
 8F B4 07 37 AB 43 CB E1 C3 99 41 64 F1 E5 39 73
 68 08 06 2C 34 90 5E 4A E9 06 60 66 94 46 27 00
 6F BF A1 C3 30 93 9F 81 CA 89 24 4F 54 ED 14 12
 9C 1F 48 42 27 77 52 1E E0 E8 B1 7A 27 83 2C 38
 A8 FB 99 4C 7F A9 57 34 AE BB 3A 28 E6 B3 75 B5
 B9 73 42 27 41 3F 34 0E 8C 57 6B A5 BE D2 C6 C2
 5D 34 71 91 93 CC 33 41 16 7F 19 64 86 3F AC D3
 B0 DD 63 D9 B7 31 50 0B 4D 59 7C 7A 7C 5A 1B C5
 99 09 26 4C 76 8F DC B6 69 48 28 E4 A5 E8 42 28
 81 F9 F6 83 0F FA 7B 9C 9C 84 4B FE C9 19 D4 A4
 B1 BC 79 47 13 E8 61 D2 12 61 AE E7 17 16 3C E3
 81 BC 22 64 17 D8 B1 35 40 93 F2 43 E5 3A 45 A7
 D5 94 85 44 39 10 B4 6A 85 3F 72 8B D8 EE C3 BC
 E6 6C AD 62 0C 38 C3 CC D3 A5 1D 0E 20 CC EF 4C
 B5 D5 B1 17 06 21 30 7E CE CA F0 E0 08 EB CD 2D
 79 88 CE 44 C8 E2 4D 60 96 97 6D 52 C2 EC B5 02
 44 D0 A7 47 99 29 D6 0C E5 EF 2F EA AD 41 7A C2
 EE 5B 66 82 73 69 14 52 AF 5E FD 06 06 20 22 B7
 E3 95 AF 72 67 EC 25 28 46 EE 30 AD A5 85 3D A7
 1E 09 27 31 89 DB 94 20 84 69 2B E5 AD AA 1B 12
 40 12 01 2D 4D EB 2D 25 B0 DA 92 FD F7 84 72 7B
 AF 20 06 2C EF B7 3D 2E 89 10 F6 48 68 A2 39 8E
 7A A7 0D 70 66 0F 44 34 DF 80 43 28 1E B1 AA B5
 6C 26 B9 7E CE EC FD EF DA 76 C8 6C 24 A2 94 C7
 BA 25 F5 1D D0 DF 27 C1 3C B3 77 F0 7E DD FE B1
 DE 04 F8 2D 18 C5 F6 73 9E FD FD E6 63 C9 C7 14
 A4 FB 1F 6D 7C 33 52 72 5A E2 89 50 F5 3E CE 1F
 5A F3 18 0A 4B D1 BD DC C6 A3 7E 6B 58 B5 0B BC
 7A 29 98 71 42 EA 3D 16 AC CD 95 EF 5E 55 3C 9B
 FE 72 23 28 AA 73 F1 FA 30 A4 A8 53 84 09 2D 42
 C0 B2 F2 4D ED 07 A0 F0 DD 25 35 F0 17 F8 1A 2C
 A1 E2 5D 5C 61 C6 4C 0D D4 15 69 BC 1E 52 B6 B6
 9E C1 FC A0 0A 9F AA 1F 30 E7 59 10 C4 04 58 D4
 05 1C BD C3 45 AE 1E 56 65 8E 9B 8E EB EE EB C1
 1B 81 8C 7A 5F 6E 56 3B 86 6F 2E 5E A5 98 A2 A8
 AB 5D EB B1 C4 9C 4C C4 F6 A5 70 F7 7E 28 71 CB
 E5 3E C0 91 E2 68 AB A1 A8 F3 99 8E BB 53 C9 65
 14 15 82 97 8C 91 3B AC 53 F7 57 DB AA E7 3C 6A
 74 10 3F E4 14 9E 5B AE DB CF 4A 9D C1 11 8E 3A
 E3 80 52 F3 A7 C8 18 6A 9A 00 7A AF 8E D1 68 70
 2F BA 88 12 05 5E 3C 14 DF F6 71 69 2C 7F 80 C6
 A2 EA 9A DF 75 B5 F1 04 5B 14 94 15 A9 A9 89 C4
 C8 81 58 F4 1B 52 87 40 F1 4A 2F 8C A9 4B 5B 1F
 B9 D9 F9 8F 5C 19 F9 75 90 0E 59 89 24 B0 E0 BF
 82 39 31 C1 50 4D 90 67 0E 67 D2 3C 4D 58 97 46
 67 E7 33 DB A7 34 91 7F B6 28 1F EA 70 0E 6C 52
 1D 17 A0 36 7C DE 6F 4D 9C ED 88 9A A3 F9 B2 2A
 F4 57 32 BE 99 16 57 75 07 DF 29 9A 72 DB EF 28
 A8 6A EE 52 41 22 B9 31 2F B2 A0 F2 FA D0 B5 2B
 FA 86 4F DB D4 DA 86 3A 61 5C 0D B6 0A 13 6D 8C
 E1 98 50 7E CB EA 5E 19 54 4F 53 C7 75 FD 7E FD
 43 1E E9 BC 02 6E 85 6E 0C 27 27 54 44 65 F9 1C
 55 7C C8 F4 79 29 28 57 FD C2 6E 4D 04 C1 78 68
 F2 58 0B F6 4D 29 ED 92 BC 11 18 0F 31 80 1B 90
 54 07 9D 9D D5 1A C7 2A 6C 5B 31 5D 83 BA 7D E4
 0B EE 4A 22 8E 35 F1 2E 71 CF 77 54 DC 4B F2 89
 54 65 CE 7C 95 54 A8 D2 A5 8C 3D 98 C2 42 75 A9
 7D A5 02 CF 4E EF BE 50 EA 32 5D 27 B6 17 F8 90
 7F 02 91 C6 3C 5F 7B 07 72 51 38 29 28 9E 84 C0
 F2 19 E2 4A 34 1C CB A1 D8 1B 36 F7 04 4F 7E 60
 34 C2 CF DF ED 19 4C 9D 24 5B 95 DB A0 37 C9 67
 AE 7A C8 47 43 29 48 1E 83 C7 63 62 DF A9 82 EE
 AC 79 6A 00 00 5D 66 A8 77 58 4E BA 59 73 FA FF
 C9 B6 C3 4A 67 62 36 DF 6E 2E 0C 72 BE FB A1 29
 15 26 9F B0 32 44 F9 DD E3 E6 0B BD E5 4B 03 14
 C2 A5 D8 41 49 8A AB 4F DD D4 D5 C4 90 6D 4E F7
 F6 6F 89 C6 5C 1D 63 DA 7F EA 8A 86 86 77 91 E3
 73 2D 2E EA 8F 21 B4 ED 9B CA 62 BD 87 30 9E 13
 4C 55 2B F3 C1 88 06 50 86 2C 23 BE 2F E2 7A 3C
 BB 03 CF 47 44 AB D4 FD 5B 4D 28 B5 1A EC 8D 36
 78 D2 AB D4 6F 77 9A 17 A7 44 97 E3 34 D2 90 1E
 20 99 A1 1E 07 16 08 AB 57 5A B2 91 38 98 14 A4
 C1 40 E2 3F C9 00 A5 D0 D2 D0 A8 AE E4 83 AA D4
 73 5E B2 CD CB 88 5A C9 94 7D A8 2A 64 CF 3A 78
 E3 9E FE 80 36 16 98 37 AA 82 03 CD A7 A1 20 E4
 2C 3E 43 2E 27 20 06 78 60 7E B7 AB F2 4A 21 FE
 3C 10 40 53 E9 FA 54 F8 F3 EA 07 19 A1 9E 8B 3E
 BA 3A 07 7C B8 9E EB A4 C4 57 6B 76 22 25 07 E8
 02 25 3C 6C FA C6 AB 11 E8 E0 3D 39 4C 53 A2 5E
 74 4A DF 00 04 E1 E2 1F 1E 1F 8B C4 91 5C 91 F3
 14 FC B0 C2 B0 66 A9 6A 3B 9A 6D 73 CE CF 8F 97
 6C 2C D6 80 B3 CF CF 74 52 A1 DF 32 1E 65 50 F5
 BA 04 CC 15 F6 7F C2 70 17 CB 64 34 07 72 31 B8
 51 5C 86 5D 95 D5 17 2C 5F 44 9E DC 8B 14 D3 32
 02 C5 F3 10 C0 AE 95 BC 1C 98 EA F7 4F A3 AB 4D
 1C 63 B1 CC 6E 84 0B 67 2F 52 D7 A3 62 30 29 40
 31 23 EE 14 EF E4 07 2B 00 29 44 9E C3 16 65 AC
 60 3F 44 38 D8 DF 76 89 98 A9 44 A2 C5 CA AF 38
 99 52 9B 8D 61 8D 08 44 20 13 AE BB C4 EB FC 45
 7B 24 5B C5 1E 91 8D 40 E5 A0 5B 51 7E 96 D1 AB
 F2 81 6A 6F EC 32 B0 BA 21 8C 55 55 3D BA FB 50
 37 3C 0F 78 A0 B2 B1 EC A1 B7 6E D0 43 B1 5B 5F
 1F 89 EC 8A 37 F5 FA A3 38 75 C3 92 8F 61 63 1F
 26 58 DF 9C E1 E2 77 D1 10 09 D5 CC A4 72 6D 7E
 31 84 D4 EB A8 72 9F C7 E0 5B B8 3E B5 02 35 C6
 D3 03 B2 F7 DD 6E 29 CC F5 4F C8 FE EC BC AB 13
 AD 05 4C D3 6A AC CB 41 52 0F DD E7 58 1B 36 AD
 94 49 CA 43 BE F4 38 02 14 60 A0 E1 88 7D 53 C5
 E2 0C 9A EB 1D 2F DE 3D E4 CA BF 11 B2 7C 67 6B
 44 7A A9 82 33 02 C2 78 2C 6E BE 78 0B A8 CD 6F
 13 38 F5 5D 5D 86 C7 09 BD 45 E0 7D 63 C7 A1 99
 6E E8 56 FB AC 09 2C AA 4D 39 D2 FE FA 5E 43 DC
 D7 B1 ED 1B 19 0E B8 5E A8 CE 2C BD E6 7A 18 50
 FD 95 EE 4B 32 FE 85 CF 67 4D F3 62 15 19 9C 6F
 E3 AC 02 C5 7B 9F 7A FD 64 E1 A3 34 C2 27 96 2B
 A5 01 FA 46 2A 73 47 73 E8 F9 CD FE EE 9C DF C4
 A5 33 43 F3 29 57 3E 49 74 D3 6F 83 89 03 26 9C
 84 CC 2F E6 0B D3 FB 75 92 57 E0 A6 F5 12 A6 4A
 72 2A E9 BB 80 BB 77 FB 2B 7C B7 18 12 0D 46 B5
 33 31 93 AF 12 8D 4B C5 12 3F 60 00 83 1F C0 1C
 D8 51 FB 03 75 BE C8 4F 3D 37 F7 42 B8 46 34 E7
 C5 A4 EC 7A 6A FF DB 6F C4 66 D6 95 32 7C DD B5
 62 79 CD 28 5A 54 26 1D 38 E0 4F 48 D6 72 B5 7A
 B0 32 35 44 87 BC FE 1D F9 FC FF 64 32 6C DC 6B
 46 4A 0B 42 73 AA 34 EF 84 2A A9 87 5D B8 4F F2
 43 AE AC CF B4 13 35 DD AE 72 11 92 AB E6 34 A3
 C3 A6 C8 83 46 EE 1C 39 77 5D 0A 47 6B C0 88 6D
 72 AC F4 4A 65 37 F8 79 63 39 0B 4A FF A8 5E 04
 B7 26 41 A2 C1 91 15 8F AE FC 86 86 55 C7 47 0E
 24 5A 69 2F D3 69 7C A8 48 2F 37 73 7C AA CC 48
 7B 26 C0 BD 6D A5 71 00 EA 6A 62 A2 F1 A5 7B 28
 9C 73 0A 0B F2 03 71 7A 5E 29 5D B5 E8 8F B8 5D
 14 18 72 70 73 67 4C 57 D6 C6 78 0B 68 B6 03 BB
 EC BC D7 D7 E9 39 BB B7 E3 88 DD 89 D0 06 1D C1
 A7 AB BE E9 89 7D 84 92 FE 28 A0 6F 0E E6 73 3E
 90 A3 6F E7 E0 84 5F 86 52 AD 1E 8D FB 58 0D 40
 54 FC D5 DC 56 A7 2D 37 71 61 0D 80 35 DA 5C 91
 91 F9 72 40 EB A0 08 14 26 0F A1 73 B2 2A 58 1A
 53 21 45 F1 DB 64 94 63 3D 50 C6 FB 23 73 6F BA
 C6 14 42 13 EB 00 14 26 F5 7D 2F 6C 71 12 56 F5
 FA BD 9E B3 3B 0B 0C E8 4B C3 7E 31 3C 8B C0 EA
 90 7A 6E 2D 84 D5 31 EC 26 1E 22 4D D7 38 42 A4
 04 7A AB 1B 78 1E B4 E9 36 D7 5C 57 B1 23 FA 1A
 C8 17 0F 7B 73 02 DF 8E FC 35 10 3F 02 EF 7A 81
 DE 83 49 6F 35 33 ED 25 81 C6 C3 50 F5 51 99 E1
 5D CE 86 7F 07 44 6E 56 90 75 37 CE 29 C0 4D A3
 45 F9 70 E9 5B 00 8F BE 38 EF BD C3 B9 E0 76 76
 E6 00 25 89 A5 FA 96 10 7A EC E7 B0 A7 CA A5 17
 3F 2E EE 4C 61 D0 72 96 38 D5 3D 30 AE 3C D8 A2
 3B B8 F8 F1 91 B3 15 A9 A8 8D DC D0 96 03 95 36
 A1 DC F9 67 D5 D7 C9 56 97 76 6E D6 E4 93 4C 98
 50 8B 42 F8 9D 2E F7 14 05 D0 08 E2 D7 43 4F AA
 FA 9B 11 93 DF ED 71 88 CF ED BE C7 4D AC B4 F1
 B9 D1 E7 B4 CE 4A B5 A2 84 E0 DE 7A 74 42 A6 B0
 82 B8 05 7D 69 66 E9 36 56 AE EA 5C 3C E9 75 17
 71 DE 09 EC C4 F3 40 63 13 D4 AC A5 9E EF 66 B8
 D4 4A 33 91 9E 18 19 76 50 7F 7B D0 CD CA 63 2E
 13 47 AA 0D 68 9F 41 74 DE AD B4 F3 F9 60 38 3A
 AF 50 32 57 9E 3C 37 E2 D7 EF 8D BB A2 F4 1B 29
 B4 30 44 87 15 AB FE BC 07 7B 84 3F 31 55 BC 00
 15 33 38 C9 16 ED 41 68 0E 13 0A 61 11 58 5A 7D
 A0 9A 29 72 5D 2E 4D 5E 1C D7 FC FB 86 02 C7 26
 FD 29 80 AF 6B BF 14 44 4A A4 03 60 93 66 C8 CC
 DC 3B 83 5D 43 FF A6 F4 D2 BC 35 A6 9D 88 92 8B
 95 9D 36 2F 44 24 D7 7B 46 4C 40 32 10 5F 2B 34
 E4 4B 6E 9F 47 2E 77 72 95 2B B5 F1 1B 89 B5 BD
 64 F1 67 AE 35 50 F5 77 4A 40 3B BF E7 20 FE 66
 8C 38 3D D3 43 F4 89 84 30 52 F7 08 A4 4E 1A 67
 8B 10 FA 23 EF C0 10 97 51 59 C1 AF D7 2E 79 3C
 A7 24 9E 63 4F C7 73 98 42 5F 2F 3A 9D 43 34 DF
 15 B2 85 2A A2 8A 7F E7 8B 00 A7 BF 7C 66 5B 2D
 9B D5 09 A1 A2 49 9E 7F 07 2E AD 74 F7 9E 6D 11
 3E F6 C7 E9 08 77 BE 16 8B 58 BE BF C6 5E C1 3F
 66 4D 13 2A 43 98 F6 32 99 6D 3F A4 1E 51 C9 FF
 D5 DA 82 3E B7 44 39 B4 BE 66 24 D3 DE 17 61 20
 67 4E 71 09 E0 70 21 4C C3 C8 9F 39 EF 92 13 D4
 A5 4B E9 23 1A FC 7F 4F 30 FE DE B0 EB A2 4D E0
 C9 5B 4E FD 6B 25 03 85 AD DB 48 44 18 5E AC 5A
 63 D0 EC B8 D7 A0 A9 83 18 DD FB 6F 57 25 BA 33
 80 83 AC E4 93 A9 61 6A 2C 08 16 18 F4 8E 8C EC
 22 24 88 AE 95 C4 12 4A F4 54 BE 61 EA 4A 2D 85
 CF A3 9C 1E 97 79 67 61 68 34 06 2C 2D 1C 12 25
 0F 6C 4C D3 97 0A 07 3F 9C F5 F0 25 D4 FB 5E 88
 DD 68 22 DD 2B 09 6D 89 6C 38 57 74 BB 2E E1 8E
 FF 93 79 64 8D DC C2 78 50 8B F9 C0 A0 01 98 2C
 95 A5 28 70 50 B0 00 57 2F EE 73 38 0D B1 16 E1
 D2 2A 58 7B AF E4 37 5F 5B FD C0 F9 3B C0 1D C8
 33 BF DF 07 28 F9 67 33 C9 71 53 2D 54 ED 0C 6B
 EF 1B 34 F4 10 33 28 E5 9E 2D 77 BA DF 1C 40 13
 2B A5 C3 28 27 7D 1B D4 0C 66 06 C8 DB F1 38 94
 33 44 A4 17 F4 B6 FD AE D9 6E 5A 12 32 DF 08 03
 3D 22 F6 97 3E 64 2C 63 E8 E6 52 BF 4D E7 B6 26
 6B F2 38 24 4C 38 D0 C8 B8 F2 77 62 11 32 32 75
 85 96 82 57 36 D1 37 70 06 B4 45 CC 5F A9 45 DF
 E4 6F 87 CA BF 1B 4B A7 99 BD 7C E8 F5 D7 A4 02
 C2 E4 B8 31 33 63 E9 44 B4 C5 7D FD 09 76 1B 4E
 1A B0 26 D5 AB 24 C2 5E 3E 82 58 1A F4 B7 2A A4
 6C A7 02 75 0B 16 62 9B 49 1B 0D F5 B1 6E 77 CB
 B4 26 D2 9C 8E 57 13 7F 59 93 D9 22 AE 7A 7B 5D
 EE 41 26 59 21 FE CE 89 71 36 54 52 FC 32 02 74
 A6 1C C0 34 AE 2D 37 5A DD 7D 8D E5 33 90 80 DD
 75 B2 A7 DC 55 C5 DA F0 0F 0D 60 AD 1C EE 6D E7
 D9 BE AD 8F B1 94 1E 60 03 1C 84 64 27 74 BE 3E
 EF 46 CB 4D E8 1B CD C4 D9 64 D8 2F 22 E8 73 02
 F3 C6 16 03 36 73 95 E1 A6 E5 13 0E 1A B4 92 94
 5E B4 F8 45 20 86 10 C9 10 50 D1 17 67 62 25 82
 B6 E6 09 65 98 93 2F 4A 88 13 B0 98 11 3F AE 0A
 C7 AB 96 D6 28 1E 6A 10 C8 4B C0 8B 96 B2 43 A6
 25 3D 66 C0 52 55 9F E5 C3 87 4F 6B 15 13 92 BB
 54 B1 2D BE FC 78 A0 7F E7 29 6B 71 EC B1 52 C9
 38 47 FC 58 91 22 DE 0C 0A BA B6 4A FC F3 9D 6A
 47 91 64 AE AF DA 10 30 D9 82 6D 16 CB 10 2F 11
 41 96 9B 8B E7 40 02 AB 97 B8 22 7C 94 78 CB C5
 24 18 C1 BF 5A EF 2F D4 3A 2E 19 4B BF 80 50 FE
 78 37 19 EB 6B 85 1B 31 5D 59 53 64 DB C9 76 51
 A6 5A 1A D4 25 AF 3C DB B0 8D B0 42 46 FA EF E9
 E4 07 DF 02 42 70 FA 49 10 76 B6 38 E6 03 38 E9
 AE 45 D8 41 AA D6 CF 4C 82 67 0D 14 E0 1F 97 9E
 F8 17 BB 54 76 5C C2 AE BD 37 E7 F1 80 72 30 AA
 71 5D F5 55 76 AB 12 A0 21 D6 1C 6E 2C B4 9C 84
 F7 59 AE 5D 43 80 7D DD 60 3F 53 EA 4F A4 6E 12
 3A 1B D7 2D 55 74 6C 41 41 5F 7B A8 95 8E F7 73
 CC 4D 00 39 48 E8 48 7A 29 FA D6 D2 3A 53 54 61
 CA A5 B9 F5 91 A4 4C D4 82 9A 5C 07 38 7F 78 51
 80 45 53 5D 0F FC 44 7E C3 D7 FF 92 E2 F1 5A 14
 5F 2C 09 C0 D6 00 8C B1 D5 B6 14 ED 4F 9C AD 30
 FE 29 7E 12 E9 CE 99 D4 9F E0 5E 95 6A 61 48 BC
 56 D9 B2 31 C6 BE 74 FE B6 1A BC 5E 87 EF A3 18
 5C 8A A1 8E 65 34 A3 DA 98 65 DC 71 76 0E 29 DC
 12 CF 37 A5 FE 15 6B 4F 96 A4 F1 18 DA E0 C2 C3
 EE BE 3F 23 D7 C1 73 BC CD FA 17 92 D6 67 03 0F
 79 BB 03 EF 09 74 09 61 E4 D8 79 45 83 91 5B 7B
 59 A8 8F 50 C4 1F F5 42 46 6F 45 A3 FC 1D C6 A4
 EF 6B F5 97 75 15 77 B0 14 39 B7 8C 50 F8 08 9E
 DE 3E 4B C9 AB CA 45 62 13 72 56 8E E2 5D 94 C5
 BF A8 B6 F8 F8 29 C6 6A D3 89 4C 0F 52 AA 57 14
 60 A0 A7 18 80 E3 DD F5 8B F2 17 82 06 CD 59 3F
 71 51 49 C1 39 C4 08 AC 03 C6 2F 96 F3 8A AA 92
 61 53 53 96 F0 40 FC 1E 9D 55 11 53 05 EE 6B 5B
 A9 9D 0A 35 9E E3 15 B5 DB 46 6E BE 5A 1E 1C 5D
 80 68 CF A8 08 8E 9F AD C3 2E 07 F9 67 93 0E 0C
 FD DF EF 6F AB 1C 4C 35 A1 28 9D 57 BB 7B 0F 65
 67 E0 AD 48 5C 91 59 99 39 C0 DD DF 3A A0 0B CD
 0E A7 99 33 E6 8C 28 3F F7 E0 16 41 34 27 B4 95
 2F 46 73 24 EB CF B1 FC 19 AB 8D 2A 66 49 30 8B
 6C 98 58 AE A5 3A E2 46 2D 16 E3 EB CF A2 EB E6
 95 1D 67 D1 92 1D 9A 7C 7E D3 CD 3C BB D1 8B 35
 5D F7 5D 97 F7 5B 1C 54 97 FB 81 9B 14 F6 7E B6
 2B 1E F6 60 71 C0 C2 41 36 43 FC F9 CB E6 01 CE
 6F 30 30 33 E9 A0 F9 C9 EE 18 96 80 25 1A ED EF
 94 1A 91 34 ED 96 09 8E A6 C6 E6 2C 58 E3 2A B9
 FC 71 7E 88 0D AF 26 58 F5 11 73 61 DC 2B 4F A2
 1F 2D F3 9F 53 66 72 75 7D 7F 1E 29 DA 78 4A 98
 27 4B 47 38 26 D9 B9 96 35 99 9C 3D 17 FB 09 EC
 9A 3C 1C 13 FE A3 C3 C5 9F 7F 3D 87 14 D3 3F 6A
 C0 2D B7 0C EE E2 23 0F 7E 7C 06 69 BA 79 2C 51
 C2 AA C2 ED 32 B8 29 7F CF C1 10 B5 BB 75 99 0D
 7F 76 4B 28 9A 86 ED 6A C0 46 E6 52 40 2C AD 3B
 12 1A 98 EC C1 FA FF 54 28 98 A9 31 50 35 51 0D
 3C 85 9C 8F 4B C2 F0 E1 6F 09 44 4C 64 16 6B 41
 C8 BB 67 B4 B8 21 BC 73 F4 68 3B 55 D1 C1 2A D8
 C4 6A 0B 77 74 9E AE A4 AA 5D 66 F0 8A E4 80 41
 43 D1 EF 10 AA 6F 4D E3 B5 57 A2 26 FD 85 83 4E
 7A A2 59 19 41 1F DE 88 05 4B 92 36 3A 9F 7E DE
 9A 61 61 FD 2D A9 DF 99 7C E4 4B 4A D5 FA C0 1B
 DC F3 4F 26 31 A1 1A F9 F1 11 5F 26 3D 18 0D CF
 50 F7 82 53 6F D3 BE 5F E0 55 12 5B 97 EA 79 6D
 57 89 93 F0 1D AD E4 95 5C B3 3C B0 96 E0 57 C1
 FB 9D 06 6A 32 B3 A3 CE 59 33 AA 39 1F C2 E3 A3
 5C FB BF E7 52 FF 58 FF FD 18 52 48 2B 96 D4 B3
 D4 26 39 31 1D 73 B0 56 3A 89 60 14 58 2D D2 FE
 F2 38 9E BD 7E D3 F4 CA 70 0A 6E A4 C0 3F 87 F6
 42 3B 42 40 12 99 A2 6F B1 43 D2 18 B8 F0 46 0B
 9F D9 05 7A 13 B5 5F FB 87 E2 B1 45 99 94 7D 76
 2E F3 E9 E6 93 35 13 E9 C4 CA 7B 1F 98 84 D4 8C
 6F 32 DB C5 C9 EE 48 CC 7D A9 8C A4 E3 61 FE 0E
 7A 04 3A 9E 02 36 5D 62 3B 18 4F 5E 18 23 12 A4
 9E 3F C3 3B 1C E6 50 C4 A3 32 57 6C 97 8B 31 A6
 CC 11 13 83 F4 8F 73 B1 6F D8 22 CB 7C E9 C8 9B
 A0 87 9F AE DC A5 38 89 FA 19 55 BA FF 44 93 6B
 8A 5F 83 A8 DB 84 E9 36 C4 59 A6 A9 EF B8 A8 D5
 45 94 8D A4 F7 66 07 56 83 53 A2 15 9B 82 54 50
 14 81 E1 98 05 A1 D7 5B B6 7C 95 BA C3 D6 D2 8F
 B0 6E E8 4D 5B 85 19 CF 2F 28 EA 68 66 D8 5E 98
 14 C1 A9 8D 17 0E 9A EA 82 CD 6D AF 54 BD 2B 08
 21 5D D1 2A 03 E4 03 33 03 66 4C BF 0D E1 7B 8A
 7C AA 97 1E ED 03 9F E7 A6 9D 1C 33 08 8D 73 8D
 D3 85 BF 51 03 AA 21 47 D7 73 88 FB 68 54 0C 14
 86 AC A8 C7 24 7F E9 A0 A4 A3 CB FF 0A 5A 6B F0
 96 D5 01 E7 BC A4 FA 8B 46 7A 00 EE F6 30 24 6E
 17 27 09 F9 1C 30 89 4B 49 74 6B 85 5B F0 76 21
 0E 1F 14 A5 A3 96 6C 1E AB 51 BF 32 94 0D C9 27
 DD 90 59 36 CF 05 EC B6 F9 22 99 99 07 25 DD EE
 92 0A 88 42 FC FF BA A1 3C CA 7F 92 64 62 70 D7
 8E FB 90 65 83 B1 1A DB A3 87 86 40 E6 43 F9 FA
 44 7A AD 59 3E 68 09 25 37 00 75 56 66 43 54 84
 9D AA 15 FF 99 4E 8F 7C F1 65 0E 32 52 60 E3 C0
 0A 5C 0E FC CF 3D 54 B5 0E 1E 25 8F F6 BA F1 CC
 BC F9 71 D7 C0 E7 35 48 85 E3 7E A8 16 D4 8C 0A
 29 81 20 7B 74 65 99 64 AD BA A9 E2 A7 7A DF A9
 E9 7C BE FA B2 FA 0B 10 4A 22 29 0F 86 DE 23 54
 81 9E 2F B8 DE BB 96 74 02 37 3B CE C3 70 50 78
 5D 58 3D 2D C6 2B DD A8 63 FF 06 40 44 D0 81 C6
 46 B6 F5 B6 E0 29 53 96 A6 A1 22 0C CA 46 4B 7E
 68 B1 9C 0E DB 62 82 81 B8 1F 63 19 04 84 68 1D
 4B E9 05 97 53 BB B2 1F 80 B1 27 CE 69 35 0B 21
 92 3A 4A 70 4A E7 65 8E D8 41 C4 CE 00 65 60 B4
 22 A2 EA CD 44 5C 6E 08 A4 91 63 13 36 3F 4B F4
 4B 7E 0F FB CF 7C 33 09 1D 0C AE D0 C6 83 98 55
 31 64 C2 2F 56 76 B5 E1 DF 5F C8 94 EF 2E 11 13
 B6 D7 68 35 AE 6F F0 1E 8F 59 17 3E 5B 79 5C 3F
 65 DB C1 5C 95 B3 18 A1 EF 65 7D 5D F1 3A 5D E4
 34 D6 CE 0B 15 A8 53 CC 05 E8 59 46 40 96 E4 76
 15 1F ED D4 27 43 C1 26 A6 BB D9 32 28 13 7A B6
 AC 95 95 C9 F1 C2 3E B7 0B 6B DB BB 48 84 5B FC
 9E EE BB E1 BC D0 70 F4 7D C6 DF D1 33 C3 33 7F
 55 E9 CF 01 6D 61 1A 0F 37 74 99 B2 6F 17 7E 2E
 B3 1E C8 9E 83 C7 1C E1 FA EE A4 6D 05 50 72 46
 A8 27 29 59 45 C8 B7 9A E2 50 C9 A0 01 2E 59 99
 0C 63 75 D7 54 25 C0 9E 80 B1 BC 15 78 56 90 B2
 37 D6 C8 52 17 84 B7 51 FE A3 86 EB 94 15 33 07
 40 59 95 29 10 81 CE F0 30 84 F7 7D 51 12 52 20
 99 31 F2 7D 8A CC 08 9D E9 BE D1 6B E7 59 0D 6F
 AA 1B 89 EE DB 47 E8 A9 44 3F F4 F9 28 31 F4 08
 B9 78 54 A5 AB 56 FD 04 EF E0 46 81 ED 58 EB 3E
 58 DF F7 CF 97 EF FF CF 9F C6 8B C4 C3 A0 55 19
 A8 96 FD 72 C8 C6 67 40 3B 89 0F B7 27 FC C8 AD
 A1 49 EB 29 2A 5A D3 3B 9F 24 B8 48 49 BA 35 F1
 B8 08 43 F8 52 D0 26 33 42 69 7F 07 4E 2E CF B9
 6C 76 94 45 97 03 9D 22 A9 27 6C F8 D1 77 B1 30
 CA 39 D9 5F 63 23 AA 11 3D 0D 1C AD 65 25 B9 8A
 FF 5E B5 8A E5 E0 64 B2 4C 5E 80 3C 45 55 E4 6F
 53 65 75 B2 08 45 F2 0F 72 D2 3E 4A DF 75 0D F7
 75 F3 DD CF 48 24 C3 BE F7 86 3D 67 C8 57 C3 AA
 64 8B FF 98 70 8A 50 B3 2E D0 58 26 2E 2A E8 36
 A0 AA B2 40 A3 FC C7 B0 46 25 3D 9E A0 EB 77 B2
 E6 EE 4D CA CF CF 3B 88 37 F7 66 EA 80 40 90 F3
 E7 50 04 93 E6 52 E1 62 FF DB 10 BB 40 23 F7 EB
 E3 89 DD 0F 05 5E C2 3D F6 C9 5F 8D 7A D9 B5 1A
 AF 32 84 0F 78 C7 5B 47 FD 42 9F B1 C4 AC FB 57
 66 82 49 9E EA 51 67 0C 77 85 65 CD A8 E7 F1 E8
 08 D5 E0 8F 3C 04 B7 D3 13 C0 01 17 8C 4C 48 9E
 93 EA FA 3C D8 3E 5A C1 81 25 AA 54 B5 43 8F 7D
 76 B7 8D 13 D2 0E A3 FC A7 9E 37 09 4E C9 74 D0
 11 DC 50 73 F4 FA 6B EF 00 13 1F 46 F5 0D 1C E3
 B4 67 57 4B 3F FB D4 B7 24 29 36 C8 F0 EA B0 45
 8E E5 46 C1 8A 18 6C 02 A8 6D AB 80 B8 84 A9 47
 CE B6 2E 2C 69 42 C6 7E 74 1F FA 2B FE 68 9C E3
 5D 56 0F 05 FD 14 7A AB 2E 82 7A 34 E0 42 32 DD
 A3 13 54 34 A1 BF EB FA 90 F2 95 AF 5F C8 10 01
 6F A5 1A 26 33 5E DE A5 FB 2A F6 EB 76 AE F8 26
 39 83 63 F5 89 15 0D C3 A6 95 CC 9D 93 23 F1 B5
 49 DC 02 86 2C E3 A3 D4 8A 70 8C C1 E8 26 D7 53
 A3 51 02 6C 09 AC 89 E1 FB 81 31 0F 3B 0F 62 10
 C2 5F 4D 1D E2 FA 15 EA AF 5E FD 60 44 9C 40 5E
 09 E2 81 9A 0F 7F 60 8E C7 2A 12 30 94 BA 86 B0
 97 C4 10 D3 CD D9 37 88 14 51 5B D3 7F FE FB 87
 5E 78 08 99 95 07 F7 80 88 14 0F 7E B4 D9 81 C3
 43 3E AE 9D 7E 88 E9 38 CD FF 31 14 D4 C7 0E 1F
 14 CF E9 6A 16 F9 0A 05 F4 95 EF 26 E5 83 EE AF
 5D 21 4C B4 91 F5 5B FB E3 F1 1F 9D 45 FA EF 20
 3C 94 CC 1F 58 0C FE D7 83 1A FA 75 14 03 14 45
 A4 25 27 9A BE 35 51 24 B5 0F F3 AE F8 C9 2C 53
 3F 2C 3F 5B 49 A2 4D 45 DD 71 1F 7B 66 9F E8 C3
 9B CF 80 40 ED 04 EE 5D D4 D0 EE 10 3F 9A 73 5E
 E4 26 B5 42 BB C4 3E 4B 7C 43 BB B5 ED E4 40 76
 39 99 E4 17 77 5D 3C AB F5 00 05 E8 89 8F FC 87
 13 B1 26 C4 96 F6 59 32 92 82 F3 EE 3F 22 90 48
 DE C2 62 FA 85 0E 57 CF E6 35 16 B3 EC F8 D0 1C
 1D 21 B3 3A 35 19 C6 A3 13 A4 E9 E0 72 60 10 27
 8E 2E FE 97 93 29 28 59 48 C7 44 FE FD 43 F9 F4
 76 9A 11 FB FD D6 58 8E 11 41 01 A4 9B FE C6 A7
 43 72 C2 AE C8 77 0B 3B 8F 31 D5 AB 85 1D 90 0C
 68 87 9B AF 3E 1A 1E 7C EB DB 91 3C F4 EA 35 FA
 EB AF A2 22 9E 0E 37 A3 95 5D 23 AE E0 BB 48 94
 60 16 C3 35 50 E0 4E A6 DA 2F 0F B4 36 C6 51 AD
 C1 54 85 A4 EE EF 84 BB 79 1F 4B 1A 7F 9A DD 68
 3A 9C F6 43 FD C8 01 BF 47 0E 1B FB F3 0B 94 D7
 0B B0 F3 57 4F 33 CE F5 14 80 D6 3C 61 1B 47 EB
 83 18 6C 86 B1 6E 27 EF AA 5B B4 46 8A E2 B5 A1
 5F 05 D9 4B BD 8F 50 BF 52 AC CF FE 00 D7 C5 82
 AC DD 83 9E 85 3A BC 7E 32 90 B9 3F 13 B6 5F D6
 C5 F0 D2 3F 68 BA 77 09 81 63 25 54 C1 16 B5 A9
 51 92 2F 70 BC 28 35 CA 57 F3 11 1B 67 7E B8 A9
 57 0C 71 B7 FA E3 2B 3B 53 12 2A DC 24 0C C2 0E
 67 2B C6 B4 B3 E8 BC A6 A2 A0 B8 4B 85 A9 65 CB
 5A AE C6 E8 30 A1 01 86 FB 9A 34 E2 63 94 63 76
 E4 97 ED B7 D0 E0 21 6C 63 E2 CD 3C 37 38 88 2A
 A0 85 94 A2 E1 84 9C 54 54 C7 E7 B3 A8 6E FA A4
 91 69 AD CA E6 8F 45 B7 0E 89 24 42 B9 EB BE 43
 B3 2B D5 84 D0 5B 83 16 22 44 33 3A 26 2D 8A 40
 61 A7 3D 3A 02 6E 4C 72 99 0F 2B 9E FC A4 22 2D
 6B 6E B1 37 84 5E 62 E1 96 48 F0 E5 26 10 05 2D
 6F 4A A8 80 2E B4 2D A7 A5 23 A9 1C 3D D5 02 88
 B2 44 5E 9C 49 FE 2C E0 D7 4D 6D 5D 43 0A 30 72
 B8 91 E8 7F AB A2 AE E8 BF 62 18 F9 1B D6 0F B4
 6F 15 EF 5F 9F 3B 03 74 18 91 EF 24 6D A9 87 2C
 6E 69 AD 8F 64 D1 97 E0 DB 1E 4E D6 5C 03 77 E9
 72 18 EA B5 D6 58 E0 CA 2B 2D D4 0A 6F 7A DF 38
 99 28 88 18 43 70 5C 1D F6 22 98 67 04 14 CE 44
 11 B2 F4 2B 3F 17 71 92 0E 4B 0A C3 59 9E A0 AB
 0E BD B8 E5 FF 96 9B 25 B9 03 DA D3 E3 7B 31 27
 97 93 E2 6A AE 74 4B E7 26 D3 E5 36 05 89 F6 66
 87 ED 72 E2 94 E2 20 18 B2 CE 7A 5C 8F 56 E8 98
 DE 96 41 04 9E 11 C6 95 35 D6 AB A8 CB 99 75 84
 EE 66 2B 86 6C 13 0B C5 8C 3C 74 1D F0 E7 16 AA
 FD 3D 32 DF 73 42 6A 3D A8 BB 2B B0 82 DF 0F 09
 9E 60 3C 97 52 DD A2 FC 64 8E D3 89 EB 01 25 2A
 AE 82 84 54 96 BA 7F BC 93 26 84 72 6F C7 BD 1B
 CA 32 0A 1A AD 30 16 66 4C 60 82 43 3D C8 67 00
 9F 9F 0A 8E 6A 58 9B C8 8B 16 F9 BE 7C 0A 20 D4
 3B 4E 8B C5 CE 7C 5F 7A ED 96 1A CE 02 EE 0C 38
 44 AA 1E 91 C5 DD 6A 66 62 C9 62 18 A6 A7 6D 27
 9B 92 4C D3 FB F1 5E A7 05 B9 9A 68 D6 8C F7 9A
 9C F3 E4 DD B3 D1 56 4E E6 A8 53 49 3A 17 87 8A
 AA 82 FB 63 49 82 14 77 5C 17 80 DC 10 AB C0 89
 95 46 8D D9 9B 28 3F 58 C2 04 19 B2 53 2E F7 1C
 62 90 D4 E8 9B AF 62 19 68 5E BE CB AF B6 12 1F
 A0 1A E5 CF 71 3D 83 FE F7 40 9B 6B 5C E1 94 C8
 45 9F AB D4 2A 9E A7 0D 6F 49 61 C9 FB AB F6 92
 42 A8 5E D5 5B 2F C5 35 F6 C5 44 22 69 48 CD BE
 E0 84 5A 8C 9E CA 6C F4 2D 59 72 EB E7 B7 FD 05
 0E A6 89 BB 92 E9 48 0E 32 69 11 3A 71 F4 A2 64
 2D 2B A2 B4 32 E3 98 20 FE 1B 51 3A 60 12 9C 4F
 CF 70 0E 5A BF 6F CF 3E F0 45 F0 BE 81 61 FB AC
 61 CA 4A 99 61 2A 54 EE EC 8E B1 5A 05 6B 1F 1A
 4F 94 31 9C 0B CA B6 C4 9A E5 A2 A1 D3 59 F7 16
 4A EA E3 15 AE 45 89 B4 98 B7 52 88 30 E2 C3 02
 14 F4 BF 25 31 C1 25 12 41 A9 90 8B 2C A1 2A 25
 D8 80 9C 6F BA F9 94 10 3F 96 6D AB ED C8 5D F9
 8B BB A0 B7 B9 D3 EC BE BA 12 B7 FD 94 C7 0C E7
 90 77 0F 7B 0F 50 A2 49 C1 75 7A F7 58 47 D6 21
 42 BA 36 51 65 2D F2 F1 84 5C F0 A5 B8 DE 1D C8
 C8 FE 35 94 1E 6E D6 92 38 13 AE DD DD A0 B9 6D
 39 26 8C 0D B3 00 89 8B 2D B4 39 AC FB 70 3A 44
 C1 EA EB 66 40 14 76 7B 8E 98 B4 A6 6D 2F 08 D3
 02 B4 F5 2F C1 8B 38 B3 93 D8 24 4F 93 FB 27 46
 7A 35 AF 78 14 2E 41 B8 B8 15 65 16 D3 7B ED D0
 3E 78 3B 2B 38 62 AD 93 47 9E 48 55 B6 5B 3F C0
 FD 03 FB 64 24 D3 61 C7 A4 5C 9E D8 43 A9 6B BF
 70 FC 09 22 77 5F 01 22 FA 1B 86 F7 3D 15 3F F5
 16 62 F6 A7 45 CA B6 CA FE 24 E7 47 91 62 21 85
 B5 23 41 37 94 13 AA 75 A2 EC 45 95 99 85 7F 29
 E6 3D 0D CA E0 5E 6E 52 2C F4 A8 96 02 5F 73 22
 9A 49 90 BD 35 59 F8 5D 0B 44 86 37 51 6A 38 E3
 DE E4 EC 19 4D ED A6 49 73 26 A6 80 81 1E F1 41
 76 BA 74 45 8E 3C 1A 46 F5 81 5D F0 FA BD 05 31
 97 E0 B7 24 84 94 A8 85 8F 15 E7 5C E1 45 3F 87
 1C B6 9F FC E7 60 C9 37 06 C3 23 A9 58 7E A4 51
 AA B7 F1 9C 2E 0E C6 AF E7 1A 28 9C 74 0F AD 64
 9D 65 92 5B FE DC 22 69 D5 09 5F 26 12 36 BD 33
 83 84 E5 D0 C9 4A 1A 60 BD BD B1 8B 53 87 1F 8B
 55 E4 69 A6 F1 84 00 05 52 A2 52 E6 64 D7 16 B2
 1C 9D 3B B6 BD BC BB D4 E0 EF 77 B7 92 B5 28 B4
 42 41 CB DD 7C 42 1D 27 9B 09 31 A2 93 1E 25 DF
 4F 5D 68 B6 B9 1A F2 3F 78 5B 0A 1F F1 47 B1 F2
 63 DD 09 EB 9F C1 9E 1D CD DE BB 3E 71 4F F1 D3
 F5 CD 9E A0 48 DA BE 3F 48 12 DE 6E D8 C3 D6 49
 15 56 15 E9 A2 07 A4 B6 55 88 FB 64 3E 22 51 AE
 54 9A EB AD 44 92 5D 43 5B 11 9C E2 14 33 EA 96
 C4 79 CE 23 CD 52 08 2C 3F 94 48 CA 0F 4D 5F 0E
 2E 95 79 93 E2 5C 8B 7D A3 50 39 41 6E 3D BE F8
 2B 3C 26 27 67 00 C0 B0 78 17 79 D2 CC 5C 09 A3
 E7 48 76 E4 2A F0 04 BA 34 41 5B 3B FD 14 E5 1F
 79 6F 63 F7 4F 05 FF 93 60 44 05 E7 1C 08 DF 96
 75 EA D9 2B F6 F1 CA 83 5B 2F 02 05 32 04 C4 EA
 FC 3B 01 5A B1 30 1F FE E4 E1 F1 C0 24 57 FE AF
 D7 EE FE 93 EE 7E B8 9B FE 1F 24 28 63 15 1B F7
 82 CF 40 67 1E 04 2E F9 8A 7E 7A 81 41 59 AF AC
 12 1C A9 EB 21 7F 55 41 BD AF 68 A7 27 CE 4B 8B
 C9 40 7B 27 9D F8 78 25 63 93 F5 70 21 0A 2F E8
 FE 4D 86 6F FA 50 14 D8 1F E7 36 00 5C 59 1C 0A
 CE 5C 02 AF 14 17 52 48 DC 58 27 D4 BD 2E F1 44
 E2 07 FE 37 36 04 40 BF C5 DA CC E9 4F A2 4E 4E
 05 21 FE A2 E0 C0 4F A7 62 8F EE AE BA 53 AE 5A
 73 63 DA E8 13 31 4C 78 DC 66 CF 0D 3F B3 92 BE
 2E A0 66 3C 98 F5 E2 C7 8E B4 F3 C3 42 98 C5 16
 96 78 A2 BA 9A 4C 97 A1 E9 E8 4E BD 9F 9E E1 E3
 16 E4 C1 FE CE 9F 21 85 75 1D C1 9B 3C 70 2C 50
 49 77 4A EC 20 8F 16 14 83 B6 76 1D 9C FB B5 6C
 68 4C 90 0A 7A 01 C8 A2 5F C3 B1 5D 51 C9 FD 5D
 42 DF B8 0B 42 6E A1 09 81 50 2C F9 27 B6 65 BC
 36 B5 54 C2 09 83 F0 EC C9 00 D3 0C 25 88 14 07
 88 18 12 35 83 C5 22 47 2A B7 8E AB B9 72 13 A7
 14 34 12 8A 9D F8 A4 94 3F BC F3 47 3D 7C D9 36
 4B 99 D4 48 20 B8 0F 28 E6 7F C4 66 9D FE CF D8
 3F EF 23 09 43 16 C6 6B 15 6E 0B BF 76 7D 3D C9
 96 63 86 65 7C B2 27 5F F9 CD 08 1E 00 61 42 84
 9A 0F E0 1E 83 83 DC 33 6C 79 F8 91 70 7B 9D 9E
 14 89 BA 7C 80 46 4E 23 06 A4 64 A3 11 BB 64 E7
 26 50 F7 16 46 56 28 84 06 14 0D F6 36 69 3F B2
 B1 2E 45 E4 D4 6C 2D 3B 5D 3B 65 B0 A1 9A 13 5F
 F6 EB AD 70 58 39 47 C8 39 FD 50 02 3C 9B A9 15
 83 F1 88 6B 85 57 63 58 A3 4D A9 33 D7 B8 C1 E4
 6F 63 CE 73 F8 97 EA A1 85 7E E5 2E 02 F5 D8 E5
 46 03 BE A9 8B C7 92 41 FF C1 6D 6B 5C F6 DF 06
 98 53 8B 0A B2 6E A3 AA FA 3D 9F F7 4C B2 2D D7
 DD 4C 2D 3F 97 19 F6 DC AA 86 E7 7D F6 00 D3 BD
 91 76 F2 57 62 8F C2 E7 6F 12 DB 98 F5 46 60 9A
 D8 F1 CF FA C1 E2 2C 6F 4F 75 8D D1 B0 98 80 A8
 DB AE D9 29 43 3E 2A 2B 92 DD E8 57 88 76 61 C1
 4D F8 3F 56 A8 80 55 74 F4 F5 88 B6 20 DF C9 12
 B3 60 95 75 F7 2A AF 9F 05 C3 97 22 62 49 7A A9
 EC 53 07 E8 A7 29 84 E7 08 63 E7 08 9F 7F B8 BF
 CE 5A 58 E5 BA 2B 26 56 F7 05 06 4E D8 16 0B A7
 10 9A 5F BA C3 83 05 F8 08 3D 7C E5 0F 0E F2 D5
 96 DC 06 D1 41 54 D4 3B 1D 1F 6B 0C DC 2A 83 60
 1E 58 EF F3 7F 37 4D DA 6E D2 B1 18 A9 5F B2 7E
 92 EA E9 40 B6 84 82 7F 35 1D 23 EE 73 9C 25 FC
 AD 88 7D 24 4B 83 C2 2B D8 42 23 2B 8C 49 87 69
 8E 06 28 E6 FF B3 DA FB 2C 4C FB FE 19 06 8F 4F
 B8 77 1C 55 CD 70 86 BE 79 79 3F 61 A0 D2 9E E9
 CB BD 85 67 DD 3E 8D 97 06 24 EB 82 E2 E9 4B F1
 2C 78 03 D4 F0 BA 26 68 5A F3 A1 08 65 C4 B7 69
 26 82 32 82 84 E1 B0 20 B6 6F F2 75 49 8C A1 DB
 AB D9 54 13 35 7B C1 65 D0 46 0B 9B 08 C2 C8 8F
 8C 6B 11 48 11 50 43 EC 51 B2 42 50 0B 85 8D 31
 BE 62 50 13 16 F3 80 21 EB 71 BA 65 37 68 5F FB
 54 5E 66 47 B8 10 10 16 2B E1 87 F6 59 23 7D C7
 0A 35 C4 59 4D 19 FA 1D 69 FD 41 27 F2 67 5B C0
 09 99 BF 6B 67 C0 83 59 CD 96 DE 95 E4 98 AE 8A
 C7 FA 80 D1 61 C3 7B DF 97 0C B7 FF 35 A5 8A A2
 22 51 F0 DB 78 DE 82 BD 7E 68 88 17 34 2E A0 07
 24 D8 39 6B FD 79 77 53 70 4A FC 39 6B 0C AF B3
 76 4D 38 8A F8 E6 E9 C1 2D F0 93 DB 91 5A 82 43
 49 24 66 A7 66 33 3E 7F 8C B0 B1 74 A0 17 FB F2
 6B A1 78 B8 95 0E 48 A5 48 9C 90 7C 0D FC F7 88
 2A 90 B3 3F A5 77 1B 33 16 99 23 5F A5 4A 1E 02
 BE F2 87 DB 05 7B 57 7D 6C F7 6F 9A 64 2A C1 3D
 07 81 E2 23 B5 38 17 10 88 C7 12 D0 83 8E 92 97
 E5 85 A5 DE A3 FB D6 D7 1F A3 0A 5D 50 52 87 A5
 35 28 4A 9E 1A 28 FF 1F E7 60 D7 86 4E EB 86 BD
 3B 7C BC 77 CE ED 11 4D 56 E5 25 48 8D 29 14 1F
 09 11 6A B1 74 59 C1 DA EF B5 42 F7 90 28 32 75
 51 5F 7B AE DB AF 2A 31 21 53 B1 18 0A AC F5 A3
 86 69 16 1D D6 A9 62 FB 24 4D 53 02 82 85 3C AA
 51 D2 88 EB E9 6B D6 E2 E4 C3 40 98 9B E8 AA BA
 CB 8C 31 E0 81 79 D1 EE 0A C5 2A E5 98 83 CE 93
 55 03 B4 AA 04 65 78 92 88 F6 76 4D 10 12 70 E1
 62 FE 8A 39 DA 4B B8 E9 00 40 14 C6 E8 AF 72 FC
 EB 01 59 16 EB 89 C3 CA 8F D9 A9 72 70 F5 3B C8
 EF AC F5 D5 E9 DD AC 52 23 37 02 87 23 CB 2B 4A
 86 55 34 10 E8 72 69 86 F3 FE 9B 6E A4 EA 76 FF
 43 F7 A9 87 E4 2A 56 63 CF FB 54 5F E1 01 64 E0
 57 25 50 DD 8A 9B DB DF 99 A5 93 1B DE 06 76 85
 9A B2 1F 83 2F 21 A4 21 A0 6C FA CA CE F0 37 22
 78 D6 C7 D4 3D 4F 37 BA 99 EE 65 2A FA 19 C8 E2
 C5 D9 67 1B CD CF 2B E7 75 32 8C 86 46 9B F5 35
 22 92 77 F3 93 09 EA 86 5B 3A 7E BA 21 75 FD 49
 35 25 8D BB 79 6A 71 09 E3 5C 2D AD 42 7F 91 40
 D0 EE A9 07 62 12 4C 6B A2 00 14 31 AB 63 A1 49
 B7 44 A5 1E 38 D9 FA 11 63 4D FF EB A0 04 4F 8F
 8B 00 95 B7 E3 3B 9E 2F 6E 7F DA BE 5C 1A C1 D8
 8D AE 20 58 10 FD A0 DE 45 AB FD B8 64 74 81 68
 7D 47 6A D0 82 3A CC EF D6 ED A3 D8 08 E7 7F DE
 E5 6F DF 94 C5 3F 21 01 00 09 9C 77 FA B6 CB A7
 BB 5C 82 70 16 59 C8 B4 E3 D4 D8 4F 7B 1D 97 6E
 71 EF 8A 84 3D A4 87 E9 14 24 F7 E2 86 D6 13 DE
 6B 15 EB 87 16 7B DC DC 44 FF 42 AF 10 53 42 30
 D4 4E DA 27 EA 64 7A EB F9 40 11 02 A1 7D 21 C9
 10 CD C9 88 D7 F2 A9 22 F6 69 36 83 82 9B FB 88
 C7 E4 60 53 65 FD 4E 84 E7 68 E3 06 14 FF 06 B3
 B7 3D 1B 28 85 E8 F6 DC 0E E6 70 22 36 72 71 64
 94 13 F6 DC 14 65 0F C8 D2 DE 81 60 09 1F 78 99
 23 BA 6F F0 EB C2 91 6D 8D B8 22 E2 CE E8 E9 7B
 17 C3 0B 8C AB 4D 5C D9 30 AB BD A5 B2 BF 10 86
 05 B2 75 DE 77 D1 84 9C 4F 5A DA 02 EE 7D 08 B9
 C6 2E 7F DD B5 AD 26 5E 04 5C BA 5E 6A 8A 06 8A
 C8 47 44 D0 30 79 B6 50 5C BA 7E DD 02 53 DE 3F
 D4 9F 20 20 2F E6 A6 D5 06 3D 30 8C 50 EC C7 DA
 44 F6 9F BB A4 EE 41 AE 7C 4E B6 05 2F D3 7D CD
 DB 9A 13 08 DC 1F 02 19 F4 40 E9 FC F1 05 73 0C
 FA 04 D2 7B A8 69 7E 1B 38 7E 0E 80 3D 45 47 2D
 1C 9A E3 7F 1F C9 65 1A 64 31 53 9D C6 99 B7 D8
 C1 D3 01 7E 16 6A 22 D9 88 0D E6 84 CE 02 0C 18
 57 14 22 DA 49 FF 97 78 98 FE FE 54 C2 6B 9C 77
 98 EF F9 34 45 D9 EE 9A C4 76 AF 10 35 D5 9C E3
 E1 D1 E1 CB C8 81 78 7D 85 A7 AF 9A D1 5B 00 96
 1C C6 82 18 65 54 BC 29 CF A4 3D 5A B3 4E EA 13
 0F 4A A0 31 2D 38 30 AD 13 52 11 50 75 C8 AF 4F
 DA 2D 39 82 A2 03 0D CB 0F 72 03 8E EE 38 18 62
 6F 1E 13 C0 8C EF E5 AE F3 20 20 BF 3C 72 AF F9
 E5 01 54 0E 8E 41 07 80 B2 94 1E D9 19 1C B1 01
 70 37 7D 9D 37 0E F8 DA 24 4A 6E 39 0D F5 8C 4B
 20 31 FE CD 2B 34 15 53 C4 41 FA 04 14 1F 30 A3
 EC CE D9 49 4D 64 A7 53 81 FF 89 78 55 BF 5C F5
 7B 80 8B 3C EF DE B2 02 FB BE 8C 31 FE 2C 94 CE
 CC 1D 09 C4 90 08 99 41 1A C4 6A 1F E9 3D 15 A9
 7B 8A A7 A5 DD F0 BA 6A C8 76 44 A5 D9 0C 0A BA
 C5 51 8B 00 0B 3C 2C 93 21 D8 4A 79 42 33 AA BB
 7F 30 4F CC 40 7E 3B B1 16 73 2F 0F 23 D8 8D 06
 1B C7 BC B0 D0 F6 B5 64 3F 6B B8 51 BE 2C 56 42
 D5 40 BB F4 DE EF 16 F2 3E BA 94 81 4F 6E 8A 24
 0D CA 9C 2D 7E 16 C8 1B 92 39 1A B1 9C A0 02 4E
 08 EA 16 1D DC 03 15 C2 9C D4 0F DE 87 F3 AF 24
 F4 22 A8 D2 A7 25 DE F7 26 82 B1 E5 9F 15 16 FA
 60 26 12 D4 96 B2 FE B3 10 D7 F4 BC DC BB F8 CE
 1C EF B3 2D 83 D4 26 CC A5 2D D3 EA 3A 15 50 01
 07 71 5F 22 79 B4 E9 11 FB 0A F2 E7 98 02 32 39
 0A B5 16 1C AF 0D 7F 13 3E 6E 90 C5 DC 0F E0 F6
 70 6E DA 41 82 39 0E 0B A0 FC 03 B1 F9 6F 15 D9
 7F 1C 17 F8 73 14 14 DB CA D0 C0 C7 3A 8A C5 F6
 05 D2 D1 20 43 E8 7E 49 79 E9 4A 0D CB 85 E8 50
 11 A3 D2 09 20 C4 57 0E C1 EA 4E 87 33 BC C8 45
 06 74 EF 60 55 16 E7 1D 1D 9A F4 44 E2 1E D4 D0
 D3 25 D7 3A FA 65 EE 57 6F 4A 16 A7 6B B5 05 21
 9E F4 D7 49 EB 3A C8 01 A2 BD 63 A3 3A 20 AD 2E
 C5 67 A2 81 F3 45 A3 B3 85 EC F6 11 2C 17 C9 6B
 41 76 BC 85 75 37 0A 6C 79 23 EA DE EA B8 25 1A
 D9 B3 1F 99 79 93 A5 64 9E 6D 08 00 86 63 36 37
 9E AD 0B E6 C7 3A 90 B7 33 C2 45 F8 25 0C FE 10
 5D 24 D4 E9 7E F5 E5 CC 78 61 1D FB 85 9E D3 16
 B7 35 4B 0A 9F 13 34 0A 4D 83 72 25 DA 14 91 AD
 A8 F3 F2 4F 73 63 B2 68 AE 7C 7F 1F 67 4D C1 53
 8D 5C 47 22 F2 2E 2B AA 42 64 79 5D 6B AA 8D C0
 06 BA 39 5A 80 BD 4F 3D F0 E9 91 2F 1E E8 A4 1C
 ED 89 49 C9 86 73 EF EB DB 71 C6 54 40 1C E2 BB
 22 78 7D 89 4E 06 2A 20 1E F8 78 DC 82 FE 82 92
 1A 68 0C 86 58 CB B4 C6 6B 75 B1 57 25 A6 92 F0
 C8 9C 90 C6 81 9B D6 9A 0E BC 68 07 B8 AF 29 E1
 EB 90 67 08 DD DA D7 D4 07 64 C0 F6 9E 2D 82 D5
 AF 0B E5 87 4F BF 0D B6 BF CA 85 48 5B 26 98 04
 95 C3 40 F8 56 DA 53 15 AB 39 A3 1D 00 99 0F 5E
 2B 20 DE 3C 95 68 D9 DA 86 5E 12 7B 70 B6 7D 09
 AF A8 51 D3 CA F2 BF 2E B0 3E DA 9E 09 B8 95 FE
 87 60 A0 90 E2 99 08 87 68 60 EB 3E 50 19 93 48
 96 4B DE B6 F8 F9 65 06 BF 59 50 AC 88 26 1A C7
 CC F2 87 90 08 D6 18 40 DD 7D DA EA F5 FE 21 B1
 EE D8 71 AD FC 6B 17 15 15 EF 80 F6 8E A7 4B 81
 D9 25 7A 97 E6 2C D9 66 EA 98 8A 2A 6D 8F 1B 27
 C4 EB 95 92 95 8A 98 EE 0F B5 DB 9B 18 BC AF 36
 AA D9 2B 03 49 4E 58 2D C9 04 AE 8E 3A 46 CB CA
 F6 F5 4F 61 50 2F 84 63 7A BD 43 6F A6 89 8D A9
 DF 96 CE 4A 9E 3D 19 84 04 1A F0 C2 6B 3B 57 13
 B0 3A CE D1 19 CE ED 2D 49 1C 45 7C 73 B0 86 1A
 92 8F DE 1A 7F F3 7C AB 2F 08 85 BB EB E9 69 27
 F5 AF EC AE D1 79 BE 04 89 EB 14 1C 92 7D 0E B8
 ED 11 ED BE 48 F8 D4 D5 6F 15 FF 59 5B 5C 0F DC
 22 EF 1F 3B 81 DD DF 0E 84 1C D0 52 B2 47 35 89
 4C FB 7B 57 77 25 BF 57 AC DD 02 E5 EF 67 AE B3
 3F 95 A2 C3 26 11 75 18 72 BA E5 F8 5D 61 64 2D
 0C 62 E5 48 E4 21 92 60 07 89 D2 B4 90 DD 79 2A
 06 73 BE 42 1D E2 AC 36 8F 6D 02 D7 D1 B7 5F 46
 DF 49 7A CF 19 13 94 33 C9 96 9E FF 40 8A F4 F2
 26 A8 6E 66 40 1D 42 EA EE CA 21 61 4B 59 CA A1
 55 17 2B A8 41 A7 A5 6D AD 5B 3B 8C 04 02 CE A4
 DC 94 79 C1 BD B8 00 B1 83 0C 4B 41 DE 7F 26 C8
 FB A9 81 D4 8B 80 25 3C 1C 6A C5 C7 44 64 0C E0
 01 15 5E 58 67 8A BD EE 4C 58 B8 A8 82 EF 70 7F
 0C D5 BF 7C 3E 7A BB 0F CB C8 FC 0A C0 37 90 51
 DA E8 6A 32 41 A2 12 0F CE CF C3 31 F3 42 E8 30
 43 37 C2 F5 57 78 2C 4F 81 F7 26 C4 4E BE B6 1C
 63 E3 19 62 66 C1 1E 04 41 18 CA 9E 93 22 29 F2
 1F 9C B2 84 86 D6 05 A1 CE 6C 09 96 5C E0 CC D2
 56 7E 31 5D 67 E2 15 FE 28 B0 D7 41 20 C1 7A 09
 E5 1A BF 6E E0 73 4E 87 B3 82 A7 26 18 60 1E F6
 40 EB C0 C1 FB E0 03 73 12 60 FD 7F BE 5A D1 79
 E5 45 3D 08 66 45 6B 86 6D 34 8D 65 00 8E C1 A1
 4D 24 BC 55 13 81 3C 81 CF B2 F2 9E 16 01 C1 2A
 64 79 08 ED 10 B8 21 BC 05 6F C4 00 87 E5 76 7A
 6A 02 DA 11 A1 39 FE E4 AF 10 26 11 91 4E 71 27
 1D 42 F1 92 77 8F 35 D7 2E 66 D8 5B 24 C4 83 2D
 EB 66 C5 E4 AF AE ED 51 57 EA 9D D0 D9 91 56 3D
 83 50 D4 5D AD 4B 2A D1 29 C7 32 9E 9F EE 62 23
 1A A4 B6 22 36 3D 54 7C E0 64 20 4A 73 ED 19 65
 5A 1C 5C 64 94 72 E8 76 9B 10 44 DF A1 23 9D CE
 B9 70 D7 CF 90 F6 BE BC 9C 8E FB A0 DF FB BF 94
 82 4D 80 85 87 D0 CF C5 8B 89 C8 C4 2D 35 58 0F
 17 E5 B1 CE 48 77 55 49 B5 4A 4D 5C C3 B3 59 D6
 24 DF 76 D5 49 FA 49 31 59 D3 3E 6E 9D 59 D8 71
 8A C8 51 D7 2E D3 60 A2 10 FD 64 3B AE 72 5D 7B
 E7 10 8C 9E E6 1B 07 67 8A 09 19 4A 21 7E F8 9A
 6C B3 92 2F C6 3A 6D 92 3B AF 03 5D 97 8F A5 A9
 3F 67 F1 57 B4 F2 14 33 81 E9 E3 E6 7E 10 27 96
 C6 B0 87 CB 51 7D C3 48 31 DD F4 55 15 31 EB E4
 EC 77 B1 F7 42 2E DA E7 9E DC 45 C4 7A 2A 9E 41
 A6 55 27 93 39 4B 84 9D DF BA 2E 52 B8 04 64 68
 3B 91 AD DC 2B 76 3D 06 48 5A 6A 5D 03 45 A2 4A
 27 D6 50 E5 3E 8C 1E E7 06 0E B6 F0 8E DF 1B F0
 0A 2A 3A C8 C5 D5 1E AF 3C 41 19 E4 1F 9F 45 BD
 AA B6 1A F4 81 AD 9D 9F 50 2A 9B DB B4 D9 80 0B
 79 3B 95 A9 01 68 67 39 44 80 0D C7 A0 1B 4B 14
 A5 6D E9 6E D8 6F 8C C4 B8 14 D8 DB 0A 9A 0F C5
 22 2B E9 88 7E B2 53 F3 43 0C EB 14 47 44 A6 18
 90 69 05 09 7F DE 7C 14 69 1E C8 DE 2C 59 82 3E
 5B B0 0E D6 91 56 EB 7D 4C 0A 30 C8 90 05 FE E8
 EE 2A 6F A7 4B 23 24 1C 79 B9 36 9A 9F 3E 44 BE
 14 D7 84 43 6F 32 AF AE 8E 7F 56 59 4D D2 3E AD
 0E 75 DA E2 F1 47 4A C1 54 49 F7 3D 2C 9B F6 76
 54 D9 FE 2B C8 7E 4B 2A CB 69 D2 1B 1E 9A 43 E2
 23 7B 15 26 BE DC 23 97 44 E0 FB 25 AE 4E A0 67
 20 9E 1F 4C E6 65 A4 56 7D D8 5D 2E 23 09 34 E6
 61 0C 8F 0B 62 04 74 D3 E1 33 2C 8C A6 35 8A 1C
 64 3B 6A 86 6C BD 8A 94 20 B3 2E CA 47 96 A8 00
 61 DC C3 92 93 E0 56 FA 42 5C 6F 8F B0 76 60 0E
 E8 AC BE 61 F6 FE 29 07 B5 A9 B2 8D A7 74 C9 28
 FB 10 E9 9B 9C 61 BB AD 65 04 E0 20 BC 70 F9 43
 8D 6C EB 90 FF EF 46 E1 B4 FD F4 25 71 9C C5 25
 E5 B2 F6 25 FC 87 F2 30 40 9A BC 87 48 AC F8 DB
 DE CB 61 A2 1D F9 F4 26 31 9D 3F 1E C0 E9 A5 84
 B6 43 FF 34 04 29 FA 6F F0 C7 00 73 4B DE AA 67
 65 1B 81 4D E1 F5 C4 14 55 E4 82 A4 10 5E 04 11
 53 6F D5 42 30 96 01 49 D5 2D E9 17 DF 70 3D 24
 5C 27 9D 6A 6E 0F 79 AF 34 05 92 62 0C 0B 6E 3B
 87 57 88 FC B6 46 1B 10 75 B6 B7 78 F1 3C 0C A3
 45 4B 8D AB CC D8 66 C5 1D D0 E0 50 B5 15 CF 2D
 31 1C B8 78 34 35 F4 F7 9E 2B EB E5 4A 7C E3 7E
 92 9F 8A 4F C0 51 CC 45 3C 65 0A 73 D9 A5 62 B0
 9F 94 DE 50 03 F0 49 F7 F4 C2 36 4F B5 3F C2 BB
 72 92 33 33 3A F0 BA 8A 8C 28 4E CE B9 0D 49 FC
 6E 5F 05 AD BD 2C EE C0 25 DB FF 74 CF 5F 20 4E
 CA A8 32 2F 33 CD 6D EC DF 73 1D B3 B2 B3 02 9C
 17 D5 CC 75 CE 5B 45 82 FA 03 8F 1A DD D5 63 94
 24 31 C6 DE 62 E3 AD 39 01 F2 14 BB 36 4B 68 26
 A5 C9 10 EA DC 4F D8 C9 FF BD D3 BF 11 43 0B DE
 D4 D9 55 94 85 DF 14 99 86 19 FB 61 2A DA 0D C6
 68 86 A1 18 07 C6 E9 DB 62 F1 1F FC 75 10 3C 7B
 3C 4C 2D A6 32 84 88 1F 3C 46 CC 5A 95 3B 31 57
 A7 75 98 A4 E0 CC AB 63 04 3C 23 EB 07 46 C4 28
 B8 2A 5D 99 3C 09 09 E0 A9 46 BC 0B 28 22 9E BC
 EA B4 E3 13 8E 12 0D EB 70 93 49 8A 7F 00 76 5D
 62 C2 13 5B 31 38 24 5B 50 09 53 57 2C 0A 65 50
 C3 6F B2 42 D4 FD FC 7F 07 7A C4 45 57 0C 5B AF
 35 42 6E 87 97 48 77 40 A5 75 06 05 6C E9 B4 3E
 66 C2 FC F7 2A 4E 0A 1F A2 C6 AB 70 FE E4 58 DA
 98 91 E4 AB 2E 91 BB 72 C9 FA 84 95 BD 79 C9 F0
 C4 22 50 22 71 05 6F DC 0E 4C DE 42 2C C0 7C A1
 C1 AD 63 00 3D ED 48 DE 4D 4D A1 19 6B 67 E1 27
 30 05 38 D6 14 3D 08 8D B2 0C FD 58 79 5F DB F8
 FE 54 D1 23 15 45 35 91 63 89 72 E0 29 A8 7C F6
 ED CE 7F D6 0E 54 3B AC EE 46 2E 45 C8 A2 0E BD
 A2 67 48 DF 20 F4 6A 27 55 1D 31 37 13 90 8B 09
 B7 D5 47 C5 11 10 5A 94 1C 15 E7 4E EE E4 FF 26
 F4 75 C7 83 AE 8C 1A 50 90 DF 43 6B 70 3D 12 54
 38 81 D9 C3 CA A5 EA 56 57 D3 D8 0D ED FF E8 2A
 43 EE F9 43 3B 73 05 E3 1F 84 72 58 CF 9C 07 CA
 D0 A9 09 B4 5D 7D EA 6B 17 54 9C 36 64 28 48 3E
 6E F7 56 63 CF 5C 06 60 93 19 57 77 2C 74 96 68
 77 0F 89 B6 82 E8 F4 95 0B 4C 52 23 02 F9 AA C0
 6B C6 31 DD 98 82 07 84 29 EC 73 29 61 C1 39 1C
 03 D8 91 5C 0F 64 B1 3D 9A 70 12 24 76 23 95 90
 69 89 2A DD A7 E8 64 EB EF EF 29 A5 48 BE 9F 0A
 27 91 D3 20 3A B0 C4 D5 30 3A 45 C4 70 A1 4C E1
 AE 0A EE ED 8C 70 63 77 82 23 49 4C 0A B1 B2 34
 06 CD D3 03 28 44 FD EE 17 4C 77 B8 80 0F 5E 1E
 9D 88 05 43 7B 10 74 0B 44 07 F6 47 D5 00 78 7C
 71 C5 F3 2F 79 72 58 98 A2 DC 4F 23 BD 75 9C 5E
 D7 2B 20 38 34 17 EC EA 73 2F CD 36 50 C5 DF 62
 AD B4 DC 9E BE 3B 78 8F 60 EE 1A E8 29 7E 3E 9B
 06 CF BD 72 B8 EB F5 9E C4 D1 8A 04 A0 DF EE DA
 91 BC 77 EC 8D 84 DD 18 07 FD 1C D7 64 0C E1 53
 BB 83 04 3A B7 BA 4E D3 5E B4 19 08 CB 93 80 28
 46 A5 70 02 4A 8C 49 27 64 24 B2 FA 0A 75 FF 85
 B2 F8 2E 67 0C 75 B6 27 1E 01 91 BE 96 DA F6 40
 EC E6 BB A7 D9 C1 7D F9 81 9D 98 29 F9 CF 64 84
 E4 F4 8E B5 7E 77 34 FF FB 40 A6 FE E5 21 24 54
 19 07 78 00 02 D2 F3 4A C0 1A 40 A1 66 C2 B5 8A
 0B 1F 12 06 54 82 4B E4 78 03 9D B1 A3 A8 CD B9
 F1 95 72 9B F7 49 62 69 75 84 D0 9C 2C FD 9D B9
 44 18 75 4E 25 80 ED B6 06 8D FB BE 0C 52 EC 8F
 74 C0 B5 25 35 D7 87 6D 3E FB 01 FA A9 2A F9 35
 E2 02 78 CF 99 73 7E 3B ED 6F BF 77 64 38 F1 5A
 14 FD 9B 90 5C B6 31 7D 3E 28 0B B1 56 E9 CB A7
 75 24 00 70 01 25 6E F6 35 80 F5 A8 D5 7D B3 15
 0C 8F 68 2A E7 BD 7F DA AE 99 EE 86 45 9D 9F 33
 B6 96 38 1F 56 75 BF D4 EE 11 AE 85 0F 6E DF CD
 A6 6D DD 88 E7 03 AE E3 0B BC 5A 8C CE 2C A7 4C
 3C 63 5A 06 70 3B B9 90 79 B7 2F AE EC 6B 3C 7A
 31 2A 7F D8 B1 F6 81 46 40 F6 70 D3 FE 9F 18 8F
 F2 E4 BA F2 1B F3 8F CC 34 93 C0 32 1B CB 3D 89
 47 73 D8 71 25 69 A9 1B A8 3A 6A C5 80 58 48 E4
 88 06 F6 A0 11 01 E5 10 90 34 31 12 E7 B3 C9 CE
 16 CB 8B FD A4 61 8B F9 94 6C E0 E6 46 5E F0 B9
 75 C1 BD 89 70 83 C7 8A 72 3C 0C 46 E6 12 25 F3
 D9 F9 31 79 D5 F3 5F AD 64 B3 29 F6 CB A7 F3 5C
 7D 34 88 30 86 07 D7 C4 BA 85 14 28 54 9A 86 DA
 34 59 DB 76 1B 92 A1 13 4C E5 A8 DE B5 5C 32 9C
 58 F3 EE 8A 17 65 D1 AC 5F 6C D2 87 50 9F 34 D4
 75 84 42 B8 4D CA 78 A6 11 90 E7 93 A0 AA EB 8B
 61 BA CE 14 AA 66 90 A6 FC A3 D0 C4 6D 5E EB 94
 09 1E 32 4E 6E 73 8D EA 08 41 58 15 66 60 33 08
 6D 1E 24 29 FA 98 E9 7E FF 51 82 97 3E 3E 90 BE
 7E 85 78 A8 E5 11 D3 14 7F A3 18 47 9C E8 68 13
 97 40 7A 71 9C 7C D0 8B B3 13 DD 20 CB 53 D3 8F
 6D 64 DC 94 D7 36 81 0B 14 83 85 11 81 C9 15 8E
 B0 8B 7B 6B C1 48 A6 CD A7 1F 5C 6D 68 E8 E0 DE
 3C C3 7C E6 9E 9D DE B7 76 20 A3 F4 8D 57 AB DF
 AF 68 D4 F2 32 BE 94 F8 B6 E6 03 6A 0D DE 38 D5
 40 BF F0 93 4C 17 12 78 B1 40 33 1A 21 93 D4 69
 C5 AB F2 D1 BF F7 1D A9 97 58 4C DB 56 B2 11 F9
 86 45 48 CB ED F6 25 58 54 D9 86 0D 5C 2E 2F 32
 BC AE 01 E4 1F D7 0A 41 40 AE 7E 79 4B FA 2A 19
 A6 6C DF 88 DF B3 CB 0A A3 BE DB 29 F3 F0 B4 A6
 BC FB AA C1 B3 28 97 EA 0D 5F 84 C7 69 FC 4B 74
 DF 78 CC 30 24 15 1F 2E 6D B9 F0 54 A9 C0 0B E5
 B0 C0 84 B7 FD 3A E1 CF FC A6 FE 91 A4 6C EF A9
 5F F2 97 00 E7 DA BD DE 48 4E 3A C4 E2 12 2C 61
 82 0C 46 C6 D8 0C F6 EE 13 89 BE E1 B5 38 27 8E
 01 02 A1 63 AF 17 77 49 8B E6 9C AB 39 5D E2 08
 B1 BF 78 6A B2 C4 25 2E 4C 99 3F 9A A2 17 4D CB
 D1 05 82 E0 8D 59 10 13 AE AA 6E AC F0 EC 90 68
 5D 02 E5 EB 24 DE 53 CF 4C 23 8D 30 B1 87 45 11
 E2 8C 89 09 4D 9A 0E 72 C3 13 59 EE 61 20 D4 11
 97 39 14 0F 17 39 32 B4 EC 21 C2 EB DD 44 19 8B
 ED 56 93 74 38 62 36 FD 83 BC 61 BE CC 02 1B 01
 87 62 A2 5C 73 79 1D 36 24 5A 17 4E 18 CD 47 F5
 AB B6 9E A7 F6 43 B6 2F 02 88 CB 49 6D 1C A0 1C
 D1 0F EE 7B 79 5D 56 27 B9 4F 2D 0C C5 89 9F 43
 43 FB AF F8 34 A5 DE 55 A1 06 CD FC 75 67 0A 4E
 7E 7C 4A 9F 72 9E 69 5F A7 49 6B BE 9E E2 B4 C1
 A3 08 50 00 92 33 15 7A 0F 68 4C 4D A5 0B 7B A2
 76 27 40 98 C5 AD C0 B7 21 39 8B BD 01 BC 3A AC
 BF 4A 63 FB 41 3D 25 13 F1 48 10 AE 8D 19 A0 D0
 A8 78 4C 36 8E E7 53 59 4F 1F 38 6D 30 96 DB 1E
 38 84 C2 7B 5D F6 AB 25 4E 7A FE 57 BA D0 1D 48
 5E AA FF F1 0B C0 F7 E2 C3 7D 84 16 0A BE C6 1E
 87 52 97 CA 45 08 D8 B0 AD 27 07 B3 47 D3 0A 7A
 D1 4C 09 CE B4 25 A9 8C B9 69 16 FC 3E 94 93 21
 04 87 8C BD 17 0E CB CD 86 6D 6B 85 57 35 DB 7C
 98 B9 4E 19 69 30 BC 80 90 62 B6 8D AF 9F 87 98
 3B 79 FA BF 08 9D 01 7C CA F5 F0 01 15 32 2B EF
 3E 69 B0 03 8C 49 9D C8 F8 46 49 A4 19 7F B5 24
 4F 7C 9E B7 BE 58 29 8E 12 9D 25 01 2A 71 A3 F3
 10 57 49 8E 3A 50 79 E0 2C D5 75 71 6D B9 CB 3B
 32 79 04 04 D9 61 AE 67 F7 A1 AF 8F 10 67 CC 56
 5F CF AB 11 27 A1 98 9B 4A DF 0D 27 73 B3 9E D7
 D2 29 49 1F C4 83 75 24 5A 70 24 A8 30 B5 B8 52
 AE 53 64 95 D9 B0 82 E4 1B BC E1 B3 C6 E3 93 D3
 67 16 4B 55 C0 56 AF 72 26 DD 7F 0C DB 52 45 65
 E8 D7 7E C2 19 DB 9A 5B 83 DC F3 FD 8B 18 E9 CD
 56 3A FC FB D3 8C 72 6A 89 B8 A3 AB 69 8A A5 61
 1B BF 1D D8 41 D7 5C B4 55 95 D4 F8 A3 2B 09 3F
 77 12 BF 5F 47 52 82 90 67 B6 FF 0C 0D C3 EF 34
 C9 DA 8F F2 24 C4 E2 69 2D 9A BB 1C E3 0C 39 2E
 3B 9C 40 D4 10 08 B2 9C 54 41 49 C9 59 D2 9C 00
 05 2F E2 8F 77 36 35 70 D1 1F 43 42 3D 36 9E 07
 E9 88 53 A1 71 01 7B 25 BF 71 DE F4 D5 D4 51 8D
 4D B9 D5 2A 99 0E 22 05 E6 EA 49 2D 20 83 13 6B
 F3 83 14 82 BE A3 4D 86 C2 AB F9 B0 BB D0 46 1B
 10 24 36 BB C5 73 42 CC 68 FB DD EC 8C D9 7A 8C
 E8 FF 7C 95 AA FF 76 F9 BF 62 D7 B8 2E E0 13 CC
 AF 8A 39 BB E0 D0 82 0A 64 A2 F7 BB A4 EB 52 89
 7B 4D F3 43 20 11 01 ED FA F5 E3 37 4E D1 BA 49
 D6 1C FD 4F 66 65 8B 7B 09 18 DD A3 56 40 D1 E1
 D9 43 D6 C7 EE A3 1C F8 80 F7 26 AD D8 08 A7 1F
 B2 92 82 58 59 8F 98 BF 2B 61 61 67 1B 9F DE C3
 9F 6A 73 F4 DB F1 9C C7 67 7B FF D4 7F EE 4B B3
 AE 22 CA 3D A1 1A 11 B5 9D 31 A7 25 62 E6 44 86
 F6 B0 4A FF 35 45 52 00 E9 DD 37 83 31 46 74 7D
 07 E9 5E F4 5B 8D D0 A9 5D DE 64 7D EF 69 2B EF
 85 0B AA B7 AD 3D 0B 3B 18 5A 04 C3 31 73 8E 9C
 A5 21 57 BC 74 B4 17 82 9B E4 97 21 7C 18 47 9C
 77 FA 43 50 92 20 67 D4 25 C9 39 11 97 19 7D 2F
 01 AB F6 C2 C8 FF 46 1F D3 0E 58 A4 3B 27 DC 8E
 50 24 12 51 C6 04 D4 DF D1 CA 2D BA AC 8A F6 2A
 42 1D 8C 14 EB 33 56 68 54 91 A9 C2 8D A1 1C 72
 6C D3 AD 0D 30 AD 94 56 2A 60 74 0A 2C A7 A8 86
 66 3A 54 27 0C 0B 88 24 47 5D 59 DD 65 8B B0 F7
 C3 21 EB A1 A7 06 BF 03 29 57 DB BA 72 21 5F C4
 BF 11 91 A4 8D 91 13 95 AC C3 12 AC FB B5 DA 31
 2E 12 91 4B C6 47 35 0E 51 00 A7 21 4D 62 4D 51
 C6 62 6B 05 68 64 7F DD EE F9 CA A5 A7 86 DE 0E
 FE 15 56 83 31 C9 84 88 F4 0D 2C D9 88 37 A1 9B
 2A 8F 0E 54 BC 04 90 10 8A C2 51 27 F8 EF 51 5C
 10 1F D8 DC E5 BE 3B 68 32 04 4D 27 B4 04 98 78
 AB E4 F5 86 04 2C 00 DA A3 E7 17 E7 14 45 CD E3
 60 11 BB 2F D0 F1 7B F8 69 BB 18 23 EB C1 58 6C
 4F AE AA 24 40 C3 95 F2 45 C1 59 6A 58 E1 87 A4
 6F 9F 21 2C F3 83 C0 C9 74 68 03 03 F9 1F E7 32
 98 D1 B4 6E 91 CE 7E 78 11 99 88 DF 00 98 E9 A7
 01 A9 A5 AF BA 4F 67 00 FA CC 29 98 F5 AE C9 DB
 2F 5D F7 0C 0C 65 D3 49 1D A3 E7 D3 D5 3A 0D 8E
 38 F7 93 CA 30 21 75 C6 80 C8 FB 2B FF 60 2B A5
 09 9C 55 70 2A 08 CF B2 5D 1A CE 4B 82 14 B0 54
 71 68 4B D9 B8 EE BD 6A 25 04 8E A4 1A 6A FB 8F
 2C FB 2A 59 00 EA 45 10 26 AA 54 E9 58 AE 7F 82
 BE 57 9C EE 21 32 FF CD 7A 8C FD DD AC B3 80 61
 80 5D DE 84 8B 8A 83 DA 01 93 A8 8B 1C 38 29 9C
 B1 F4 8B 52 77 F3 D2 3E 66 BA 7B 28 54 93 7C 9D
 CC 3A B7 CB 6A DD FD AF 21 72 DC 83 5B D4 3E 89
 49 72 2B BB 66 F0 18 A6 62 A6 17 E1 3F BC 13 6D
 96 1C 66 06 09 03 A2 9B 7C F2 F2 64 92 C8 D6 55
 13 93 04 6C 99 73 EB A7 24 B6 6C D4 3B 20 D3 A8
 66 8C 72 14 C8 C9 47 4A B2 35 F5 DB C0 69 87 C4
 4B FE BE B0 F2 AC BE 7D 61 8E 78 12 19 60 F7 8E
 92 B4 D6 6C F7 13 56 07 AD A7 B9 A7 03 25 5C 6F
 EF DE DB F1 CA 37 BC CD 2D 42 4B 51 8D EF E6 ED
 CD 1D E3 EE 2D D1 57 7C DE 7F 68 1F 95 E6 D0 39
 F0 DC 69 CB F5 F8 97 AE 6A 39 EA E3 8D 62 80 17
 28 79 93 70 0F BF 9E DA 98 A6 9E BA 90 F8 BA 73
 0C 5B 02 DE 3B F3 8D 62 4F D6 96 33 44 49 96 A9
 45 3C 51 45 E5 FD B5 10 8D BB A8 73 F7 28 6B 0A
 AD D6 40 8E 8D 2F 4A F4 43 13 DC 5B 1B 80 19 A1
 01 2F 06 53 C2 6C 2D 13 8C 1C 78 96 E1 D2 1D 0F
 11 74 9E 1D 76 EE FE 09 CD 1B 95 DB 98 D9 FE 9C
 8B 14 E0 D0 A1 49 EA E1 E2 79 3E D5 C5 D5 46 F4
 C7 66 47 40 13 1A 3F 8A 5D 8E A4 FB A9 81 C6 17
 94 23 1D AF AE 68 B0 5C FC 20 69 9F 01 37 13 83
 81 38 C1 2A 59 FB D0 43 B1 F3 D9 C6 B6 E1 E3 35
 F6 AB AB 03 6A 2C 9E C7 6B 90 EB BE 6E 02 E5 38
 A1 4A 86 53 4F D6 38 77 71 36 49 2D B4 23 76 4F
 5A B0 44 3D F7 2E FD 59 91 AD B0 EC E5 81 AF 77
 38 AD C1 54 05 3A C9 5B 0E 14 CA 29 AD 9F B8 CC
 AA D4 00 A5 88 C5 B5 10 22 7C 90 2E 82 E0 0C C5
 81 72 1A B6 89 94 76 F9 A0 31 AD 69 63 71 14 B8
 1B 14 43 E5 FA 26 53 72 B9 8E 77 1D 6A 83 DF 35
 26 92 D5 D1 39 5A 51 8C 6E FD 41 AB B7 7B 1E 0E
 84 90 21 B9 D2 3F CD 58 47 CE CF 67 1C 94 30 E5
 21 E6 2A D8 AC 48 0E EA B8 CD FD 94 B2 C3 FD 47
 7A 90 BF C9 29 28 22 98 0D 38 29 AB 66 93 2F FB
 E5 66 59 6C 2D D8 BE 63 A7 50 7C A8 D7 38 35 2A
 23 78 BB 66 B6 06 2D 61 71 69 B8 4D 85 A9 B5 A3
 CF 49 80 4F F6 D5 BB A1 AA B7 5F 84 BC 9C 99 2B
 E1 05 5A A7 4C E2 1A FC 48 E2 93 DE 05 EA A4 AA
 30 E5 30 0A 4C C3 CB 23 83 2E 3D 3E A7 3A E5 7A
 9A D6 65 14 DB 6E 2E BD 8D CA C2 14 5C E9 F8 7F
 D4 0A AE 1D A4 98 E6 E7 CA E7 EF 95 EF 2E 99 1E
 A3 FF 99 09 CC 7B 8E DB C2 6A 82 99 82 66 96 30
 20 F2 47 F9 DA 1C 52 FE 37 52 BE 4D DA 30 E0 08
 6E 96 C8 82 67 CF 6D 55 FA D2 2C F3 DB EA 32 10
 53 0C 17 C0 FF DF 38 97 94 C5 5A 74 ED 14 A7 50
 F1 D3 EF AB 84 8A 14 58 26 45 BD BB EA 10 68 C9
 C2 79 E1 96 AF 50 26 A2 5F 6C CD 9E 17 67 79 98
 69 D2 36 81 26 56 DD 75 91 62 FE 03 28 92 8C F9
 57 27 D3 76 B4 34 6A C5 F3 FD 0E 27 D8 D1 58 86
 5F 40 0C DE BF A5 04 FE 54 77 0E 4F AC 4F E2 50
 50 49 F3 8F 2B 0D D0 A1 1E 39 38 C6 6E 97 D4 07
 A7 15 F7 9A DE BA C8 D8 F1 EA 63 DF EE 06 53 DD
 38 18 A2 18 F3 32 22 62 06 B3 8C 69 CE 34 23 D7
 16 51 43 A5 3E E3 F6 1F 2E 0D CF A0 92 29 A5 E3
 DB 5A F9 95 62 25 50 51 E6 EE 84 B2 D7 47 89 8B
 98 FE EC A6 4F 4B AC 9D 51 25 0B AD B3 BF 92 6A
 49 96 2A 77 9D 9F AC 82 7C 11 43 3B 52 2F 5F 6C
 9E B6 AC 41 41 3B 8E 5D 8E FA 47 AB 66 13 BC E9
 7A 63 37 35 03 2E 74 B2 23 95 C8 DA E7 BB 1A 1A
 63 09 89 AD 5E 76 C6 66 55 B1 DC 09 A8 9F 62 25
 79 3A 78 31 1C DC D5 A1 DE 43 96 BC 68 6E 72 62
 B5 B9 D6 7C 42 9D CF 8D 12 41 CD F1 E3 5A AE 90
 8B 42 10 9A 25 0E 2F F1 C7 53 A0 A2 30 2F 56 5E
 7F 25 F6 C9 45 09 46 F1 3C 3F 6D A9 2E A8 31 A5
 7B C0 D7 EB A2 D8 73 C2 B9 B5 87 BD D5 EF 8C 21
 74 B1 1B AE 25 A1 1F E4 5F 6A 8E 02 CF 26 F3 7D
 85 E0 D2 65 C4 89 1C 14 A1 6B 47 48 58 C3 0B 54
 29 89 4E 00 79 AD 05 6F F5 B9 3C 0E 84 EB AC CA
 BB 7D 67 34 F2 E7 AA FC 12 FD 1B 46 A8 C5 39 FD
 94 45 B0 81 9C C0 E0 81 15 AE 1B 10 C3 41 3F 41
 5A 51 4A D5 38 25 2C 5A 32 B7 C1 EA 02 6A AE DD
 D9 1C 31 61 80 77 1A 8B 4A FF 93 85 03 23 D1 C7
 CD 2A A8 75 6C 3A 13 75 6D 42 93 FC F7 B1 BC EC
 74 19 8F D5 F2 0C D4 87 07 6C 78 1E AA 49 BA E7
 4B B2 39 B6 1C 2C DF 0D 04 D3 8F 88 6D A1 1A 8C
 43 D4 5D 8F 65 39 73 3A 6A 18 70 22 CB B1 3E 26
 3A 5F 6E 0F A0 88 6F 60 96 4C 91 78 AE 31 54 F1
 5B 98 26 3F D7 52 55 C7 28 9B 18 C4 26 CF 5D CB
 57 64 BA 9D 24 39 B3 75 CA C7 72 E6 05 D7 4F A6
 3A 7D 87 B4 6C 66 C0 B2 91 01 64 18 37 A6 D3 C1
 B9 C0 F0 5B 47 40 5D F9 3B EC DF B2 66 87 4C 8A
 E0 3E C2 7F D3 CC 18 5D BF 17 38 7D A0 75 34 2F
 D2 08 BA 2A B5 FD 6A CB D3 D2 C2 0A 3B E4 F2 78
 70 47 C0 3F 8C 9D E9 1E 65 DE 82 C6 10 93 53 CF
 8C 1D 75 0D F2 85 4A 51 5E 8A 9F D0 4E B9 D3 7E
 81 D6 29 B1 CF AC A2 39 63 69 A1 99 2B DE 2D BB
 29 BA D6 F1 E8 D1 EF 4E 35 16 21 7A 9A 6A 75 45
 C5 46 C9 CE E0 CF 46 E0 8A 76 EF 2B B4 AB 86 82
 88 3B D9 EA F7 71 96 64 17 24 28 29 D7 E7 AA 53
 E2 33 90 F1 FC 52 FF D8 F8 92 CF 92 B1 53 23 37
 A7 13 BA E7 60 1A 80 99 17 E1 AE 1A B4 73 48 41
 21 54 C0 81 09 0C 27 EA 9D 4F 5D 70 EB 77 D6 CD
 8F FE CF 7E E3 A8 E2 26 5C 2F 88 15 FF 89 94 0B
 9B AA E4 50 EE C2 1F C5 0B A9 5F D6 E6 E3 0B 47
 E8 B3 C8 B6 43 3C 1D 20 10 CB AF 8B 14 E9 D7 48
 B6 DB 6C 11 A4 27 DC EE 16 B5 D0 C2 C5 F9 5D 2F
 DB B5 8F B1 05 B1 D7 C8 84 C1 6A 44 FF 95 B8 2D
 A2 E3 7B 34 4D 26 97 E9 F4 0F 24 8B 89 1E B6 FC
 C7 2E 89 27 EC 6C B0 19 42 0C 8E FB 03 1D 2B 8B
 3C 8F 14 0E E7 8B FC A1 2E 75 B1 07 6E 00 CB EB
 80 9C 76 AA F6 C0 3B A6 D2 C8 2D 0E 72 90 F2 C6
 02 D8 E6 32 6D D0 F6 C0 51 05 D8 69 88 12 32 F0
 F1 9B 7C B2 DE 97 4E 2B 25 F9 40 0B 5C D3 D9 41
 B6 33 CD C3 ED C3 23 3A 48 3B 8F 99 0B 03 2D 4C
 FC 56 80 38 F3 88 13 DB 66 68 E2 44 81 BD 58 AF
 66 D7 55 F3 51 DD 03 94 69 85 CE E1 99 3E C8 97
 6A CE EC F5 E7 F9 57 1E 8A DC B9 55 82 EE 78 9B
 90 10 21 D1 1D 72 AF 70 C9 17 A0 B4 E5 41 B7 0F
 60 60 74 D1 8A 5F AA 7E 40 C9 C0 E9 B3 9D 02 7F
 AA E1 7A AC 09 91 E7 64 88 7A 8A 00 8A 92 23 0F
 C0 E6 C8 8B 0C CA CF 88 95 51 08 BE CD 21 FF A8
 3E C0 09 FE FD 42 4B C9 70 37 B3 5D 04 41 F8 C7
 8C 73 FC C0 A8 1A A6 8B 82 06 A3 F6 6C 1F 7A 8A
 BF ED 7E 0C F8 3F 9E CD 43 C1 02 37 F4 9D E4 A4
 05 32 EB 10 A8 20 40 DE D7 43 91 C3 F7 34 7F 62
 59 E5 07 6A 50 3C 1D F5 03 C8 14 16 52 FD 47 F8
 E5 3A 9E D1 67 CB 69 93 11 9E 78 DA BB 0C 29 89
 56 3D 28 7B 63 38 90 26 A1 5D 03 69 56 F7 FD CE
 A6 04 74 E2 F3 1D E1 DA 8D 5C B4 A0 91 B2 4E DF
 CE 90 F5 89 07 75 18 2E BB D5 CB FF 12 A2 66 D4
 A4 B9 9B D4 F1 0B AA 13 F6 8E 7A 13 0A 33 11 45
 E0 67 A9 95 BD A3 B0 B2 FB 7F 9F D5 D1 F2 B9 D5
 41 7D F8 39 21 64 B3 60 34 1B 28 1E DC B7 35 67
 49 27 58 55 A5 68 69 44 01 99 33 EA 4A 13 FB AF
 05 B7 D2 FC CD 1F AF 4F EC 44 BB 27 85 BF 57 F2
 64 13 FE F1 52 35 90 E2 E7 0E B3 26 21 97 C8 69
 6B 2F D1 02 D7 07 C7 5E 41 1C E5 42 BA CE 50 D9
 BB F7 72 74 8B 22 C4 D1 14 73 82 E3 7A AB 30 BE
 BC 5C CB E5 DF 90 73 CE F9 FB B7 2C A3 EC 94 C9
 11 49 C6 4E 48 E6 E0 E1 E5 EB 77 0B C2 52 40 63
 56 48 DB E9 F5 C7 3E DF 44 CA 8C 34 D9 72 89 13
 91 84 C5 B2 68 36 D9 92 C5 D5 42 BD 11 9A 79 F3
 98 3B 79 01 41 B6 6A 5A A6 66 C3 E8 9A 57 AA D3
 6A AE 60 3C 20 DD E9 26 9E A3 7D 0B 5B 64 A2 31
 BE 15 FD A9 50 73 72 A6 DF 87 5B 52 9F F7 10 1C
 12 F9 ED 88 F4 82 72 45 5B 24 F8 F2 B5 7B F9 E5
 D7 04 28 D0 DC C0 8E 28 81 42 59 43 63 FF 0E 2E
 A5 57 FA 4B 2A 89 90 E6 03 B1 C0 BC 59 DA A6 BB
 24 12 B1 86 54 32 26 37 2F 58 AB 24 41 77 FB 9C
 0B 24 63 FD E4 DC 17 37 1B 83 29 D2 D4 C6 A3 E0
 AA 37 11 19 85 8C 3D E3 A3 1F BA 5B 83 0A 15 37
 70 52 60 D5 C6 A0 33 0E 07 2D 60 72 47 09 8C 97
 F7 3D 3C 75 E4 A6 05 A5 A2 A1 F5 91 83 EA 6D 99
 A4 4B ED E8 6F 39 3A CC AC 51 B6 A3 41 75 F1 85
 EE 04 71 0D BD 45 EF 6F 28 91 EC 23 5B 04 F1 D6
 E8 52 26 33 69 AB 87 E4 28 D6 2A 63 6E 05 C4 A7
 04 A7 90 55 AA 80 C0 48 6D 8E 9E 2B 3F 5C FE 2F
 E9 4E 36 AD 03 52 B3 72 2B BB DB 7D EB AF B4 AD
 94 FE D6 94 2F 06 60 2A 63 7F 57 3E 8D 96 0F 56
 97 45 C0 86 5D A3 E6 DF BB 32 2F D6 84 06 4C 99
 1B 6D 44 61 3B B4 D3 40 94 46 83 63 44 B0 8E 51
 61 AF 65 8D 28 F5 BC 33 C9 99 A0 0D 1F 0C 93 90
 C8 8C B6 F3 7B 82 44 3F D9 67 18 0F 86 B8 C2 17
 98 68 1F C4 69 23 1D 75 50 DB 54 CD 51 A8 9C E9
 17 4E EF 93 FB 6F A8 46 1D FC 43 0D 69 48 10 41
 02 FD 97 46 DA 9B C7 DD 83 DE 35 E9 B8 8A 62 DE
 2B 6C F4 5E D3 4A D4 AC 36 FB 7D 8B 22 63 FD 40
 B3 A6 82 2F 0D F5 8E 92 DD B8 1D 56 B1 8F 49 D1
 49 DD A0 75 B4 16 1C 32 FF 53 E0 72 28 34 A2 3A
 27 1A 21 C3 7F ED 47 8D E0 12 BE C4 44 61 FB 75
 8A 02 F2 C7 DB 51 48 4B E3 25 B4 F0 DC 45 8D 20
 92 AF D8 FA 2F 57 BD DE 99 00 5B D2 89 FF 30 F6
 19 2C 08 C7 1B D5 09 13 02 41 32 E0 08 21 4D 4B
 6D 63 B5 22 5C AE A8 AC F6 98 54 C1 9F B9 C4 E6
 B1 6B A9 BD 91 52 97 4A 65 07 64 AF 8A EC 9C 58
 30 45 9A 3C 11 F5 1E B4 EA 8C 1C 7B E8 6B 32 E7
 05 EF DB E4 BB 17 4C 50 63 84 88 4C 7D 0E 99 D6
 D2 A7 52 73 F4 29 07 21 CB DB FC 2B 76 6B 06 CC
 9A 6A D3 30 4E AB EC A0 0E 7E 45 35 A2 5C AE 3F
 E9 A0 B9 71 3E 73 59 1E E4 60 42 C0 A0 57 F9 05
 24 0B 7E 4A AB 48 67 5C 02 5B 61 5F F8 D6 65 53
 EE 78 07 67 27 B6 AE 6D B6 F7 77 0D D3 9A 34 08
 03 7E 6C EA 21 BA 8A E4 C1 D0 A5 54 A0 F1 48 EE
 86 33 BB 7C 98 94 2A 53 9C 6B AF 15 57 B1 05 57
 A4 B8 53 7A 60 96 A4 AA 30 E8 47 D0 07 1A C4 E9
 93 2E C9 F0 30 49 65 0C E6 8D 02 1B 19 C6 46 8F
 EA 1B 1C E0 9E FD AF 1E 8D 62 6E 32 62 B4 1C 2D
 7D 85 38 42 AB E7 89 A1 05 84 2C 8F 87 2B 66 35
 EF CC 52 56 68 8B FF 50 3E FB 3E 6D 47 59 9B 6A
 63 39 E3 31 20 7F 47 EC AE 2F 40 73 3B D7 C6 9B
 0D FF 2F A9 54 79 56 22 78 9D C1 70 07 97 C4 3A
 2F EF 8C 02 C0 81 13 B8 83 75 06 E5 4C F1 1C 72
 EE A3 39 B9 CA E1 87 0B B0 F3 D0 AC 2B 3B A7 36
 48 06 69 7A 8B 42 2A A0 70 24 43 E9 CA 5D 50 89
 93 B5 C7 DA BC 97 74 79 1B 9E 6E 12 98 FD 93 13
 74 4B 2F 37 58 9A 23 27 50 00 94 BF 00 DF 8F E5
 D5 B0 4D D5 99 44 D6 DE 73 BB 42 60 CA 3F AA 9E
 B9 53 70 BA E2 69 FC B2 B2 E4 CC 9E E4 9E 8B AA
 BE C7 82 A6 FE E7 EF 08 DA 80 01 8B 47 AC 9F 40
 4B F6 00 AF DE 8E 37 BC B6 88 03 1B D6 C8 8C 02
 BF A9 1E 14 A8 13 43 8C 42 F9 8C 58 35 ED D5 9F
 13 D1 6E 97 A7 59 75 70 3E 6D 7B C0 7F 51 B6 60
 DC 29 BF E2 72 FE 05 C3 CB DE 61 A0 BC C6 5D 6C
 4C F0 32 07 BD 50 95 D7 49 3A F0 93 6D 9A DC 12
 DD 45 26 5D 47 5E 11 74 4E 49 05 42 DC 77 B6 CD
 C8 33 54 52 9F 27 E7 CB 81 5B EE B2 84 E3 3D 4F
 3E 2F 5E DB 6E AC 30 10 F3 3F F0 0A D4 1C A4 CE
 2C 9E F1 78 D2 D2 8E 58 42 BF 71 51 23 74 CE 09
 AA 22 35 FE AE 40 2F 86 75 11 07 5E AB BF 46 BB
 3F 55 FB 5A F2 4E E9 85 88 50 C7 5E FD 3A A3 32
 59 D6 FB 21 47 52 EC 49 17 53 75 7E 07 8F 6F 45
 1C F5 53 03 B8 1F 2D B7 F1 51 22 98 36 36 8C A5
 BC F7 CD 20 2A 84 79 06 82 F1 BB CB B2 6D F2 EA
 A0 48 6C C6 F9 99 BE B6 EF 27 8B 5E A3 43 24 69
 48 32 01 7E F1 5F A8 18 26 3C 3D 5C 70 C2 D4 B9
 5B 30 39 7C ED 7F 9D 06 73 81 C0 81 36 A0 A3 C4
 B1 52 C7 7D BD 57 3E CC 4F 74 FF 87 5F 2D A1 D5
 4E C2 F5 4C FB 02 5B 07 2E 5D E4 BC 73 C5 95 04
 D5 0D AB C0 A1 E0 07 70 B6 10 3F BD AD 20 10 A5
 FD 8C 33 DA 2C B8 94 FA 64 48 E8 96 E9 BA D2 EA
 A2 58 EE AB 9C 2F B4 F2 03 DD BE 72 B8 92 AA 7D
 8B 64 2C DD 89 E3 7E 05 40 77 27 E6 13 CC DE 8B
 69 B0 4E B9 EE 6F DF 3B 47 BB 14 A9 A5 4D 11 45
 8E E4 84 37 8D 7B 20 2F 14 96 5B B9 14 FE 61 A1
 73 38 EC 86 81 2F 78 C8 6F 7D 29 93 DF 93 3F 21
 78 3E 88 E2 A8 55 87 AF 1C 58 33 4C CC CC 42 95
 85 42 3B CB 50 28 48 59 EC EE 70 12 CD 2F FF 40
 FF 45 D6 13 84 CE 5F A1 CF 09 67 9A 83 4C 7A 7A
 28 25 D8 AC B0 66 2D BC E3 58 58 91 52 60 49 50
 77 59 61 4F CE 52 1C 72 07 B9 94 0C 6B 1D 0B 03
 3C 4D 61 85 D1 F3 53 80 AD 3F AA B0 DC F8 BE B2
 52 13 0D FC 01 57 3A 90 44 D9 15 07 16 6F D4 E3
 98 84 8F 74 43 99 23 8C B5 5B 4B 8C 4C 87 7F 12
 B1 CC A4 C2 34 BD AA 37 35 F3 5C C8 A4 07 A9 4D
 74 39 81 08 5F 2E 82 C7 CD 37 B3 FA 3F EE DE 98
 73 F7 02 AD 4E 96 F8 FD E2 79 1D 2C 95 B5 D7 04
 5B B8 14 99 B1 3D 2C 18 DE E4 DB AB E8 45 D0 83
 F6 25 26 C9 5C 3D 5E 3B FA 2F 0F 86 05 54 BF 38
 86 E3 E4 DB 3D 02 A3 95 8A 37 A0 3D FF C7 E4 4E
 CE 60 7D 49 44 B7 9E 17 7B 02 4D 33 44 3E DE CD
 CA FC 89 A2 40 0A D6 59 56 95 A6 55 96 96 93 0C
 5B 9D 9E 6D 31 CB 22 8D E6 EB 5F 7A 3C 61 03 1D
 AD BD 58 CE 87 B2 76 44 3D 68 BE 51 4A 34 F5 11
 6A 8C 34 83 79 74 53 8A 17 5F 51 5A 2B EA 47 AD
 36 96 99 CA A5 04 BA 14 72 F4 FA F6 10 E8 9E 73
 D5 78 15 4D 59 6E F9 14 8F ED 78 FF 61 E4 9B 2E
 4A DF 6A BB 0F D0 C5 D1 9F F9 47 4C 79 B0 51 33
 6E 78 C1 26 C6 59 BE 62 ED BE FC 67 63 4B 2F 9F
 7A 5F F6 0A 6D 85 13 59 EE 99 16 8A 7B E9 2A D4
 22 A7 EB A5 71 62 03 77 49 DE 22 95 39 4F DA 66
 B0 E2 07 E2 93 0D D8 D5 66 FC AC BA 27 3C FA 9E
 30 19 4F D6 58 E3 CB F1 AC 1B 4B E7 A0 D4 F1 20
 47 EE 81 1F 13 A4 B6 A1 71 E9 E2 BB 94 32 51 04
 C5 23 5C 7E 14 DE EE 04 50 11 B8 84 10 C7 5F 94
 78 F2 0B 81 9E 78 08 25 AC 91 0A 96 16 84 00 10
 19 56 16 1A CC 50 FA C1 D3 2F 68 BF 35 95 2A D9
 CF 6E F2 42 2F 11 0C D5 9B FE C7 F4 14 C4 A7 98
 3A E0 20 28 6C 88 99 E0 33 96 5A 55 E5 92 82 5E
 66 8A 12 C8 6A B9 66 30 0B 4C 8C 57 24 19 2A 25
 45 4A 50 71 B7 8D CA 34 F2 A6 80 AB 1D FD 80 3A
 1E A0 F2 2C 38 D0 5C 96 03 51 A2 6C 3D 38 69 A5
 04 14 64 28 E7 50 A1 6B D3 06 D2 96 E8 43 8C A0
 BD E9 B6 50 DD 68 F2 CD 03 12 AD DC E3 F3 A1 83
 CA 27 AB 67 7D B3 F6 CD B1 7C 0E BA 3A BC 3D A4
 A2 14 DC 38 AF E9 2B 8C 44 BB 3D 49 FC B3 2C A7
 DA CB B1 B7 21 BE F1 2E A5 DD 7C DE 37 EB 21 99
 A5 B3 A8 50 DD 88 A4 59 BF C7 33 16 10 3F 43 5A
 03 B7 03 21 28 18 36 C1 A6 DE 42 AE FB 3B 72 E3
 2E D9 AA 38 F9 0E E9 5A 8E 29 08 17 0E 8F 8F 1E
 CA 64 D6 C9 FA DB F0 2D 6F B2 3B DD 60 E0 68 BB
 13 42 9F D0 F0 29 BB 7F CA 88 6E 0C 50 56 A9 E7
 E0 CE B6 8D 3A 82 02 B7 7C 3D 2D FB 73 29 48 36
 50 79 D9 81 FB EC 94 7D 1B F6 34 21 7C 34 03 3D
 0E E1 50 22 C4 CD 50 B8 EB C0 AC EC 47 0A 6A C8
 AF 9C DC 6B BA C9 51 18 27 EF CF 27 E3 F1 9B EB
 B7 C9 0C B6 66 7F CD B9 8E 95 E8 FB E1 6B DC 76
 BB 6B 17 E7 A2 20 73 8F DB 14 3E 92 B4 21 70 86
 05 A0 FA DC 9D 13 FD 33 EA B3 00 52 27 15 5D 75
 E3 BC D8 2D 3F DB A0 69 6C E0 18 B5 E0 51 10 63
 D5 76 7E 77 C8 53 E7 7F B4 B8 83 BD 7C B5 D3 CE
 FD 50 28 C0 53 49 76 D0 63 F8 1A F5 23 FE 4E BE
 43 8F BD D4 42 82 6B C1 C1 2B A9 03 2F 67 1B 5F
 02 A3 93 E3 B6 ED 73 84 5B 7D 49 C8 6D 90 59 C7
 87 02 D7 02 A3 C0 63 A6 25 D3 77 05 C1 05 34 EF
 83 BA 3D 25 96 33 3F E2 47 1A A6 90 EB C2 DF AD
 9E 96 8D 8B 87 AD D0 3B E3 1A C5 17 C0 1B DE FA
 B5 03 43 81 82 9F C2 9A 59 13 A5 43 A6 79 2B 3A
 E4 FB 5F 36 56 67 7B 7B 91 39 A2 00 7D 83 3C 29
 6E 10 9C 5E 3F 97 FC 1B 3E 62 A5 94 65 DB A8 1F
 1A B9 C4 D7 F8 00 B8 6C 77 D1 30 AE 51 9B 30 21
 0A F1 B6 48 39 E0 98 D1 30 4B 17 77 EA F3 92 D6
 9F 70 50 BF EA 67 25 80 57 54 04 5D 0B 19 19 7B
 79 8E 9D 63 B3 16 EB F9 CF 54 D2 55 A5 3E B6 6D
 07 16 D6 51 E2 7C 80 E9 06 68 82 4D 1D FE E0 B8
 DE CA E8 B7 36 AC 5E 05 72 46 73 3B 61 17 66 DE
 FD 32 31 8D 9E CC 3A A4 A1 AE DE FF 4A 6A C7 3B
 9B BC BB AD F6 4C 46 85 21 C6 FE E2 50 6B BE 70
 C8 B0 67 BD 73 22 74 E0 07 C2 21 1B 0E E1 AC E6
 28 3D 48 9E 2A A6 DB 79 FE EE D6 45 D5 5D 9F 81
 21 BC F6 E9 41 05 35 B1 19 89 C4 37 40 B7 93 E6
 AD 5F EF D8 D6 4F C1 35 7F 16 D0 B5 0E 22 F8 1C
 0D 33 37 05 64 C3 A7 EA 14 7A F0 2B 93 5F 45 2D
 58 9B EB 65 34 62 B9 26 D5 A8 56 CC 84 CE A4 6F
 38 5B 11 35 18 88 14 7D 17 B2 3C E8 4B B6 3B 53
 91 FF FA 79 7A F1 E0 BE C2 E7 8E B1 40 2E 90 CE
 5A A9 A1 F5 4F 10 F7 9A 2C B2 C5 3D 0F 4D 76 95
 61 77 DD 74 ED 62 D9 52 B4 19 2A 21 9B 0F FA 81
 1E B6 2B BB 43 35 08 E6 62 22 57 45 18 0F 0F A5
 BA B5 98 41 AC 06 5A 66 50 2D F4 D1 43 33 33 C4
 99 2B A6 D0 DD C3 27 E1 11 C3 FF 0C 55 D5 8A 0D
 08 6A 25 D0 5F D5 A4 B3 D2 49 6E BD 50 42 AA 5E
 7A D6 67 AB 32 9A 9A E4 6E 2F CA D9 96 9D BF 8A
 8A 52 04 C4 D9 36 CD B9 B3 0F 41 B5 02 AE AC 31
 57 36 A4 1B 33 1D 1D 60 ED 5D 5A A7 18 3F 8F CE
 23 BB F8 CF 37 F6 9A 41 D7 FE E0 44 A6 90 A5 29
 35 41 D0 73 1F DF 53 33 69 29 28 6A 58 95 6B 9D
 48 8F EB 7E 5F 1A 82 B2 39 2B 37 FA E3 BD 33 E1
 11 64 AC 72 D1 77 B8 6F F2 A9 02 AC 64 20 7B 82
 3D 95 31 AD 80 E5 C5 52 C3 31 6B AF DD 0A 23 3C
 AC 85 EA E5 8C B1 FA E9 2F FA 6D B3 F4 31 5A 2E
 F2 6C EE BC 3C 9F F4 4A 5C 39 7E 0D 4D 23 9D 69
 C1 B6 6F 35 5D 89 71 CE E4 BE 48 A4 13 FE 61 84
 76 CA 80 F0 06 FB 29 3A B2 0D 91 DF C4 70 59 01
 A7 08 6F A1 46 22 85 9B B8 28 10 EE 05 9D 1A 4D
 41 DE D2 4F F9 79 24 8C D4 CB 12 5B BC E7 A6 FE
 A4 EF 4A 64 4C 4F 9E DD 62 2D 14 B8 D6 EF B1 32
 04 FD AD C8 EE 85 CB 15 B7 A5 01 2A 6C 5E 62 6F
 D6 C4 8C 7D BF F5 B0 43 DB CB B8 0E 7E A8 14 10
 F6 44 D2 49 2D E0 D3 10 37 A9 81 60 DE 06 D1 06
 E9 44 CA A2 F6 8B A6 E4 E4 1F 51 4F 00 E9 25 FD
 25 DC 1C 74 58 CE 79 7A 07 46 04 0B DC B6 8D BB
 6C BF 0F 96 D4 FE 7A 05 52 50 AA C2 DB A0 F5 FE
 44 83 05 DD A8 30 55 82 80 6D 82 8F 83 8C F1 C2
 19 DA 65 6E 9C 29 3F 60 07 77 40 9E 7F F4 79 06
 EF 06 D3 D4 38 84 29 88 91 29 2E C6 4E EB 29 25
 A1 D6 A5 22 DF 18 1E D0 50 2B 2D 16 D5 0D 76 3C
 99 A6 F0 71 B1 A1 82 1E 54 56 2D 99 A0 A7 05 14
 B1 3B 9E B3 8D 9D B5 40 BA E8 D9 FE 61 04 FD 78
 BF 52 B9 A5 2B 05 79 5C 4A 08 9E 1A 3F 3E E7 BD
 44 C6 A1 E7 B4 0F 32 1A 3B 41 40 45 45 4E F6 DE
 7F 7D 8E 24 33 A2 BF 24 DD 90 BE D8 D3 74 1A C9
 EB 0B A7 ED 3F A3 DF 79 67 A4 CB B6 E1 7D 20 F4
 A2 59 EB 6E A9 A1 6E D0 BF 6F 6D 15 0A 5B 4B 3A
 DC CB 3A 33 38 B0 58 69 B2 98 A1 C1 6A 10 30 12
 5F 4E 37 55 BF 05 5C 53 F2 7B CC 35 42 03 95 D1
 15 69 7B D8 5F 13 DE E4 EE 5A 8B E1 F8 72 6C BB
 81 C8 22 D8 89 2D 59 07 69 02 85 CF 66 BA 74 D2
 AF 35 11 C0 21 A5 0D FD 4D 4A D4 2E 4D 42 26 00
 30 94 08 D6 14 DB 2A 35 75 A6 28 7A 0B B7 63 EE
 B7 BF EF 41 30 38 B1 B4 51 85 DF 32 F5 E6 09 12
 7C F5 F6 BE B0 43 A1 E6 CD C2 8F 46 D3 D7 02 59
 65 A9 CC 46 F4 33 74 44 C7 A1 96 F5 D5 0C 9B 16
 BB 9F 31 8E 61 87 24 5B AE 1F 4B 83 0E DE 2E 4F
 28 2E 1A EF 13 77 F8 58 50 D7 1F A3 1A C1 FF 6B
 8B 6D 2C DA AC 26 0F 92 55 2C E7 F3 9E 02 E0 2B
 E5 2C 86 11 58 03 20 39 1D AC 38 4A 7A 6B BD 6C
 7D 03 40 93 09 01 7A 6F 49 86 6B CA 30 E8 52 DC
 2F 82 AE FC 4F 92 F8 13 D4 49 B6 BA 08 F4 8F 99
 25 6D 02 73 60 8F B4 D8 1E 21 4B 19 BA BB 3A 4E
 E8 3E 75 CB C7 A5 9C A8 44 71 0D 6D 4C 7C 9D FF
 EF F2 D2 EF 3E 2C F4 9D DA 0A 2D 8E D3 AA F8 8E
 9B 0D 6A 60 15 B6 C9 24 5A CF 0C 9D BE F3 43 0E
 D5 B9 9E 6C 78 1F 1B 1D 47 EE 2F 02 E1 7E 3C D9
 58 BF 46 40 D5 60 B1 64 30 FF FA 80 07 D1 5C 2A
 7E D0 AD 8F C5 2B 4D A8 AC 14 6E 35 05 48 25 11
 77 1B B1 E4 D1 30 FB 19 DF 58 47 F6 08 96 DC BC
 8F 89 01 AD B7 FF D8 0F 7A 85 52 E0 28 57 83 42
 E1 A9 FF 12 27 C0 79 06 48 0D 93 9B 12 43 25 92
 E0 AF 76 2F 46 D8 E0 B3 77 DA 4E 16 50 7A 18 A8
 C4 7B 41 48 DC AC 5E 70 5D BE 4C B2 29 F4 C9 9C
 61 C3 2D 60 A0 DA D7 9D 43 F1 BE FA 53 62 80 3E
 B3 FF DA 31 09 DA 3A B5 6F 0E 35 C8 5B 24 64 E1
 0F 7B AE 59 CB FC 25 C8 18 CB 06 6C 02 BE 7E 09
 85 97 DC 77 F4 68 36 38 F5 C8 B5 90 A1 B5 FA 99
 8D 0C D9 A5 30 A1 F6 C6 1A 0E 2D BF 46 A0 9C 59
 C5 51 77 A5 9F AF 4A DE F2 67 72 30 79 DF F5 7A
 C5 FE BD 85 B8 8B BB 3C DC CF 23 67 10 2E 9A 3C
 AB BC 67 18 1D 30 8B F9 B7 5E 20 59 0C DB 7F 54
 06 23 D9 46 25 52 E9 09 25 6F 12 94 C5 22 92 CE
 72 4F A4 2A D5 02 CA F4 89 37 DD AA E4 35 C9 8D
 3F 0A 18 51 D2 EB 51 E3 D3 5B E7 9C B0 07 05 80
 44 8A 00 D0 9F 9B 62 FA 63 C6 92 FA 8A 0E 23 92
 E1 DB 16 47 2A 8F B2 4B 22 49 42 BD F6 E0 ED 87
 A4 02 22 D2 6A A2 E6 5A A5 2F 96 0B CC 70 99 5E
 DE 3F 5C 33 6B 57 0D AA B7 BF 9D E4 9E 3F 62 19
 25 6D C3 FC 39 78 F1 85 8D 59 27 A7 91 28 0F B3
 59 D3 EA 30 94 A6 D3 24 4D 2F 07 77 30 2A 74 F0
 12 50 00 FD 81 12 A2 15 37 5E 71 67 DB C4 FC 09
 4F DC D3 D7 57 62 65 00 81 A0 0F 64 3B 63 28 73
 9B 2A 9D C8 FD FF F7 F1 DF 4C 72 80 99 67 DB 1F
 D0 8B E4 3F D5 10 23 CA CD 41 23 34 3A 29 CD 6A
 68 34 DB C3 41 3A EA C6 43 DA E3 1B FC CC 73 D3
 32 FE D1 55 5D B9 1B 2E 81 69 DE A9 D3 85 17 C2
 30 03 61 BA B4 F1 86 3B 48 86 BB 98 76 48 7F E5
 B1 B8 A3 64 34 F7 85 BD 29 1C 56 8D F0 61 82 17
 F9 4F 87 BC 74 80 26 DE 25 F6 45 74 B7 2B 91 3C
 1C 4E 8B 8D 48 68 3E 48 6C 5D CE 04 30 9E 1D 4A
 9A 18 EC 93 0E 09 D5 2F 18 52 3E 3C A3 F4 DE 3C
 F1 0C C0 6E 13 D1 37 AF DA 91 FA 04 AB AD 58 44
 F5 14 49 A8 9A 69 57 0C 9F 07 28 85 D5 9E B3 8F
 FC C6 48 51 5C 7E 7F 16 66 AA 27 7D 72 91 03 E3
 14 6D C1 DB 61 EC B8 93 65 33 C1 C0 C3 9C E2 33
 6C 95 E4 81 1C B6 26 95 EE 68 52 FA 30 23 FE A7
 A8 54 C0 15 DD A8 C3 B1 98 71 FF AA AE 0B 68 D3
 54 1C 13 42 E1 0E 15 69 78 4D 97 2C 8F EF 6D B3
 08 F2 FB 08 21 BF E5 19 01 0D 7E 96 8C D4 65 E7
 01 CD E0 D0 A7 96 0F 7D 12 E1 4C 91 7B 9A A9 3D
 92 50 E1 E6 EA 2F 67 A5 A5 FC 88 D2 AC 59 AA EF
 CA B2 EA 2B A6 67 4B 2C 3A CA E3 ED F6 E8 CA 03
 C6 0C B5 08 4B 00 A0 70 47 2E 85 17 5A CC B1 2F
 0D 1C 13 75 DC 92 C1 79 31 E2 63 0A 8D D1 D4 91
 0B 26 49 CB 2B 2A B7 AD 1A 4B A5 69 F5 D5 03 53
 5B 5D BB 55 BF FE E6 96 D1 F2 C5 07 C0 88 CD A2
 E1 A0 7D 80 A1 CC E0 4C 59 7D C7 AF 5E A5 83 3B
 CF 3C 7D F2 BD BB B1 87 FF 77 DC 09 AA CF D2 EB
 4B 4D 39 A7 47 B8 6B AE 8D 83 CF 1D C6 30 43 D1
 E6 2A B1 B0 C7 9A 04 9E 4F EA 15 C9 C9 88 FB CE
 F4 21 E4 31 3B 65 13 03 0D 87 AF 3E 59 FA 7E DA
 77 77 F1 1A AC 39 C1 E8 DF A7 AB DB 6D DA 24 D7
 DA 68 17 87 DE 03 07 A7 52 F1 75 90 30 D4 9E 65
 8C BB 63 2F D2 FC 5B 04 AF 2D BC E5 18 98 08 A9
 8D 9E 60 78 F3 96 77 FF 06 0A 85 17 80 96 29 54
 5C 76 6F 3E 31 4C D3 E6 4B 58 63 E3 75 BC 5D C5
 DB 83 29 EA AA 77 0C 05 DA F8 A3 09 78 78 BA B8
 83 9E 48 6B 28 0B B3 F6 02 D5 28 8F 7B 50 09 B1
 57 50 CF FB 87 9A 65 20 57 0E 52 80 CC 86 C1 BF
 FB CE F6 7E BC D8 09 AB 4A 1C E8 C7 FF 98 4B 93
 1E 55 BA F1 54 90 AA 8C 6F 30 17 D6 16 06 86 15
 D9 BE 93 F5 A4 1A 17 29 54 EE 5F 71 7D 9E 20 9C
 70 12 AC C3 3D 8B 4C 46 5E 1D BA 90 4D 57 C9 7E
 43 F0 35 8E DE C2 32 53 7D F6 E3 35 F9 F3 1E 7A
 F3 CC 52 0F 28 78 7B FB B8 4B 30 E0 A0 59 A3 06
 A0 87 3A 06 A0 88 D4 4C A9 2D 90 64 6B 21 A7 16
 8E 8E BE 3C 20 7D D3 5C 49 E0 35 D7 AC 79 DA 3D
 61 ED 24 67 0D 34 71 72 8F 42 DE 43 A7 BD 9F 3A
 C3 06 B3 03 1A 8C 17 73 8D 76 E7 F9 AD 60 E9 B5
 64 AD 14 54 6E B6 70 4D 5C BA 86 B8 AD 47 03 78
 8C 31 6F B6 D6 6D C6 3D 6D EA 94 70 EE DA B2 84
 E5 16 5F 18 AD 43 97 2A 44 7D E5 B2 40 0C A5 5C
 50 4E A1 74 55 D9 C0 22 F3 42 0A 2E 31 A8 7B FA
 43 89 3C 8A 83 02 AB 69 9F 62 08 2D F5 FD 14 A1
 4F A1 F3 5D C8 15 F9 B2 69 2D F6 F8 73 04 D1 33
 6A C6 83 10 D7 E4 D9 F2 21 7F BF 29 D0 F0 92 BD
 C9 FB AF 0E 83 D2 40 4D 4C 08 83 74 79 F1 90 DD
 40 D7 20 0B D9 63 A9 F1 AE 10 4B 79 3B 64 2E 8A
 50 D2 E4 C3 A3 CB 7F 91 72 AC 27 B9 41 23 24 8D
 7A CF E4 2A C6 0F 21 24 99 B1 5A 0F 14 CC 8D 00
 B2 32 CA 44 BF 2E B8 73 7B 09 1A D3 CD B8 52 48
 3D E9 44 81 70 81 89 C1 B7 04 0A 0F 1C 8B C8 71
 A9 9A 31 DF 54 8E 03 CD FA A7 E5 32 98 BF 1D F7
 93 36 E7 76 35 48 AE E8 D8 44 A0 38 BE CA 9B 75
 3B 0A 22 4C 8B B5 7C DC 45 D4 76 D2 7E FE E5 37
 BB A6 2F 78 FF 99 24 AF 5A 4C D6 A0 E4 47 81 9D
 AC 13 46 92 60 9C 72 C2 12 CF 69 E1 BC 32 6C 49
 A7 C0 B9 C7 07 AA 6A 54 71 CC F0 0A D4 00 5B 83
 A8 66 C3 76 18 C4 F2 95 3A 80 A4 EE 6D D9 22 14
 12 54 FC 47 94 F3 93 0D 0F EA E4 3D F1 A8 D9 F6
 9F A2 E4 7B 44 58 DF 85 0C 6C C9 8C F5 76 B7 7A
 86 F4 AA F6 AD 59 40 25 65 C3 1F D2 E2 74 BA 69
 09 D9 B0 F9 AF E6 FF C5 0B BA 21 F1 99 41 D6 DE
 1B 10 93 7A B8 4F CD 2E 60 BC FD 39 0F 01 13 C8
 B9 6E E1 DB 08 6A 93 AD 3B 72 95 7C 9F 88 DA 24
 BF 67 DE D0 A1 B4 FF 60 C2 3F 9A 15 62 09 98 36
 AA D8 41 24 8E 3D B8 11 E8 34 A1 35 C4 C7 E2 57
 0A 92 27 DD 08 87 01 6E 36 27 40 0B F8 A9 CF 41
 48 F5 ED 91 AC 34 B6 7C 34 7B 42 05 5F FE 53 89
 CF 2D 08 41 2A 5F EE 69 77 65 F8 DC CA F4 47 C3
 27 7F CC 4A 41 B5 82 EA 62 C3 C4 85 0E A9 B0 2B
 15 96 B8 F7 B0 C2 EF 1C FB 8C FA 99 BC A5 E8 B1
 7A 79 85 F3 91 B3 83 35 9D 55 3C 8C 42 EF DB 17
 40 06 CD 80 16 E1 0E 17 65 8B 85 5D 66 42 B5 89
 62 4C A1 54 BD 1E 11 57 82 E2 5D 12 C3 6B A3 5F
 0E 97 F9 A7 E6 82 E0 15 8F 27 B8 83 F0 26 F4 73
 40 11 CE 7D AA F2 04 3F E2 F8 41 AF 90 E6 1C 00
 DA C8 C3 C4 DF BA E2 22 65 11 B1 9F 5C F3 3D 18
 D5 6B 91 EB F1 BF 91 64 A5 D3 1B C1 15 1A EE 8F
 D7 D6 36 E4 C8 E3 85 DC 48 F3 31 B9 45 74 18 7A
 5C 48 AC 02 33 4B E8 D2 27 67 FE F7 DB 63 37 CF
 C3 09 F9 12 08 0A 85 F9 0A B4 92 2E E3 C9 56 28
 4C 81 77 B6 EA A6 74 24 2A 2E AB 45 3E FC 38 80
 7B 83 A2 A2 E0 E6 18 1D CA 15 F4 A8 BA 04 DE 7A
 FF 1A AF EC 0B 28 44 AC 61 51 F4 C6 B9 59 F7 90
 34 9E 5C 20 BA FB C4 F5 23 C7 25 1D 02 88 C7 92
 18 8C B2 D4 7E 49 3E D8 E9 D6 59 18 E1 85 D2 A5
 F9 7F 5E 76 18 4D BF 3A 9F 19 E1 0A CF 89 B0 56
 06 5B 18 37 B9 C5 F3 BF 73 A8 7D D5 0E B6 E4 9D
 ED 07 32 C3 77 06 93 F3 72 45 18 50 7F C1 8A 47
 83 9C 96 6A 48 0A 8A F5 BD 06 7F 4C BF 3B 1E 60
 40 43 6F E1 14 B0 2C A7 07 C0 3D 18 5E FF 86 2A
 DB E9 A2 97 D0 B8 8A B9 C8 BE 50 1D AA 0C 65 2F
 41 76 64 68 C8 5A F5 4F E9 FD 47 2F 26 FF 29 5E
 43 69 37 8D A6 00 DB 23 41 10 06 5B 77 FC F1 BD
 F7 F6 CE 36 BB 78 3B 6C 96 DC F6 AE 72 D7 63 FE
 28 E4 BF 7B 50 CC 26 D0 48 23 59 BC 3C 15 66 64
 0C 2F D6 7B D6 5C AE D1 F7 01 5C BC F1 82 C8 8A
 08 E9 6A 1F E2 4A F3 6D 0C 1D 92 33 3B C8 4C D0
 A1 94 EB 7F E1 09 1D 34 C0 33 83 B8 03 09 DF 33
 92 45 26 29 53 46 8A 19 BB 33 14 C8 4C 0F AB 65
 8A 32 B6 98 2D 75 A5 D5 1C 70 6B 5D 69 57 D4 A4
 78 58 9D 86 21 D1 BC E3 37 AA BB 7A 95 42 09 E4
 4E E2 6C 71 79 73 12 07 48 52 2A F9 B7 D6 B9 ED
 39 1F B9 A1 A9 30 36 16 02 EE 04 E6 04 99 03 8B
 C5 C8 E8 16 7F 3E 89 82 91 58 B2 F6 4C 0C 22 4B
 D7 40 48 DE 4E 77 41 24 41 F9 53 CE 0D CC 0D 8A
 B1 EA BA 18 5A B7 A1 A5 EC FB 1D 23 65 9E 38 1A
 18 9A 3E 3E 4B 71 82 FC 20 DB 99 4E C7 79 2B C3
 45 E5 64 F2 21 F6 1A 4C 67 2A A7 86 FC AA CE 5C
 EF F5 8F 03 7A 23 49 5B BA 4C AE 96 C5 D8 1F D1
 DD 58 B5 20 76 70 5D 1D E5 C4 03 26 FE ED 92 0C
 D8 AD B6 7E 21 60 F5 DA 16 15 12 56 A2 C9 B8 4F
 26 B8 E3 6D 7C 06 97 D2 8D B5 33 C5 6D 2B 5F 19
 A5 C4 70 D1 0C 50 B3 19 67 10 6A 43 6E FB 02 90
 80 13 B4 78 8C E4 81 9F CD E9 E3 BD 51 63 1C 67
 D5 F9 EA 51 4B EF E9 AC 10 60 26 7E 2D FA DC 34
 A0 C6 E0 79 17 8B FE 37 40 F4 6B 74 96 F2 F4 B9
 0A 7D 87 9D A4 8D AF CD 2D E9 9E DD 69 39 4D 84
 35 88 41 35 00 97 0E 81 70 97 47 E7 85 88 8A 40
 DC 4C FA 14 AC 82 15 0C D0 20 E2 57 21 43 73 12
 BE AA 85 D6 7D C5 92 7D 7D 19 F8 E5 44 25 2D 1C
 DE 17 9E 13 C9 4D BF 2F 8B 84 FD A5 5F DE F7 44
 BB 2D F2 39 12 D5 75 BD 7B D9 E9 5B 29 AB DB 18
 EE 23 E2 CC D1 50 8C E1 62 78 E8 88 6D 55 CF E4
 12 CA 37 5C E3 71 31 11 31 E6 5C AF 05 43 0E 97
 5E 0B 16 B6 2A C1 49 E7 4F 4C 3A 39 1A A9 2D 0D
 36 FA 16 EA 20 FD 1E 5A C2 E3 72 80 C5 E3 1B EC
 06 43 5A 18 EE FF 6B 04 31 1E 0B 02 63 2D 2B 7E
 E9 EA AD 78 50 9A EB 06 3E 09 D4 9C 12 EA 00 9A
 99 BC 75 8E 33 C0 35 53 78 28 58 3D BA 9F 3F 36
 F6 0A DC 65 72 3A F5 3D C8 98 B5 28 1B F0 5D 15
 BB F8 C8 7A F6 FF E5 A0 2A 4F 58 6C 02 B1 38 33
 FE A7 89 A6 72 38 24 41 14 99 1B 25 79 FC 83 61
 95 C2 B1 08 86 91 88 05 28 36 F6 7B D7 E7 BE BF
 46 67 F9 75 B4 9F 9F CC D3 84 99 D6 FB C0 FA C1
 8E 8D 9A 0E 3C 8C FF BE 1B 0B 98 40 75 B5 25 7F
 BB 49 08 F7 53 88 76 B5 24 68 D0 FA 9E F9 C9 5F
 FD D3 BE FC CF 50 7D 61 CB BE E7 4A 33 8C 91 B8
 20 98 5F BE 95 7B 19 13 D2 CA D0 0B E7 D3 5A 91
 F9 E7 FB 5B 18 31 83 94 0A 44 18 88 21 9F 6F DB
 6A 85 00 1C 7B 97 54 EC 74 B5 59 2F DD 63 E2 68
 58 A5 40 1A 0E ED D6 36 83 31 BA 38 CB 67 80 54
 BB DF E2 73 C7 E0 E4 13 4A 86 33 C2 FB 5D 81 23
 A9 62 0A 02 A7 C7 DB D3 60 D4 F5 38 3D 47 BD 3C
 F9 7B 05 1C ED E4 FC FF 32 CB 45 BE 01 63 48 0A
 85 86 2E 97 F3 1B F7 B3 7F F5 61 4B 31 50 9F 10
 45 CD C4 2E F1 45 91 54 60 AD 58 9F B0 CF 93 EF
 D1 A1 28 26 FC E9 91 62 01 18 22 FF DE 9C 6C 77
 19 51 E9 94 97 26 A8 C1 DC 5E 91 34 36 D8 24 4E
 7E B5 15 F1 F3 27 FB 61 DC 05 E8 1A FC 15 F2 13
 0A A4 0D 5C 20 E9 53 9F A6 1E D7 56 F6 BE BA 45
 A4 DA 5A 02 10 B9 91 9A E6 BD 6C FC C2 E7 FD 83
 4C 46 77 74 F0 56 E5 5B D3 00 DB FA 5F D9 4A FB
 75 F9 98 32 B8 69 4B 50 8F 39 79 16 1C 61 5F D2
 FA F1 A9 78 54 BE 56 B5 B1 61 A2 56 AF C6 F4 56
 E8 5C B3 FD 58 7A C9 6D 54 2D 48 DC 6A AC F1 70
 D0 5A 16 2E 41 18 BE 62 CE 51 5A 57 DC E1 D0 EA
 7B C0 41 6B BD EC A2 17 90 0F E4 C9 A2 0C 19 27
 FB 0D C6 F8 20 CF 8B B8 DA F8 31 BC 68 0C 30 6F
 E5 B1 5A F1 2E 3C 7B B2 80 63 20 03 1F 71 EC 7A
 5E 1C D6 16 1E E8 FF 88 1A 5B 74 4C 4D D6 5F C6
 56 62 74 BB D5 F0 A4 B0 6C EF AE 2B 2B 4A D4 03
 64 BC 26 D6 5C 26 DC 04 15 58 CF 2C 8D 8F C4 B1
 D4 4D 7A 44 39 12 A2 6A 2A 34 CC FA 4F A3 10 29
 C8 6C 31 57 87 CF BC B7 05 25 81 7E 74 5E CB F1
 C1 F5 2F 5D CA 74 1C 54 F2 C2 30 97 B5 4D 16 D5
 64 E7 2D E1 07 23 43 A5 2A D2 8F D9 D0 A8 E3 6C
 0C 20 53 B5 E1 E8 7E FE 56 A7 52 B3 91 5B 60 A3
 17 7F 11 D9 88 D8 47 E1 B2 F3 32 0A 57 D8 6A DA
 F6 69 14 BF 62 1F B2 1A A0 B1 8D 5B F3 D8 51 5C
 C2 9C 08 5F 3A 90 95 2F CC A1 3E BD EC C9 56 E7
 25 07 E1 D9 98 76 D1 13 20 58 EE A0 AA B0 96 04
 E3 6D A8 EF 6D 2A 19 F8 50 3F 2E 08 40 A0 59 94
 3D 23 A0 57 6E 2D 14 E2 C3 0D 7E 14 24 AD 81 59
 E1 A9 70 72 E4 1A D8 FA 82 EC DA 93 42 27 10 32
 BE E0 11 EB DC 73 64 B3 B7 46 FA 4C CF F8 7F F1
 AD 2E F1 07 16 94 C3 3B 29 ED C5 48 8C F6 C3 59
 31 94 51 FF CD AB 7E 14 F3 78 BA 84 6A 25 3B AD
 FF A9 98 FC 53 5B 3B 1F ED 74 5C 5D AB 68 52 1C
 47 36 AA 7B B4 6D 02 BE 5C 2C B0 A1 46 09 CF 96
 0D B5 77 25 D6 42 D1 99 1F 79 05 7C B6 99 10 C9
 3C 26 F3 94 B7 F5 6F 27 94 41 CF 49 49 5D FF 2B
 B2 06 2A DC 31 AC 83 D9 86 D3 B9 DB 87 F9 4C 4D
 0C CF 59 FD DB B7 0D F7 CE AD C2 DB 3A 64 1A CF
 61 0C C4 FA 14 68 F4 78 D4 77 DD 85 3E BD EA 6A
 30 46 8F 58 DB D7 9C ED FF 60 95 6F B3 68 C6 FE
 E9 01 2D 3A 35 83 F5 ED C6 6E 26 96 D0 B4 D8 A9
 84 13 3C 02 EB 10 9D 11 B4 21 DC 21 9A BF 18 32
 5F 40 7A E6 0F 1C 50 AA D2 DF AB 9F 3E 87 1A 7B
 58 D3 C2 88 11 F0 EB 18 E9 D0 59 0E E2 F2 62 71
 86 A3 6E 28 F4 61 2D 7F E7 AC FA B6 69 27 A0 59
 26 6F B7 C1 85 1A D4 34 D1 AE 1A 90 A7 CC 47 FB
 36 70 47 C6 E8 74 52 4E 79 D0 EB 98 B0 C7 56 64
 BA 49 BE 9C ED F0 11 71 9D BB 6C 8C B9 B6 3D 70
 9D 59 7E 56 3C BD FA 28 71 4C 02 0B DE 1B 6F 00
 DE F1 DD 77 ED 47 4D F9 AF 24 DD 82 02 A9 7E E0
 9D E7 76 C0 22 38 14 7D ED B3 1F 91 D4 EF 5A 9E
 85 C1 DB 40 51 4D 45 DC 5F E9 6D 98 DC 22 A7 98
 EE A0 76 07 28 1D 49 1C A9 32 4B 60 8E 05 66 52
 39 CD BB FB 32 A7 C7 95 22 CF 77 E6 EB 90 FB 8E
 ED 95 9B 0F 00 AD 50 A6 51 D7 A2 96 A0 0D DA 76
 E7 0F 29 AC B0 AF 26 9C E6 8D 5C C7 5F AD AE ED
 BC E8 16 39 27 E1 8E D5 FD 72 CE E1 35 51 8D DD
 DA 43 4C 1D 88 DE 4C B6 7E 43 79 64 56 CC CA 3F
 68 5C 0B 50 33 37 ED 81 EC 26 4D 3D AA 08 16 04
 B9 29 1A 0B EF 48 2E 6A C6 E8 E2 04 A3 94 D2 D1
 C5 C0 6E 40 0F 09 46 75 43 09 63 0F 11 69 42 F7
 CC CF CA 5A 65 0A 1C 14 58 5A 27 8D 0B 3A FD EC
 18 4D 6D 54 44 4D B1 CA 74 4C C3 DF 2D CE C3 FE
 A6 54 E7 6C F5 0A 9B 36 74 0C F6 96 97 04 27 ED
 99 CC 8D 34 4B E4 ED 3A 4B 92 95 97 03 74 E4 A7
 57 7D 3B A7 79 8C 58 3F AA AA AD 4F 0B 8F D2 05
 2D B2 BC E5 84 A4 C8 3D 54 62 F0 F0 C4 8E ED 64
 74 7D 32 30 77 EA FD FB FD A1 68 76 49 0F 5D 16
 97 A6 D8 E3 AB 35 32 A4 F4 C8 04 CB FE 08 D5 E1
 75 51 1A 2B 8E 48 E2 CD 4C 87 83 B5 4E D2 0E BC
 86 1A 66 CA E7 48 11 FD 6B 4C AB 07 D5 98 EB 62
 53 07 AD 48 4F B4 5A F8 34 52 EE 71 DF 74 A3 C9
 A2 F5 11 81 B6 12 25 5E 01 23 2E 78 23 AC 7A E9
 36 E1 8A E6 30 56 DE FC A9 C9 52 8A 46 53 49 2A
 69 FF D9 10 88 37 A4 BF F6 99 35 EA B0 8C D8 44
 76 3F 87 8B 21 99 6F 05 9C 68 25 FF 30 41 90 6F
 3F 82 6F 42 4C D6 8F 78 D1 AF 00 D8 17 64 9A 08
 65 71 E1 1C A8 F9 90 FD B2 02 7E DE D9 73 E6 D7
 1C EF E2 D4 70 D3 29 80 CB 93 68 A9 A6 03 32 E2
 BF 8C EF D0 B1 0E 9D 53 BA 8B FE 09 AD 6C 11 0E
 B2 18 58 F2 95 98 A3 A4 8F E1 3A 27 C1 B2 08 39
 37 F0 FE EF 2C B1 89 52 18 14 A9 57 87 41 6F 18
 33 A0 C9 4F 2E 10 04 13 82 13 C0 5C 61 E4 CD 3D
 BC 3F 90 7C 5E E2 22 32 C0 A0 11 6F 47 42 8A 3F
 EE 69 59 A7 10 D3 A4 25 AF C9 EE ED 31 D9 B1 15
 91 05 C1 27 FA 67 12 95 A2 96 7C BB E5 E6 DA F1
 19 46 E2 5C E7 BA 43 52 91 BB 2C E9 B9 EB 74 60
 F8 83 05 DE A7 7C 06 BB D2 39 9D 09 48 F9 81 5F
 31 C2 3C CC D1 4F 89 87 7B BA 1D 7D C9 C4 27 CE
 ED 22 A3 4C B5 1B 47 74 4F 4B 26 8C 5A 38 E9 12
 4E 25 D7 EF FE FA E0 FD 01 97 FC D8 39 AF 6E DD
 24 20 32 5B C3 54 C0 20 8F E3 73 91 0B E6 E3 65
 4B B2 8C 2C C6 9D 2F DD DB 25 A3 83 76 7E 66 D6
 9A B8 5D F3 24 F2 43 D4 77 47 3B 97 9D 3A 0A C0
 EA C5 B4 04 43 75 76 43 01 49 93 64 FD 83 C2 40
 25 0B 92 02 95 90 58 61 76 8F 42 24 DC 5E 37 F0
 03 C7 55 CE 4A 37 41 C8 9F AF 68 46 BA BD 83 FF
 72 D7 39 21 25 40 A1 FE 6A B2 B9 D0 FD 28 93 E0
 29 99 50 DE 8D B6 BE 21 C9 A5 4D 99 34 AD B7 48
 F6 DD 7E 9D EE B1 CB CF 7C CB 0B F9 BF 38 53 BD
 A3 A2 55 DC 53 1D 12 BB 8F 29 1A FA 38 27 C5 C6
 7D 89 BE 4D D6 D9 58 59 9D 39 7F 92 93 21 A2 B2
 11 D6 D0 5E C8 DF 32 EC B9 E8 8B 8A 8A 40 A6 D4
 2E 41 B0 0C 11 A3 5D B6 EC 28 B4 C3 BE 4C 1B 99
 56 93 CE 9B E8 F4 2F 03 B3 58 B0 57 F6 86 EC 83
 57 DA 1C EA 2B B3 EC 07 1A F9 30 E6 C3 E5 A0 1C
 D4 11 72 A5 C6 A6 E1 7A CB D4 E4 06 8B 20 0B 69
 90 F8 48 43 F3 8D D8 B4 9C EA 4B EC 7E B0 6E 7F
 72 FB 45 36 CC AE BB 90 1C 08 69 3C 59 E7 CA 25
 8E 1B 0D 46 8B 33 D9 09 D1 02 22 C1 91 2A 6D 58
 29 24 31 CF 8A 19 37 35 1A 1C DD 3C 20 4F D7 4C
 27 35 02 F6 58 51 54 48 D7 D0 11 16 4D 05 A6 BC
 A8 8D 16 17 56 B2 35 28 54 9D D6 B2 34 86 91 72
 48 72 64 FE 55 4E B3 F6 07 D6 8F EB E1 10 9A 22
 C9 4E 1C EF EC C9 3F 59 B5 01 40 E4 06 0A B5 D3
 0D 22 67 87 DC ED C5 3A D5 48 89 8D 03 8B 42 02
 18 D8 2A 71 16 FE EE 56 0F 43 DA 65 E8 6C 53 F6
 E5 72 F3 82 B8 FC 87 6B FB 5C 10 76 CA 0B 76 70
 19 33 17 25 7B 0E 3A CD A5 83 62 84 56 F6 0D BD
 2D 68 B5 AD BE 2A BE 83 12 B2 A2 58 AA 3C CD C2
 9E 78 9F 1A 15 22 CB 3B FA 66 9A 62 E3 E7 5B 6A
 E1 3B C6 82 00 EF CC 90 21 94 64 F1 39 CB 49 F5
 4F 93 00 EB 69 30 55 5B 08 4D C3 D5 AD 11 5F D3
 7F 7D C6 5A E5 BF CA 37 D8 68 6A BF 43 0A F2 60
 31 30 70 2D 20 6E 3F B6 75 2A 52 BC 5B 6F FD 32
 43 C2 76 9F 65 CB 6F 87 5F 22 D7 8A 5E B6 F5 02
 5F B7 D2 53 55 D7 AC 34 E6 AF CB FE A9 8D C9 32
 66 49 D1 18 1D 2A F7 52 57 D7 A7 E4 0A 97 A4 37
 5C 90 EA FF D4 C0 37 2E 47 57 2B 41 57 F1 7B AC
 F8 B6 3B 25 3E EF 2E F9 5E EA 77 CA D8 B1 14 16
 B1 39 34 36 0D 61 2D 2D EE 75 04 73 F9 65 4A 0E
 16 06 FB FD 77 8F D5 9A 03 D1 7F 47 A0 73 FF 56
 17 2E EF 6D C9 4D 09 2E 3D 7C 95 30 81 CC FC DE
 98 99 13 B3 45 BA 29 D3 0A 11 CE 1D 09 72 A9 A0
 F5 C5 58 A4 E4 AB 3F 21 15 8E 1A CF 49 37 60 88
 FF A2 1E CB 5D 0A 5D C1 72 53 E7 11 4E BF 88 1C
 2F 83 22 ED 1D 38 2C 21 DB 4A 61 3C 7E C5 0E 03
 F4 43 F1 CC A1 6E EF 1F 22 EE 45 57 BB 9E 90 51
 86 AB 03 EE C1 79 94 B0 6A B0 05 FB 2E 67 6E 45
 DC D6 40 CA BA 07 18 29 01 8E B5 6A ED CF DF 3F
 EE 1A 0E BC 20 6E 0F 79 C8 95 13 44 6E 84 11 8F
 CA BE 3E E3 85 CA 7A F3 DE 56 1F 97 56 75 0D DB
 D8 4F C1 90 88 A2 8F AA BB 34 E0 F8 D1 54 AC C3
 0D 70 C7 5F 1D F7 7A 54 40 E7 FB A9 ED 37 88 E2
 3B 53 9C A9 75 0A B8 75 4D 9F BD C4 BA 68 B3 51
 25 30 AC 54 34 32 3E 9A 0F 16 DF F9 5D 0B 41 47
 4B 86 1F D0 BB A9 12 06 A8 D8 B3 14 F1 BB 5A F1
 03 B7 F6 67 F1 F5 FF 04 0C CE 75 C6 24 75 EB 5F
 26 C8 C4 B1 99 57 6C C9 C4 74 0F 66 63 D2 C6 E3
 EB 90 1A 63 D2 AC 96 2D 06 D4 74 E4 22 C4 88 CB
 CF 00 C4 C0 97 45 58 71 09 76 0D 95 21 3F 40 8C
 F4 ED 2C FA 57 20 9F D6 5A 6D 76 55 EE E0 35 02
 F0 97 FA 6D D7 0E E0 6A A8 7E 6F FE E3 51 0D 3E
 EF A6 3B 74 25 3E 64 D4 C1 31 F4 2F 0C 9E CE AF
 ED C5 34 70 B1 E5 F5 07 75 8E 60 2A 9D AD 45 DF
 6F 14 6C 0D 46 19 89 0F 43 A6 4B A9 36 A5 45 7C
 3C D9 1C 91 C8 1F 2A 0A E0 EB BF BC 03 FF AD 08
 BC 7F 79 0A 65 5A 54 1E ED 16 F3 9B 6E 1A 76 01
 4F 0D 79 6B 98 D6 00 16 05 81 52 2F B2 40 2B 5A
 C5 E4 53 3F 29 29 4E 57 74 B0 99 76 2A F4 0C D1
 60 6B 44 8A 6C CE DB 56 1A A1 2B 78 B2 A6 E3 02
 97 FA 43 26 CB 91 43 6F 55 EA D0 A3 FF 81 D6 27
 B6 F5 5C C3 5E 5D 50 84 8C 73 72 27 18 76 DA 4B
 0C 3F 2B DD 3A 8F C6 A1 4D C7 D7 15 02 57 B0 44
 17 FE 5E CE 63 50 A7 82 8E A6 31 39 0E C5 E4 A9
 5C 02 52 58 E9 94 D1 2F 2B E3 9A E2 1E CA FC 10
 6B 1F BE 27 1D 85 58 A0 14 69 FA E7 63 A8 9C 7D
 06 CC D9 A0 A6 CB 77 0D D2 44 E8 9C 99 B8 2F A8
 01 DB 5E C2 7D C4 8F 21 DD 26 A0 81 08 7D E2 90
 3B 61 C0 F4 23 8B 31 26 F3 AC 6C A4 75 30 3B 49
 05 10 CA 61 8F FA CE E9 A7 9C 20 1E 1C 8E 00 74
 A3 18 FE EB 58 AC 5F 2D 14 17 0A F1 FF 02 95 FA
 5C C8 2C EF 96 C9 60 63 8B 39 03 DA FA 43 6D 82
 8D 4C 8E 31 3D 16 83 29 82 E7 CB 44 3B 6B 4C C9
 C1 0A EC 9F B5 38 A8 06 B0 40 11 52 0F 54 77 34
 93 49 4D FD 61 81 F6 A5 20 CE 0C 2E 57 8C 09 0E
 E4 4E 01 96 18 D6 09 FE 01 F7 EB D3 05 77 0E F9
 CE EF DE 3B 0B 6D E5 B5 C9 89 7A C9 8D 74 2C 42
 5A ED 76 17 82 63 8B CC E3 D1 20 43 66 49 7D E3
 F8 16 2E 2F 4E 75 C5 02 8F 79 75 2B 29 EA 87 A4
 1A 73 42 D0 7B 95 50 6D 56 BB 3A DF 47 BF F2 4E
 70 60 CD B6 67 19 98 DF B7 EF 9D 38 4C 00 CC A8
 86 6E 58 E5 27 25 13 30 16 31 69 20 97 E8 7C 95
 40 BD 44 E8 33 AD F8 D4 6C 31 32 C2 B3 1D 11 36
 43 32 E2 48 3C F0 46 9B 64 13 90 51 8D 3E 68 07
 ED 86 CC 2C C8 58 6A DD 57 4C D9 30 10 90 42 45
 5E 8F 9A 38 68 41 93 AF D0 75 B9 8E EE C1 A3 FE
 C4 3B D0 9F 8F 71 70 BB AE 73 18 47 96 03 3F 4A
 96 40 26 9B D8 F6 08 DC CB C5 57 07 C3 CC A7 75
 E5 21 E6 7E 5B 35 DC CA B2 66 27 A3 CC 70 45 BF
 8D 4D 60 5F 1B 96 25 7C DE 77 04 64 52 67 43 79
 E5 05 6D 35 AC E3 A4 4E 91 DF 85 E9 B0 DC 95 25
 5D E1 60 33 43 EB 59 3B 81 05 07 3A BB 55 D1 08
 2C 26 64 B4 EB 8A 65 61 A8 B3 38 10 13 A0 50 EE
 F8 BC B3 71 37 9A BF 26 7B D6 24 B8 3D 05 22 C7
 18 C1 13 87 56 5F 99 01 FF 2B 8F B2 11 40 9E B6
 7C 72 8A 3F 61 EA A3 55 9A 5B D8 7E 3C EE D3 BB
 7C 78 9D 6C 3C A0 30 36 2E F6 CC 80 86 16 C5 7E
 71 D9 5A AD 96 49 67 F4 5E A7 5D 7C CA 74 7A 75
 C1 6D 35 AB 9F 53 5E 03 DE 2B 1B A3 F9 EB 05 D7
 D7 CA CD 61 0B 85 2F 93 DF D5 10 0C 20 1A 0C 75
 E5 D4 D2 05 8E 61 0E C0 97 2C 44 98 30 86 A5 69
 D8 1D FB FE 4A BD 28 DA 86 32 7B 72 89 BD 41 4B
 DF 68 09 47 B6 F6 C4 30 63 09 CD D6 F2 FD 55 97
 D3 5F 68 DA C7 7B 92 90 AB 33 E4 D5 AE 78 B8 EB
 F3 32 61 54 98 D5 9A 5E 26 50 AF DA 94 9A A7 4C
 D7 36 76 86 F2 F2 BD F7 AE EB BA 9E DA 9B 8D 3C
 94 0D 09 E5 A9 F3 3C 0A B8 EE 2C 0B EA 05 8B 34
 64 A4 DF A7 67 26 FA 2E BD 0F CE 74 CD F5 0A 81
 6A 3F 4E 68 EE 55 E8 50 62 82 16 85 50 2B CC 32
 F0 36 09 81 57 78 95 00 68 1B A5 40 C0 CD 69 AB
 2A 68 5A 8D 20 70 6B 3C FD F7 B5 E4 F0 C3 FE D7
 4B B9 3A 9F D0 FE 6B CC AB A5 0B 5E E9 EB 55 4A
 85 1A EC 72 95 37 11 ED 19 09 87 C7 31 6D 6F 44
 74 CD A8 33 0E 02 0C DC A3 83 D2 1C DD AB D4 30
 92 F0 04 53 CF 5F E0 FF 6D 40 62 FC 2E BA 39 D2
 4B 90 99 25 5A D7 1F FB 2A 15 99 F9 81 79 61 B5
 F4 CA 7C 2D 19 E1 56 0A 40 39 D3 27 FF EA EC 76
 37 D5 F1 18 6E CC 00 C5 14 74 5A 5B A1 B5 9A 8D
 20 40 C2 00 14 B9 31 99 C2 96 3C 59 D6 B6 28 43
 9B 80 60 E9 F8 C0 39 3B 7B 8B F7 5D 46 79 A0 1E
 D2 B0 94 09 80 F9 E6 39 42 D4 20 52 D5 F4 EE B2
 A1 7B 00 C3 6C 08 B8 EC 21 8A 62 11 AF D6 E0 AB
 19 AE 5E C2 CC 79 B5 B2 E4 6C 79 33 B6 76 19 87
 0E 6D 00 C3 90 99 02 98 04 2E CE B1 55 C8 48 30
 AF F2 73 5B 02 D4 16 48 77 42 B1 5B C6 9A FA 7D
 19 25 AF 48 34 E6 23 E2 4A 9F 00 AA 91 6A 3E E6
 61 7D 1D F7 3A C6 7F 29 68 1C F4 DB FE 45 AD 4E
 8A 0D A0 B2 B6 CE 95 1F 2B B0 73 95 C8 18 A6 71
 0F E5 71 1B B3 B3 77 4E 6B F6 FC E5 2B BF AE F6
 E1 42 14 A9 99 01 68 36 84 24 BE AC 75 D5 4A D5
 8C C5 C3 BC 1C 05 6D 64 62 62 32 09 DF EC 39 48
 21 94 E8 C6 AE 11 A9 79 41 51 15 5B 7B 46 D1 58
 19 E2 5D B4 E6 DA 42 33 E4 8D EC 4F 7D 3D 47 AF
 D0 0C 61 7B E3 A7 32 05 FB 86 51 EE E2 3E 5E E7
 C9 07 9F 1E 7E F3 78 85 46 96 E8 FB C4 F1 55 B1
 43 E1 FC 21 A0 BF 18 9C F5 5A D4 7D 8E 07 48 26
 07 E2 9B E7 BF 5F 25 81 70 14 35 C2 C8 C1 44 74
 B2 3F 26 C4 E4 93 93 F5 23 F1 F9 B3 AA 30 49 6A
 29 DE 5E 2F 68 52 D1 89 D8 4A BB A2 22 8A F0 CE
 B2 F4 D7 87 BB 34 F1 94 7D D2 BD D0 A5 58 2B B5
 72 58 3B 42 BB 5E 8E FB CE BA 73 1B 55 8A 7A 71
 FD BD B1 75 E6 7C 61 F3 3E B2 46 39 9F A9 8A BF
 51 EE F7 B4 E7 C0 F1 09 F5 AF 9B 9C 37 87 29 75
 3F 0C E3 58 DE CD E9 32 1B CF 30 5A 64 77 27 3D
 CC A8 98 61 41 F9 AE F7 8E C2 E7 0D 3D 1D 8A 18
 32 72 C1 30 A9 47 3F AE B5 40 BD C2 D9 7A 9F A9
 58 79 4D 7E 5A 74 A0 B8 D8 33 9E DF 81 03 B3 62
 E4 3E C6 18 8E 0F 71 11 9A D5 63 27 11 24 A0 52
 55 10 73 E3 53 53 32 17 D9 5A 89 50 30 9A FB C5
 04 2D 45 B6 DC 96 BD 33 DD AE 0B BE 88 D5 75 26
 1B 47 B0 B4 F4 91 A7 B2 84 A0 26 03 00 11 6E 9E
 49 A1 A4 19 6F 91 74 EA F2 B3 43 58 B4 D8 61 BB
 FF CC 8D 7C 02 29 7F 02 2F 4F C7 E2 62 08 24 5D
 8C 5A F0 CE 92 87 01 83 16 2F AA 95 49 19 F6 2A
 28 5A B1 41 1E 92 39 42 B9 74 8E 04 CF B4 EF F6
 87 DE 32 DA B3 CA 18 51 AE 4B AF 2B 48 37 A7 EB
 F5 77 C3 DA 92 E5 12 B3 07 79 A4 0C B1 B3 78 57
 CD C0 DA 48 B6 81 E4 49 1F 06 74 A1 ED B9 CB 54
 09 A2 33 61 90 EF 04 89 73 1D 8D 35 EB FD FE 6B
 3C 94 8F 2C A3 4A 9C A7 D8 33 1D 11 5E 92 83 BC
 C2 7C 01 E9 58 3E 2B 97 1B 64 5E C4 70 C0 E7 D3
 C4 CD 5A 8D EA 76 92 45 D0 C8 9F E4 D5 22 6C E1
 64 61 DA 78 0C 4C 55 FB A8 B6 40 40 50 14 FC 6E
 C4 63 3F 49 64 6D 78 07 5A 4D E8 DE AD 0E B0 2F
 DF FA A7 AA 1F DF 13 62 36 75 B5 C2 38 2C 7D A1
 2E 65 72 37 12 2A 9F 4B 50 F5 73 3D A3 74 8D 12
 71 49 3A D0 54 CC 5B E1 3A E5 E8 A3 DF 70 16 58
 DC A2 88 BE 2B E1 BA CD CB 24 C6 81 C3 AA 96 55
 AA 9C 02 38 71 03 60 83 BF E8 71 0A CC AE 63 91
 99 A1 50 D8 6E EF 93 D7 54 C0 5D 1C 64 76 51 EC
 E8 D3 08 EA 75 51 99 34 A5 EE 3D 3E 0A 60 1C 55
 64 37 3B 14 0A A2 B5 75 C7 B3 53 C3 5F 72 15 4B
 E6 1E FB 8C 33 8E 73 D7 2E D4 AD FD CA 33 0D 12
 2C 54 CF 35 8A 92 74 44 DC CF F7 CB 29 6E A8 30
 5C F2 92 9E 8F DE 00 33 1F 21 32 DB E3 3D E4 75
 8C 0C 7E 9C 63 AB 4D 0E 79 41 C3 CE A1 99 C7 85
 6F 37 C7 06 CD A2 6B 79 F5 BC DA F8 34 53 29 91
 35 F4 AE 81 9C 73 1B 76 E5 9B 10 64 9C CF 86 BA
 4D 82 19 FC F7 49 0C 00 43 8A D1 98 C9 B2 A1 E0
 57 DA B5 6A EC F2 82 3F 41 2C 65 E1 19 5A 3F 94
 83 21 A5 22 02 13 DB 07 AF E3 07 AD 2D 54 E2 61
 8A C4 53 82 DB 7F B8 D5 65 01 08 21 7A 6E A2 C2
 6E E9 8E 57 A4 63 79 EE DF A6 F6 D2 E5 C4 FD 22
 6D 78 FD C9 47 E4 27 33 64 E9 A7 7A D7 8B 77 1C
 44 CC 3C 6C FF 43 7B 5B 97 6D BB AC 5B 5B D3 40
 21 FE 70 41 82 7C 77 CE 3E 2A 48 75 7C 3B C3 69
 A6 DA D5 DD 26 19 92 0A B4 9D 5D B9 F0 79 C2 F4
 A5 96 DE AD 7A 21 3B 8B 4F 21 3C 58 7B DE 26 A5
 B0 39 C2 0E 06 48 F7 3F 29 8F C4 C9 67 96 F5 2A
 3D 74 C8 14 31 9E F7 6B 83 DC C1 87 11 3F 20 D8
 68 C8 D2 38 7B C1 D4 D0 2C BE FC 71 2B B3 1E 33
 CC 56 63 8E 4A A8 A1 22 B5 62 38 51 4C 9B DB 61
 4C A1 C1 B9 12 57 15 B0 AC F6 DC FD 8C D4 28 58
 E1 8A 43 48 E8 89 99 5D F2 F1 96 D7 ED E0 67 49
 05 69 D2 73 71 9C B8 DC 7E 9F FB 07 FB AB E1 74
 3C 4F 99 08 37 D4 45 71 EE 65 AB 9E DA E8 76 8B
 8E C2 8F 5C 7E A4 49 5F DD 11 40 6E 00 BC 1F 71
 B6 00 D7 5C 07 DF 01 B0 44 B6 25 80 04 1C 46 B8
 03 41 C9 21 17 12 C8 DE 96 EA CB 33 B3 0D 94 1A
 A9 F4 49 6B 72 9E EA 84 14 30 4F 9E A2 27 E7 D5
 F2 CA 0D 0A 11 4D 0D C9 08 22 80 BD 13 3B 40 B8
 01 DB 15 AE 53 C7 0B A6 BA 40 16 5F 4B A8 EE D9
 95 A3 C0 78 A6 F4 ED 8F 6C 43 03 9C 97 5A 64 C6
 D4 04 73 6A B6 F0 04 74 AB B8 3A BD 21 69 F7 EB
 90 C2 2A 0C D1 9C 0C 5B 79 DB 6F 04 63 F1 0E FE
 42 63 81 F0 E3 AA 40 88 54 4D 5C 69 8F 68 47 98
 E5 2B 37 35 60 98 4C 8E 9C BD FD B2 5C D1 70 7B
 C3 BE C7 D6 FB 9A E8 13 BD 04 A7 DE D1 BF E9 01
 89 F0 18 8B CF AA BC FD E2 9E C1 66 E1 4C 4F 5B
 71 0B 85 86 C9 AC 17 47 78 7B 5B 89 06 36 E7 6E
 54 98 9F 7B 9B 45 3D 17 73 28 2D F2 49 A2 0E A5
 E3 D4 F7 52 87 85 44 0D 15 91 0C D6 72 15 97 74
 BD A8 68 9F C8 87 A6 B5 B2 29 B7 B2 98 D1 4F 06
 59 84 DE CE E4 28 E5 8F 82 7D 05 3C 1B BD 09 3C
 66 49 0E D1 44 9D 6A 72 FF 3F 10 5F F3 C7 C8 B2
 B3 55 31 5C A0 7E 26 5E 4C B5 BB BD C0 59 68 0C
 DE 43 26 1C 56 CC 50 0F 65 9C 84 B4 68 F1 AF 9B
 B9 31 F8 28 E8 E1 1B 2E 6D A1 A7 8B F2 58 94 D0
 7A E0 76 93 8E CB BE 9E 2C 7A B7 06 B3 85 4D 2B
 43 BF EE 35 14 21 06 C3 38 E9 4F AA 92 29 23 84
 FE FF FD 29 60 62 4E 7F 37 FB 7C FD 28 B8 06 08
 73 E7 62 C3 83 68 A6 22 A3 D9 4F 76 A4 19 47 6D
 65 66 CF F1 CC 02 C8 8D 55 14 1F 9C 4D A7 88 34
 EF 19 95 EB 31 59 B5 4B 21 2D BC B6 ED 9E 2F 0A
 8C 2B 4B CC 20 9B 58 65 C9 85 8B 99 10 0F 3A C2
 F1 D9 47 56 87 D3 37 36 09 50 41 7E FB 50 1C 63
 CF F7 BE DC 76 54 48 A7 E9 7F B3 00 57 33 16 3D
 2E 31 A2 49 3D 6A A6 99 7D 1F EC 2E 63 58 80 08
 D3 0D 12 CA BB 03 03 49 51 E4 A1 85 2D 44 FC 8A
 8B 4E 25 66 10 EE 56 2C C6 60 F4 40 96 BE DB B0
 0F B9 46 15 85 25 3E 01 58 6E D6 96 C4 26 48 02
 4B 6A 8B E9 F6 01 65 D8 79 9D 0B 61 DA B1 34 E7
 9B 56 91 E2 E4 1A 98 C2 FE 19 13 F8 AA 7D 01 07
 26 A9 41 7F 63 10 65 18 69 31 38 1E C1 97 34 63
 25 00 88 7E 6E 66 B8 22 74 A6 06 47 50 98 95 27
 5D 69 A8 01 62 BF 6A F4 9D A2 D5 5A E4 94 F1 22
 B0 31 05 2D 46 58 9F A2 90 A5 FB 8B 6E 91 22 12
 E2 61 22 03 A6 09 03 A4 D2 0C 79 6B 07 FB 38 38
 E0 6A AD 40 C6 F3 B2 D4 6E A4 29 E3 53 78 F4 12
 7D 69 86 59 EA AB 95 0E 7F 77 DE 83 C1 8B BF 89
 9D 28 72 8A 29 67 0C 2C 1E 60 FB 38 91 64 9F 8D
 13 AD 90 32 B4 27 CA C0 52 DC 8D BB 0B 9E D0 52
 C7 CE F3 8C A2 20 E9 BB 2F E6 33 3C 04 A8 7E D5
 2D 02 C5 2C 6B 07 51 FD 6F CA 09 65 8B 61 C2 8D
 33 70 E0 91 AB 27 7C C1 CB 70 12 C0 39 A3 74 58
 2F 0F EC A2 13 7F F1 69 6F 0D B8 39 EA 0F B0 A7
 4C 29 EB 3B A8 CC C5 6A 12 D0 62 C6 65 0F C6 91
 77 6D 78 F4 76 F4 42 EC 30 BD 0A EC F9 27 10 B2
 62 27 B9 EF 60 CB 50 0C 33 10 30 24 01 44 AE 8A
 E5 74 33 17 85 4F B4 BC 9F DA 54 20 60 A9 0B FD
 46 47 4B F5 68 AB 03 2A 08 AE A9 77 D6 EF DC E5
 C1 0D 03 EF FE A4 FF FA AF 19 9D 6E 6E 37 E2 8E
 61 20 07 01 F0 1E D8 C3 FB 08 E0 87 6F 2E 33 A8
 E5 B8 3E A1 B0 95 58 99 8B 67 D6 7F 10 5B 21 53
 29 60 A5 07 5C 57 81 FC 40 B6 2F 26 43 A3 2A EE
 D0 26 13 9C EA 75 AB 0F FA 9A BE 9A D3 6F 74 4B
 5A 91 49 07 2C 6F C7 81 38 3A 88 50 EF 4B A1 F8
 63 39 AF 74 9C 55 4C 62 40 C6 56 78 2F A2 3A 67
 6C 94 F2 7E 81 44 F6 8B CB B8 35 BC EC B0 A0 F9
 31 47 51 70 73 3C 6B F7 C6 53 F6 C7 67 C1 45 74
 DC 25 80 18 07 C6 9A F0 53 3A CD 75 02 E1 3F A9
 5D 9F EE DC 34 23 47 F8 C6 D0 DB 11 A4 B9 17 8A
 69 1E 24 D7 AD 3E 8E 07 DC 9D 9D EC 1B F0 2D B6
 B5 16 A3 16 0E C5 E0 90 4B DC 62 E9 61 3E 4C 85
 82 7C D9 6D F7 A6 C1 5A DC 7B 22 DE 70 E4 1B 68
 79 51 81 34 2E 2F 1D 24 82 F2 55 9B E4 43 75 99
 A2 FD 63 33 BF E5 E0 F8 B1 19 50 7F 72 4E 14 67
 9A 64 AB 05 01 C4 8C 20 2D 6B 7C 59 C8 DA 1C 46
 A3 3C D2 FF 1A 3C 3F 72 90 32 0B 2B 67 80 18 1C
 C3 76 E7 FB AF 78 B6 CC 63 54 FE E4 AC 1A 19 0F
 1D 99 B4 A0 00 73 D8 41 87 51 05 EC 2F 49 46 75
 8D 0D 6B 5A 94 2A 0B E5 58 67 09 24 62 45 14 52
 78 82 85 D0 B2 9A EE 35 F9 1E B8 5B D7 53 8C F4
 4F 3A F2 0C 85 7E 58 F9 1F 60 1C B1 01 21 1D 69
 86 DF 7D DE 94 D0 63 E9 63 0F 36 D9 37 69 95 DF
 C6 EA 88 72 B0 EE 31 7D 00 6C 2E E9 2A 2B 73 F8
 A7 9B 15 F2 D1 3B DC FA C4 46 6F F3 12 66 84 0E
 AA 55 E2 3B 02 A6 8C 11 CC E7 67 B8 77 13 C9 13
 CC CB 17 96 33 99 72 39 2E 8B 53 EA 68 98 48 A2
 24 BC 9D BF 5E 4A 52 8E 25 B5 3D CA C5 6D AD 63
 D1 6C B7 95 F7 EB 98 38 DC CA A1 3C 23 56 C5 4F
 B7 3A 79 37 63 5E 7A 8F FD C8 ED F9 F6 28 3A F7
 BB DE 1F 05 D9 5F 24 9F 57 EF FB 5B 54 3F F5 43
 07 41 F9 AE 57 BA 2D C8 58 17 D7 D3 E4 DA A8 BB
 56 08 9F 84 B3 CC E3 F2 C9 D6 AD 70 A5 8E 3A 37
 E7 E2 55 92 D5 A0 CB B0 18 07 F2 E7 F0 EC 65 21
 34 31 B7 6E C4 54 98 A9 E9 80 EC E7 0B EB D6 73
 4E 0A A4 DD 5D D5 71 38 55 8C 75 D2 06 A4 0C 28
 67 DF 0E 43 92 BB BA 2D 7B E0 81 C3 10 55 B1 48
 D0 1E 88 1D 21 FF 87 93 6C A0 CC E9 A0 F1 81 D0
 9A CA 24 2F CE 6D 43 A7 34 70 CA D4 E5 6C 23 21
 23 6A FE 6D 91 34 1E 7A 4F EC E1 B9 A1 E8 63 5F
 DB F8 36 4A A9 53 12 71 E7 52 9B EB 38 78 90 13
 3A D5 6D BC 32 3F 7F A3 F6 54 69 86 72 72 D1 48
 11 B7 90 1D 3E 70 8E 66 26 13 9D 18 81 33 0A 91
 16 C0 C5 26 88 14 1C 75 8D 0F 2E 89 11 70 23 06
 6A 9C F9 08 70 91 AE 6F FA FD 99 0C 81 93 EE C5
 7D FD F2 FD 1D 82 EE 65 FC 5B 2E 81 44 CD A5 01
 BD B0 B1 21 FB EB 88 DB 8C EF 5C 4C 0A 92 75 DF
 B2 E9 4A 32 9F C5 A6 B5 6B AD 92 A2 59 B0 13 F6
 31 D8 12 BF FA C0 8A 1C 0F 93 12 E9 0B 83 0D 34
 9B D6 E0 D9 A6 1A 44 D0 CA C2 19 AA 04 85 88 AD
 1A 19 68 35 E7 B1 BA BD 5C 7D 87 52 8C B7 5A AF
 45 19 D9 E9 19 32 AA 38 66 08 B6 10 19 AD A7 86
 11 AB 8A 9B 9C 4C 50 EB 03 8C C2 D1 47 77 16 09
 AD D5 35 BA B3 21 BD C0 61 4F E1 BE 5B B0 05 F7
 79 02 BF 2A 4C 47 8C 72 E7 6D 0C D7 7A 99 C3 79
 B0 76 8E A3 E1 46 E1 8E 7D 8D DA FD 69 5A 2C 48
 21 8A 2B 44 D5 18 3B 83 0F D6 31 3E D7 78 7E 2D
 08 35 56 C6 E9 B7 65 E8 D2 EF 49 42 46 CA 9A 6C
 B9 46 A4 1F F1 6A CF 03 EC FE DA C9 1A AE B1 D6
 20 DA 6B 7E 9A A5 DE EF F2 AC 73 AC DD 7B 60 65
 3A 0E AD 74 F4 1D 09 8F 79 C4 48 21 F1 97 C2 1D
 84 B3 65 73 45 85 1B 52 E7 30 C3 3E 8A 09 79 3F
 A7 87 96 FB A8 12 2A A0 D5 4D F2 2F 42 1D 2B 44
 62 E8 F1 29 9D 2B 95 BD 28 73 22 2C A1 F7 8D FE
 07 01 5F 1C 85 93 53 E4 FF A4 3B 70 B6 1B B8 00
 C0 79 1B A4 DF 8F A1 D1 11 8E AB 17 74 04 98 B9
 33 D9 59 B2 37 B5 84 D6 97 58 DA D0 F3 1B DE D3
 37 31 7F 86 C1 93 3E 6F CF 90 6B C4 A3 A6 70 94
 59 6E C5 F7 F8 8D 86 45 76 A6 1A 85 37 E4 6B 23
 7D 04 CB 98 20 D9 CB 81 16 82 A1 F9 74 D2 AA 6A
 BF C7 23 ED FF 82 AC B5 CE 6D D4 A4 D0 90 58 3C
 4A EE B9 EF 15 7B F3 2C B8 63 B6 20 4F E7 59 FF
 20 04 0C 5A 54 75 DE 5F 8F F2 08 6E 2D E4 A3 C8
 AA A3 FF F7 94 4F F1 BF 1F DB 6F B3 73 B6 84 8A
 82 EF B5 B0 58 EE F0 C1 64 99 06 85 4F 4B 40 88
 8F 86 9E B2 0F 85 72 81 D7 DE F9 7F A1 EE 53 EE
 AF 8F 64 35 CD BE 23 E4 6A 13 65 29 2E 72 0B 7E
 9E 60 BC F8 1B 9A BB A2 69 85 C3 77 9F 3E 14 A3
 A8 61 9D 2A 42 C8 74 8A 7A A9 E1 C8 52 84 C0 B8
 33 79 17 17 18 82 D6 94 FE B8 5E 72 BE A9 06 40
 DA 57 83 6C AF 86 B5 1F D1 3E 28 3B 4F B3 76 07
 C4 B7 99 CF FB F3 C7 6D 23 83 2C D0 4D 1C 32 34
 62 32 E8 44 E4 2A F7 BB E0 EC 67 9A F0 CF 04 A4
 AD 80 C6 77 C7 6F D3 F6 A6 A9 39 15 1F 4E F9 BC
 76 5F 69 15 28 DD E5 58 CA C3 14 71 75 85 5C 84
 42 2D 9A A7 E8 76 4E D5 5E 0C 5A 8D 93 8E 1C 90
 C3 63 69 6D E4 8A AA 18 81 9C 53 ED 1B 98 C9 87
 BF C7 C0 58 E0 D8 7F 49 9C 59 B8 1C F3 C2 4B 43
 58 E8 54 09 6E 85 DA 26 AC 45 EC 9E 77 73 F6 76
 E9 FD C3 45 A8 0A 66 A4 D5 D2 19 BE 53 1C 05 AF
 EB 1B 28 19 58 1F 4E 0F B5 0B 71 A1 78 3C A0 B5
 7B 61 A2 CF 4E 37 68 07 D2 87 09 2C A7 46 AE A5
 AE 9F 6B AE CE BE D3 E3 12 22 6A E3 86 C5 80 D4
 38 35 86 E5 D6 6C 03 B8 7A A5 9D 52 98 78 6B D9
 47 6F EC 7A 89 7E E0 29 62 24 AA DF 3E 5A 51 9D
 69 89 F7 1F 4A 3C 9C FB 1B 9F 53 AF 93 30 D4 73
 82 E7 4B 31 63 D8 34 A8 45 94 31 0B C7 68 64 0C
 C9 E4 64 C4 15 30 20 7F 82 D5 48 71 2E 67 B1 37
 CB 7A 7A B6 5D DA AD 62 B9 4E DE 9B 5D AB 62 14
 E7 63 D2 A0 B8 38 A0 CD 2F CE 08 B0 7C 7A C5 10
 3E F8 ED 17 9A C9 36 5F C9 33 26 87 23 36 11 7D
 38 E5 6B 59 CE 7D 00 99 A4 CD 3A 77 7A DA 08 45
 5A 28 76 0B 46 2E BF 3A 4D 0B 7D 91 2D 72 01 D8
 03 17 AC E6 5E 6F FC CD BE CE 27 17 F1 1D ED 8B
 CE 1E F1 E0 C0 33 59 B6 E3 FA 11 92 DB 21 94 01
 F3 0E 03 E6 F2 BE 56 31 51 5C D7 46 E0 57 5F 9F
 97 16 B0 3E 37 F3 BC A8 C0 CC B7 91 A9 5B F4 27
 21 8D F1 D6 10 E7 6C 05 67 EC 16 5F 76 17 6D F2
 37 F4 E4 CC CA 4F 53 19 3B F2 BD 60 F3 00 CF FE
 2A D9 9A 6B CA 43 1A E3 9B E9 F4 09 A5 1F C3 0C
 89 EE 9D B6 4C 7F 0A 3F C8 5B C1 65 DF D9 4C 1A
 56 0F 8D CC EB A6 48 45 92 42 C4 7A E9 2D D1 C1
 2F 33 A5 20 CF 10 3B DC 66 C4 8E DE B7 DF 0D 6F
 B5 A0 BE 95 4C 5B 73 0C 93 7B E8 2A 6E B6 BC 25
 D7 80 61 D4 BD 1B 4E 9F 08 40 77 27 59 4A BD 3C
 C5 70 C3 EC 29 0D 1E A3 55 C1 5A E3 BA 3D FC A7
 1B 52 18 4E EA FB 80 E7 47 63 24 AA D9 4E AF 30
 60 12 AF 91 4F E1 A5 39 4E CB D3 13 0B 74 F2 44
 96 95 69 AC 44 B8 33 FC FC E7 4F A0 4B 0F 3B 1E
 B7 C7 1E F2 8B F3 D0 AB E9 89 03 A4 47 56 4B CB
 76 90 4E 5B BC F4 FF A8 5A 4C F6 DD 6E 7F B9 D3
 0C 9E 1C 0D E9 DF 0E 18 C7 51 F9 5F 23 AE BD AB
 B7 FA 31 5A 2B B9 2C 7B 62 35 8D 3C 36 DD 19 12
 ED 6A 93 B7 DF 88 6C CE F3 3F 75 DE EE E7 A8 6F
 57 AD 8E 47 64 D2 0A C1 EC D9 07 87 74 B9 A9 09
 32 99 BA 21 4F 61 C4 6E 36 ED 23 9A 30 58 93 43
 AA 1B DB 2D 80 DB 29 14 71 46 EF F2 D9 09 3E 50
 F1 3E D4 BC BD F0 B5 0E 48 3D 79 F2 30 1B D7 57
 E2 A2 5F 6F 8E 5E B1 22 3A 6F 71 B8 DE 4D DC DC
 55 47 49 2C 53 6B 6E 2E F3 53 FC F0 B4 2B E5 DA
 5F DE C5 64 B1 9D 62 16 EE 4B EC D2 3F 93 9A 01
 F1 C5 21 20 D1 15 27 19 59 5C FB 0B 01 99 A0 F6
 63 DD 97 49 E0 30 C8 86 A0 8F 28 7A E0 D0 E7 BD
 D8 CA 31 87 3D 95 DB 7D DB 0E 78 3B 33 86 EB C8
 5B B6 11 04 B2 FA 47 88 A2 F9 B7 59 13 43 4C 9F
 0E 56 7C 73 D2 A2 EC F5 93 34 CF 6C B3 05 4E 75
 74 C9 36 97 FA A7 BE A7 81 C2 71 16 77 61 00 95
 3F EE 60 A0 4E DD 5E 1A D2 06 82 FF 3F D2 93 FB
 8B 48 03 6F 76 F5 AE 96 02 0F A0 70 37 61 0D 06
 47 00 70 B8 81 7B BC ED 75 64 0B D0 E2 90 68 29
 52 EC 25 02 A7 87 31 C6 4E 97 9C 53 99 D5 79 2C
 78 AB 1F 63 20 A6 A1 F7 35 97 36 7F 4F 4B 46 C4
 C2 69 6F EA BD F0 83 09 B2 A8 51 FA DB 26 B6 FD
 4A BB 66 B8 18 99 26 6A C8 AE A8 BB ED 9F 25 7C
 DD 09 88 C6 1A A1 3B 07 BA 9D 23 69 D0 02 29 45
 FF 04 D7 6A 22 22 6A 7E 6A B6 48 B7 0B F7 38 53
 B6 3A 61 9E 3C 91 67 AA 8C 7E 8C EC 7F 88 E4 71
 A0 24 A4 6F 74 E0 49 CC C4 B6 C7 A2 88 A3 AF F7
 A5 47 61 B9 BA 22 1E C4 3B 6E 7F AA 7C FC 28 D3
 87 FC 53 86 86 14 C0 76 9D 60 DE 00 AD 12 E6 78
 B9 76 49 4A E3 1B 5C DA FD B9 E7 04 5B 4C 72 B6
 3F 5A F6 AB D7 06 E9 3C FB E5 DA 31 12 AB AF 79
 4F BB 16 45 D9 8E 82 51 4F 83 2B B1 12 D2 21 BA
 CB BF 37 C1 F9 E5 84 D7 A8 8D 2E B5 72 3E 16 83
 AF EC D3 22 D1 27 CC 29 08 35 B2 FB 36 98 5B 37
 47 81 F6 CF 20 33 59 81 C3 9E 56 17 C4 2A 9D B3
 60 62 D2 3B A6 1B DC E5 88 60 B1 D7 19 6D 48 35
 F9 EE 6F AF 2D F4 F1 20 18 E6 A1 C2 50 71 B5 B0
 01 87 3D 4E E0 0B 51 A6 03 70 42 6C 42 C2 70 B9
 8C 53 C0 C4 BB 8A B6 47 25 1F F1 09 9C 4B 10 5F
 09 B0 B0 6D 50 1B 75 7E A7 77 A6 E3 E7 AC 50 9D
 BF D3 B0 88 45 F5 5D 48 BF 85 24 5A 16 1C AA 6D
 D3 51 38 AE F3 A2 A7 9A 86 F2 A2 62 D7 9F 3E 36
 AF 26 05 A3 B6 53 75 D6 B7 9D 6C 13 B9 9C 9C 8B
 18 BE B0 29 5C B8 A0 B1 09 B9 CE F0 93 BB 44 40
 9D 7F 6F 35 AF 8B 25 B4 60 03 18 2D 34 55 F8 6F
 A2 3A 62 0B 6C 29 4B 3A FA F1 E3 2C 92 E7 E2 28
 46 7E 36 2C D7 FA 64 C5 8F AB 44 10 00 6D 25 77
 40 74 5A D2 6A 5A 86 BA 02 B4 E1 29 2A 89 89 F2
 89 81 52 0D 98 CB 04 39 CB A6 79 11 E5 CE 68 22
 41 58 16 80 CC 89 48 96 84 73 97 0A 55 92 5C 90
 01 6B B4 65 C6 54 59 9D 28 B8 DF 07 8E 96 16 1A
 D5 7F 9A 5F 73 A1 E5 99 C8 4C 32 C0 43 0F 15 CB
 8A 60 A1 F7 A2 87 30 90 3D 1F 93 7A 17 E8 DA 72
 65 F9 56 7A 30 11 DE 55 53 40 4E 4D B7 3B 24 32
 7C 59 C3 73 D3 D2 C5 F2 80 8A 37 3F 23 19 D9 40
 17 72 F4 DD 57 D2 55 F7 B5 BD 0C BE 54 70 7A BA
 CB AA A4 9C E5 F9 7E A5 DD A2 E8 CC D1 C0 5C 7A
 CB 5C DB 50 1B 0E 0A 73 38 1D DB 40 6A 45 A2 6E
 1E BB D7 36 00 55 3F FB 1D 87 D2 18 D6 C4 60 77
 C7 C9 EF 80 4B 73 8C 73 FB 46 E6 5C 2E 01 69 A3
 A9 04 98 1F 91 79 15 87 9E 1E 91 BC E2 7C 94 33
 6E 1C 2E EA CE 3E 8F D6 17 5E DD F1 09 64 55 3E
 2C 34 11 D1 4B DB 23 F5 AB 2B B7 9E 55 4C 0B 8F
 9A CA 44 AF F8 EC 79 46 B3 67 CB D4 AA 1C 3E DF
 7C 7B BA 70 05 B0 4A D9 37 E6 15 8D 43 5C B2 38
 CD 79 0A 88 F1 23 C5 6C E4 0C 7C D4 F6 89 BA 65
 A8 A4 38 1C 64 EF 77 F4 79 E8 CD BB FF 8C E8 AB
 79 5B 92 C1 C1 C7 80 E0 38 E1 5F EF C9 E0 EB A5
 34 0A 0F E0 04 22 3C 11 3E 10 23 A5 F2 0F 60 70
 D9 C5 63 9A 10 08 69 8F 70 9C AC 51 1C E4 70 A7
 C1 8B 62 84 E2 4C 63 8D 10 0B 27 6D 42 0E E5 76
 FC F5 FA 04 05 76 39 39 BC 38 C4 E4 0E 46 0B 28
 17 D7 38 03 DE A6 1D 21 94 7B 05 9F 30 5F 19 68
 10 06 E8 CF 56 45 2F 2E FE 68 F3 83 BE 0A E7 B4
 E0 92 6E 32 68 F1 03 02 57 18 5D 07 AE 6C E7 A3
 F7 76 1B 52 0E 16 BD 51 02 63 9A AF 0D 41 76 AF
 C8 C2 8B 39 2D 4F F2 F7 F9 DE 5B 7A 97 DC 33 6D
 16 82 D6 22 FD EA E7 6A 1D AA DE 5C 5D 81 D5 14
 5E 16 28 E2 84 72 13 FD 75 7E 8B BE 21 77 3E 04
 57 74 C1 47 B2 F9 8C 47 3C 32 82 7B 6A 67 0B 4E
 47 FD D4 C5 24 2F 12 C0 58 20 10 08 B2 26 04 F7
 4C 00 C6 3F 98 EF E1 35 F4 EC 96 BF 4D E4 1D 02
 D3 45 F4 A9 38 B9 F5 49 02 05 D2 37 A6 76 0B BF
 73 1C E2 80 0C FF 73 43 23 95 48 37 1A D8 1C 31
 F6 DE F0 AD 76 13 A1 7F 48 51 6E 9D 6E 1E D9 7F
 A5 F6 C5 45 3F C0 F0 CD 44 9C CE EF FC 11 75 D0
 47 43 A9 AB 31 AD 28 3C 50 C0 07 E5 1E 82 65 A1
 A0 86 1A 5F 53 07 6B 78 F6 41 FE 54 C3 75 0F CB
 1A 78 84 69 DC 92 7A 96 5B 01 C7 09 7B AD 06 4F
 36 A5 A7 59 69 07 04 AB D4 D7 F8 00 3B F5 C4 8A
 C2 E2 E3 F2 F5 86 D6 FA CA 2D 8D C0 E6 F0 D1 E8
 00 67 03 B4 B4 59 BA FE C4 77 BE 31 95 C5 9C C0
 43 36 90 F8 3D 94 BD 34 20 34 25 1D 40 1A 79 A8
 16 C1 60 3A FB D0 E7 8F E6 ED 26 65 7F 73 DD D1
 DA C0 2B F0 A4 91 79 91 E1 AD 49 E4 7B E5 4B 43
 35 E5 A3 34 E9 0C 1B 69 48 99 34 95 91 39 E9 5C
 56 2A CB 37 AB 31 F6 3E E7 C3 1A A9 0A EF 6D D3
 4E 48 E4 B2 DF 65 61 DE 75 FE B4 F5 85 66 E5 CA
 D7 40 59 7B 44 D3 09 20 03 0E D9 AC 25 B3 90 7E
 BB 00 A0 EC B3 FE FB B8 B5 5F D4 51 FE 43 19 D5
 94 2E 95 CA C1 54 F3 5C A2 6F 6B 12 04 90 47 EB
 C1 6A B6 7C C9 82 02 AB 7E F0 D4 C5 F4 C7 9D 3C
 76 7C 0D D9 3A 5C 82 92 1F 6D 8E 19 40 B2 C5 D0
 5C CF 2D 1D 6C 0C 41 F1 4C F4 CF A9 AB 7F 5A 53
 00 47 34 20 58 A1 2A 69 42 EC AF 02 F2 1F 7E 61
 A9 B5 7C 41 0B 56 09 0E 19 39 0A F7 1F 7B 32 0E
 5E 1B 93 3F 16 6D 42 D1 A2 95 DD 47 E0 96 DA 8F
 9F 2E BB C4 90 EB C1 F3 FC 62 1B A6 79 79 60 25
 11 4C 3C 24 EB 06 5D 7D 91 23 F0 2A 16 4A 23 BD
 42 9B 7D F0 C2 38 4B 50 B4 BB C0 70 1C C9 09 DB
 D3 4C 12 5B F1 91 C3 A0 0D E7 B6 EE 79 68 94 82
 2C EE A1 B5 D9 A0 06 66 91 85 54 95 78 E6 B8 18
 04 6B D4 C2 52 B9 69 7A FD EE 2B 51 6F 49 FD 73
 34 1C 00 A4 1E 11 FA 73 20 D8 F1 25 4A 58 99 8F
 7B F6 27 CC 7B BD CC 93 0D 03 3E 87 67 F7 7C 40
 A5 1A 90 D1 C6 5A C3 24 53 9E F7 AE 3B ED 0E 81
 32 F5 D9 BC 3F BD FF 20 1E 13 DB 3A F3 B0 E6 CB
 B2 AC 37 C8 C7 52 E0 E9 1A 08 60 A3 5D 3A 16 52
 DB 37 93 6C 13 51 63 A6 27 8B FC 1C AB B4 37 10
 4E FF 36 08 D0 D5 57 BC F1 B9 10 D6 48 37 10 49
 A8 30 D3 7A 31 77 36 46 0A 89 B9 6A 69 2C 0A 5B
 9D 05 35 10 81 CC 75 A7 2C 8D 6A 33 39 98 66 F1
 A8 5C 01 ED 24 C5 DC 95 9F 27 77 9C 10 16 20 8B
 69 91 63 AE 68 EF C4 C2 6A EE 8D 18 5B 1B 99 DB
 24 BD 5C C4 11 CB A5 29 95 E0 D0 FF 89 AC DD 0F
 75 8E 1F 6A 59 94 E0 47 D9 29 37 90 6C 3C 3F D6
 17 42 64 46 2D 6F C9 DA AD EC 8E 0E 1A C7 C3 62
 62 6B 3D 87 28 09 C5 F3 F5 0A FF 86 BD D6 E1 76
 CC E0 39 82 01 B7 A5 62 BE 6F 05 C9 83 48 FF F6
 A9 BC E6 E8 1C CE 25 48 48 8B 8C F6 4D B4 5C 23
 0B 57 6B E6 B8 37 51 A5 2B 01 4B 0A D7 D3 8A 5E
 FC B6 6E 0F F9 5E C5 87 C5 54 ED 60 8D 42 5E DA
 5E 28 74 88 74 1B 39 2F F6 CE 0C 4A 2B F8 52 4E
 78 87 A5 DD F4 89 FB 29 9B F3 D1 AB 40 64 A6 7D
 14 44 7C 95 5C 9F BE 0A 17 C7 05 38 AD F8 F1 83
 5B 5B 04 19 4D 6B D8 C1 95 6C 30 01 93 1A 13 E6
 48 FE 26 01 37 25 82 B3 6B CE 8B 5B 9C 83 96 6F
 0A 36 7C AA 19 1A 6E CD 7B AB B2 B5 FD 93 BE 4E
 B6 1C 35 C0 51 4E 3A B2 98 26 0B BD 06 98 95 09
 13 16 55 70 39 E5 0B 56 F0 CA 9F 2C 95 F1 1E C5
 34 49 20 BD FC 77 D4 27 6C BB E0 FF CF 74 29 C2
 8C 41 BA EA EC 28 FC CC 68 F7 7A 5A 43 F3 80 14
 3B 63 60 E2 2A 52 86 05 A2 C0 4A 11 F6 F3 BA 86
 E8 B8 94 E4 95 55 3C 74 79 57 C2 A8 3E D5 0D 3B
 A8 18 21 62 86 DA 04 D5 65 12 AE 78 49 57 81 41
 CA C2 DE 8D 2D 7E 3A DA 00 50 E9 06 E8 CF 07 1A
 ED CD 6E 92 C2 6E FE 93 93 AC D9 CF 3E 45 D0 1C
 E6 D5 1B F3 2E 62 D7 E7 5F E3 DA B3 BB 46 0B 3F
 0F 9F 2E 0C 67 24 60 FC B3 73 F4 39 DE 64 77 2D
 4D 58 06 C0 A7 15 3E 80 6B 78 33 26 6E 42 EC 70
 F0 EA 92 C9 2B BF B3 A6 89 19 82 8D 3D 22 6D 29
 BE C1 22 CB 55 20 EC 50 B8 98 0E F7 0A 4C 45 81
 8E 48 2C DA F9 4B 6E 7A 97 39 33 8F E6 44 64 22
 C6 AD B0 32 1A A0 88 78 8E F3 CF 1C 81 18 53 7D
 89 40 20 2F 7F 49 62 A6 D1 A4 39 E5 3F 34 2E 2E
 72 43 DA 31 57 F9 DD 67 40 7B FC 63 20 F5 14 D9
 E6 C5 FE 78 94 15 E0 AB A0 3A 96 58 92 04 D4 D8
 49 89 EF 16 BF 0B 16 53 BB 48 33 64 FE 0F C3 CC
 E3 10 1E C7 2E E1 66 BA D3 7A 59 CC DD 67 A5 5C
 29 89 BB 11 59 2A CE 37 96 13 1C F4 D6 45 03 CB
 61 6B 8F 4B 06 4F 50 E9 CD AC EC 52 15 29 F8 0A
 14 5B FF 5D 23 69 0F F3 3A 86 F0 19 EE 90 20 03
 18 E2 8A F9 6D 97 FD 93 E5 E5 B3 BF 15 29 59 F0
 E4 CF 85 8E 18 EA 16 F2 85 E3 63 41 FD 09 E6 E4
 82 15 00 F0 54 DC 59 8E 57 12 6C B1 F0 91 10 B1
 FF 21 45 DB E7 8A 2E DB 1A E4 6F 7E 89 BA BB 20
 A8 68 A8 89 E0 23 FC 43 52 B6 CA 41 19 13 45 4F
 7B DA 3F 43 A6 CE 76 60 93 4A E8 50 A6 A0 07 F0
 7B DD 8A 88 7E 2A B4 A6 56 F8 E3 D6 33 75 C9 DC
 73 72 57 13 02 56 56 59 0B 2A BA 33 57 F2 87 3F
 92 22 DE 2E 67 B5 37 B8 7E CB 34 40 4C 22 69 12
 93 E4 AE 4C A2 CA 57 30 F9 CB 38 50 FF 90 12 85
 C7 F8 70 8C 4B 5A AC 15 75 5F 3B 7B 6F 83 83 95
 7F 90 4B C7 93 D0 E5 11 B1 9A 98 9B 14 48 60 CA
 77 9D A6 2C D2 25 56 99 E1 65 0F F5 2A 07 E5 C0
 55 41 19 DE 3A 58 68 0D 33 2A 04 1C 17 2D 7A EA
 AA 0D 6E 0F F8 F5 2B 15 F4 D3 E1 1C 30 28 ED F8
 D2 B0 70 CE F7 55 5A 84 88 15 37 B6 6B 86 0E BC
 8D 3B 83 29 44 A6 83 39 A5 34 7A FD 62 F6 07 E9
 44 B4 0D 68 EE 69 5A 81 5B 73 47 0B 40 9F 64 1F
 19 79 A5 CA 6B F9 A4 6B D1 3A 41 91 50 9E DF A6
 A0 2F 2D 25 66 05 90 89 BE 3A 40 42 FD 1C 14 B9
 40 D4 80 8C 73 44 D9 7B 53 59 1E D9 B6 3C 63 44
 88 FA 0B B5 CC BD 59 AD 7F 52 9E 52 90 A3 81 C0
 4D 37 22 B4 48 C6 1E 45 A4 4A 28 4F F1 09 B0 51
 FE 24 1F 25 98 B7 07 AB 67 3A 3A B2 6E 28 E3 FE
 8C 36 AF CA 8B 96 3A 1A BF AD 52 53 32 3A 0D 4D
 70 8B 7E 34 7D 8F 6A B3 E1 B3 92 CF 28 27 7C 2A
 7C 35 07 62 7C DA 62 D8 1E 98 70 A8 87 29 FD CA
 F0 3D B4 A8 36 4F DD 34 6E 9E 9F 3F A9 AF 65 EC
 25 80 9A B7 13 96 D5 09 BA F8 78 89 E0 62 E6 D9
 E1 16 EE 17 EA F5 78 DE 79 46 29 B3 9A D3 DF D8
 FA 8B C5 5D 94 E5 57 3A AD 62 59 F9 27 61 89 15
 68 E4 53 70 46 A1 9C DB 46 9D 85 A5 9D 5F 14 96
 FC DF FB F3 EE 97 41 84 8E 10 B3 F4 57 24 F7 C3
 46 AA FE 87 92 9D 9C BC 0F 34 67 A5 7B 6F 07 68
 B3 51 B7 14 2F B8 49 33 3D 4A FC C9 7D D2 31 73
 83 49 63 5B 02 A5 D1 C5 37 71 C7 FB C1 BC C2 A0
 9F 74 B9 37 69 70 93 F2 4F DF F5 85 96 29 EF 1C
 51 5A 99 45 E2 0B 7A 65 2B B2 89 70 77 BF F5 94
 86 A1 8C FA B7 FA 77 00 C2 96 DD 29 76 05 51 F3
 31 98 DC F6 EB 00 53 AB 99 68 55 0D 81 E1 0E E1
 D7 8D AE 25 7D E3 B7 24 5C 87 E9 C3 EC A6 AD 71
 86 B2 99 2C 41 5D 93 36 3E 84 45 38 7B 50 44 60
 26 04 F5 65 70 C7 9C 3C 3B FD 50 BA 9E 01 F2 10
 15 C1 78 9B 2D 01 12 83 91 00 68 6F 0C A8 0B 36
 7D 85 73 F5 4D F2 78 95 4A 33 AD 26 1B DA 79 4D
 B9 45 EE 6B 4F BC 04 42 30 51 B1 48 97 8D D8 82
 0B E0 1E 5F FF 68 89 1C 7A 04 97 58 F5 EB B6 2D
 12 36 02 5C E4 97 C8 42 A8 19 F0 34 32 4E 31 15
 0D 83 0B E8 A8 9D 3C 13 4C E2 BE F9 70 71 E2 A9
 CC F3 7A 95 93 DC 76 59 B2 C7 B0 2C D5 59 44 FE
 4A 92 A6 F4 EE 2F 4D C0 DE BC FE 89 B9 F1 88 B1
 7D C0 97 89 61 D4 3D 36 63 18 AA E3 52 FC A9 5F
 66 E2 80 99 43 76 AE E8 F7 71 64 2C EF AB BE 8B
 1C EF 95 A9 5B 45 88 61 13 65 71 13 D0 1E B2 33
 59 1B AB F8 69 9B 7D 2A A6 BF 91 1E 0A 4B FE 9C
 F8 5C ED 95 3D 06 60 60 CB 5D 11 58 23 C6 9D 1F
 A5 FC BE 08 B9 1B 8A 23 95 20 A2 AB A6 2E AF 46
 1F 0E 35 B0 CF F8 A2 50 72 D4 1D E1 EF F4 82 D1
 B5 04 80 B1 45 98 A1 D2 91 38 5D 88 C7 A8 C6 E5
 A1 D8 72 9F AA E1 52 E7 08 17 4E 61 70 C9 D7 4A
 1A 01 AC AE F9 7D EA 3B F1 B0 F2 CF 19 26 D8 12
 FB C5 4F 59 28 A0 7D AE CF 08 50 9C 92 78 77 C3
 B1 D4 A7 7B 9C 49 AC 32 2B C3 D8 FC 81 DA 85 90
 12 A8 B8 6B 4B 54 90 55 13 EF C3 45 D9 A5 EB 2F
 AC 3C F7 B6 D0 F3 92 CE 6C 1D 57 D6 97 19 1A A7
 B8 5C 83 A8 49 A6 46 2F 31 17 3A 6F 53 43 22 BD
 43 E5 1C DB 16 30 28 57 21 64 22 1D CA 2E 82 DA
 2D 2A 18 69 26 4E 9B E5 45 83 AD A7 65 DF 0C 6F
 87 8F 68 5E AA 22 21 6D 1B 09 A1 7D 0A F2 EA 94
 49 79 E0 4C A0 C5 A8 D4 2D A5 A4 3F A2 61 F2 0F
 F5 A7 4A D7 04 7A CC E2 A3 90 C1 02 6C 50 C1 6B
 09 33 32 E7 A7 24 E0 4F 4E A9 7D 14 29 AB 4F 32
 B7 00 75 82 DD 0A 57 D9 48 4B AB 53 EC C5 01 74
 A2 90 54 0B A8 A5 7D 83 6F 20 D4 2A A6 F9 82 9D
 26 EC 44 28 A5 AA 74 C7 A4 17 47 1B 02 6A C2 BD
 F6 B1 F1 4A 85 CB D4 2A 41 25 C3 AE 81 74 06 3A
 0E 7D A3 35 79 23 66 B0 FD 4B 5C FD 17 34 4C D7
 45 CE B9 56 C2 F0 3F 78 59 4A 8C 9F D5 99 91 0B
 E6 5B 4D 06 DD CB 6B 63 87 F7 B5 2E A3 90 39 32
 BE 47 37 1C 88 33 1F 84 18 B8 42 8D FE AB 0C 71
 EC 0C BA D4 31 45 31 AC EE 35 64 30 AA CA AC 6A
 2E CB 3B 86 50 42 6F E0 F1 3C 93 5F 6B 56 E8 31
 34 7B D7 A6 2B 43 AD 7F C6 49 89 7E 1F 5D 00 B2
 E9 78 6E F6 5F C4 93 A8 6E ED EF 20 12 75 67 F4
 2C 50 AA 42 24 ED 23 F2 62 96 7C BB 27 BE 46 45
 20 62 59 C3 DC F2 2D F2 50 D3 0D 2D FD 48 ED 4A
 B2 D5 0C AD 6C 2C 4A 11 FF CF 9A 65 D8 3A D9 26
 53 8D ED FC 72 E9 5A 46 F7 C4 BF AD E1 A9 02 B3
 C8 17 A2 EE F5 48 AB 50 2E 37 52 FF DC A7 6D 67
 E1 19 F1 4B 36 88 98 18 4A 08 FD 94 21 94 53 F2
 B1 8F CE 02 2E 55 96 5D 82 39 DE 2A BF AA 53 44
 D9 D5 FC 97 4D 6B E0 02 F7 EB C6 E7 20 F2 35 A6
 D1 47 66 DC 02 E8 EB 19 7D 95 91 F1 93 CC 98 6F
 30 9E 0C 90 1B 7A 13 F6 CB EB 65 09 E9 07 AB DE
 0B A7 07 03 B5 77 0B 1F 9A 6A 66 D8 F2 26 BB B6
 85 96 F4 11 7C D3 97 7D 45 48 A2 CB A7 05 EF F1
 67 D6 ED 59 4B D7 12 9C C4 2D 61 03 58 75 BC E6
 B3 DE 77 A8 49 1D F7 CC 4C BD 15 79 31 55 AA 9B
 21 08 E8 62 CE F9 FC 86 54 70 14 9F 86 D1 B4 4B
 9E A6 A9 E3 0E 78 0C 30 41 86 93 53 B4 16 C9 FC
 68 D9 9E 5D 32 7D 64 6A 8E 0C 60 BC 02 05 FA 95
 5E E0 3D F4 ED 92 DC 45 E0 AC 12 57 2B F8 F0 90
 9F 67 6E C6 67 74 E4 CA 3E 46 01 B9 65 12 58 83
 92 EC F6 DF FE 77 A7 DB 0B 16 70 73 05 99 77 5C
 E8 0C 39 B4 F2 80 6C F5 76 E4 61 13 66 C2 D0 96
 87 5A DA 4D 2F 2D F4 55 2B 51 77 04 7F BA 02 57
 D3 31 89 D9 C2 A8 72 99 03 8E 37 62 40 37 E3 6A
 47 FA B6 91 F0 D0 EF 3A EF B0 BC FF FC 9D 61 59
 3B C8 C5 BD C4 6A 79 EB 17 07 B1 48 AD 8C 14 99
 BA 7E ED C5 88 F8 5B E0 5B DE 17 48 A3 53 50 46
 05 73 E5 36 88 6B 90 8B 74 DB D7 B8 79 7A A4 39
 31 7E DB BA 20 1F 25 85 DA B5 CA BE 6A 19 CD CE
 F8 B5 0D 7D 95 B5 99 07 67 36 50 7C 28 6E 1C 90
 16 F6 E1 F8 E1 FE 71 52 EE 2B 48 37 83 FB BC 3E
 E3 7B 34 B1 5D 95 B7 83 7D 33 E8 D2 3D C0 26 42
 AD 0D CA 84 F0 F1 28 0A 03 5C B2 62 47 27 63 A4
 D0 81 11 64 90 A0 4F B1 C6 65 F4 EF D9 E4 EE 79
 A7 82 6D 94 80 44 75 B1 89 36 CD D9 5A 46 52 A9
 DE 7B 67 09 96 66 3A A1 FF 00 F7 15 D6 D9 A4 72
 15 D6 D1 46 64 A4 F9 89 CE EA 78 74 27 51 8F 04
 47 D3 C3 7F 0D 3F 05 B5 43 60 08 DA 4C 42 50 80
 40 A3 B6 8D 9F 3C 4A DE ED E8 10 29 A0 2D 0E 17
 F7 82 F9 D4 74 91 D3 32 D5 D8 B9 40 9F 87 7B DC
 95 0E A6 5D A7 05 7E 24 F6 1A BD 8D 1C F4 CE EF
 1F FF 9E EE 42 61 CE 3A 3F 34 83 6D FC 74 EE EE
 22 33 46 B7 4E DD 4D 6F 2F 6F 6F A4 E3 EC 59 79
 AB 59 C0 60 7C 03 DB C4 83 CC F6 AD 9D 06 2C EA
 14 60 02 DA 42 4F 26 76 41 AE 16 A1 E4 BA 0A BA
 5A E2 4B E8 01 4A 2F 0D F0 D3 E5 5D CE BA 41 AB
 8F 51 E5 2A 81 9B 48 53 91 1D 7B 17 43 71 9C AB
 52 D1 4D 22 A5 46 DE 85 BC AD 36 C7 E4 A4 06 F2
 35 42 45 86 99 E3 8E F4 C6 8B A4 E6 48 BA 60 29
 5B C8 11 38 A9 5B 5D A8 F2 8A B9 7B 7F 91 36 88
 F1 6C 5F BB 1D 48 E5 1E 2A 11 E6 E8 0B 17 00 25
 CC 5B B7 D6 46 11 A3 55 B5 51 EA 17 8B B3 CF 41
 C9 80 91 9F AC B1 B2 9C D7 68 7A 5B 67 A9 90 80
 61 AD BB 03 09 29 6B 84 7B 43 35 76 52 38 78 B0
 C9 D2 96 E6 23 03 28 5D 44 EC 63 8E 72 19 C2 0F
 3D B8 DB 56 24 47 64 79 48 47 23 13 3C 64 26 D1
 AF 4B 39 98 4F 5D 27 62 0C 26 90 35 8A 4D 08 A0
 5A CF D7 25 8C D6 CB 9B CB D0 58 70 26 36 80 90
 0E 2F C9 6E B0 49 AE C5 20 CC 40 30 81 D4 B6 F6
 86 47 7B 61 E4 24 D1 BF E2 08 09 DD E0 59 00 2C
 99 14 62 FA B5 5D 1F DB 1D EC 14 DD B5 8B FD 03
 83 67 45 FC F9 98 CF F4 8A BD 95 68 54 DB E1 0A
 17 EA 3B 08 76 AE 89 D0 64 B8 2E CC 5C 7C 59 A7
 BF 18 90 79 CB 10 AE 02 55 2D 1A 5A 09 11 CD 46
 89 EB 62 B9 65 28 30 4A 91 31 AB 92 0B 52 80 45
 BE A4 61 A4 FE EA 13 50 BB B0 E0 1F 40 02 D6 92
 A9 34 B6 49 DD 2F 23 7F 5B B9 E8 7D 34 9A 53 24
 BC 73 08 19 02 B3 FA 67 6D 4A FA 9E 03 4E 75 95
 29 44 D0 61 7C 4C 18 A6 D1 4C D2 30 23 23 4F BB
 7D 4F 6E 02 19 F2 6B A3 DE A4 57 70 7B F2 79 70
 4D B1 22 BC 70 8E D5 87 F2 3A FD AF 18 01 1F 8C
 8A 2B 95 BF E8 7E B4 6C 48 27 D9 2B F2 35 74 17
 0F 4A 0C F7 F3 11 38 E7 BD 81 00 6B BD FA 57 14
 BC B9 92 0D 98 BE B9 E4 A9 6D E1 F0 01 73 F0 64
 C5 7B 6D EF C8 91 0B 79 75 F6 C0 18 D1 DD 84 B5
 A0 C4 8A A0 34 0C 0E 63 69 60 FC BF 1F AF F1 15
 EF F5 B8 48 C7 1E A2 82 32 CC 63 E0 D4 87 F5 B7
 22 D6 3B A2 9B C1 E6 36 46 10 0A D8 52 1D 83 17
 79 6D B7 66 0E E2 02 40 BB A9 56 94 AC AD 81 29
 76 5C F9 C0 BC 71 25 90 FC EA D5 2E 91 8B ED 45
 00 96 4F EC 39 55 15 A3 80 EB 5B 48 16 CD 3C C8
 11 4B 8E 9B 89 39 D5 34 6B 1D C8 70 3A E4 D9 DD
 28 7C FE B4 EE 89 E1 67 D4 09 C5 5C CA 7E 7A 16
 EA 6F DD 7D DF 9B 44 15 95 B0 E2 D7 ED A2 BE E9
 9B 9F 87 9E 3C C5 34 0B FE 39 A1 8A 87 B4 01 DB
 B5 BB F6 B3 68 76 38 92 A6 43 7C F5 E5 C0 7D DB
 D1 CF 8C 24 87 B8 19 80 F4 23 9E 19 EF D4 E4 87
 16 B9 70 A6 3F 7D C4 34 51 AE 8D 3B 76 3B CE EF
 0C D8 CA 44 C4 F7 0F 71 FC A2 91 AE 1C 3C F0 D1
 2F FD 94 FC B2 C8 C2 A7 08 67 9E A7 E1 BE 59 E7
 C8 8E 57 65 72 67 BB 4A 85 AC 47 4C A1 94 59 5A
 C0 D8 9D 9F EE AC 49 94 DC 0F 46 A2 A1 8D EF 0E
 57 17 61 38 45 8E B1 5B A1 5E D1 5A 75 96 21 0F
 FF CA CA 27 71 B5 41 D6 FE 3D A0 84 2B 47 EC 6D
 33 AB B4 7D 5C 3F F7 24 6C 40 59 B3 4F 7E C7 42
 CE B4 5B 11 A1 70 35 6C 9A 86 14 BE A5 B1 E4 68
 87 0A 2C 54 38 34 BA 1B 27 26 3A D3 03 2D F2 C4
 42 91 71 7B BA 78 44 FC 9E 22 3F 62 93 87 09 27
 44 FB AF C0 53 61 8F 57 95 1B F1 A4 2F 18 4B AC
 85 68 AA 61 37 37 8A 0A 3B EE 03 08 AF 24 DA 7E
 47 49 1A 1C 88 31 9C F2 43 12 E5 F2 FA 54 C9 E2
 E1 96 57 C7 6B 8C 26 3F 8A B2 FD 48 07 C7 98 B4
 78 78 AE A0 F4 84 05 51 CA E4 A4 45 80 48 D8 80
 E2 22 66 71 75 06 D8 FD F7 0D CA C2 38 A7 E9 8F
 11 69 4C 03 91 87 EA 54 B2 1F 4D 52 4F A7 7C 6F
 05 1A 06 A3 F5 77 4C F6 E8 B0 E9 05 16 53 0F 51
 23 43 59 99 2C 3D D6 30 5D E5 45 B0 17 67 76 1E
 5E CC EA 3F 20 23 B2 FC 34 7A 05 34 AA 21 4A CA
 56 8A E2 08 27 E9 59 07 4F 02 B4 EB 17 96 DB 2C
 C0 F2 A2 AE 81 D8 66 7F 7F 63 67 10 12 B1 2D 38
 C7 DD 94 37 1F B9 A0 7E C7 E8 58 3E 27 34 FD 10
 86 8E 9B 93 1B AE 73 3E 64 3A 9E E0 95 09 AA 41
 CD 92 2E 13 93 5E A5 AD 84 63 76 99 DC 5B 81 36
 44 62 A3 27 2C 06 73 38 94 78 02 E4 5F 4F 47 88
 96 DF 9F 86 C5 DD 50 BB C7 7B BE 90 94 FD BC 12
 35 BD 90 A9 07 29 BE F6 0B 2D 6E D9 2F 3E 0E 10
 EB EA 1A 70 DE 09 B4 8B 53 72 80 8C 9B 20 A1 29
 2C 72 DE 23 C9 00 88 31 72 96 C7 BD 74 43 A4 C3
 8B D3 AE 07 99 98 2E 90 97 6E C8 8F B0 1D 82 89
 65 1F 57 84 09 1A EF 75 BB 5F 1F C2 09 C8 0E 50
 94 B9 8E 46 B9 F3 75 47 46 BB 7D F2 8C 98 BA 79
 58 B5 E1 89 A7 36 62 7F 08 EA 72 91 EE A6 1A 7B
 03 17 C7 65 10 D4 FF 60 8B E3 CD 8E 14 C3 5A 13
 D1 5B B5 0E C3 98 D9 FF 46 EE ED C7 BF B0 66 C2
 43 58 F3 B3 70 5E D9 89 9B 52 EC 93 3F 15 A7 2E
 8E FF AA 3A F5 0F 82 8F 4A AF B1 C7 0D D4 2A FE
 0E 39 EE 3D AD FD 31 56 F7 66 21 E6 01 FB 51 D1
 E0 7B 7F F5 B1 67 81 FF 04 03 A0 A3 6C FD D9 F8
 1E E7 7D 8D 8C 3C F1 2A 43 B0 59 DD 4E 4A 76 51
 E5 77 33 9C C4 6C 12 EA 35 59 F1 88 C0 62 4F 15
 AD 18 38 09 5F AD 88 AC EF FB 9C 2D B5 35 AC 5D
 72 F3 CF B2 48 0B 87 3E 43 D9 27 E2 7C FC BB 0D
 79 F9 CF 35 A2 56 A1 F3 AD 59 43 FD CC 51 60 DD
 1D E4 19 BC 97 A6 73 BF 69 F8 12 EF 3E 35 2A F7
 1D 7B 9A 71 19 FF 99 04 32 5E 4A B9 1F CC 55 9D
 AD E5 95 C1 44 AC 64 AE 51 3D FC 7A BC F9 8F 5F
 21 39 3C 12 80 38 E4 9C 48 BC 04 75 BA 29 2A 78
 5C 81 23 2E CE CD A8 DC 1D 06 AC 21 08 F6 4A 03
 D5 9D 79 A7 23 7C 6D B9 E3 D4 0C E1 01 7C B5 9B
 A9 28 8F 24 BD 07 48 B6 C0 0D BB D9 33 FA 61 D4
 57 5F C5 10 37 FA 07 13 40 E2 CD 12 A3 14 60 84
 0C B6 F6 1E 3B F3 65 AE DC 1E BF A1 10 E6 C2 30
 98 97 C2 2A 5B 80 F1 64 8A 1C D2 6F C2 B3 8D DA
 A6 09 69 6E 26 48 88 F9 A2 54 9F AD FB F6 EA 44
 DB 8D 1A 27 AC 79 AF C2 9A FA 66 CA 1C B4 78 63
 D1 2B 53 47 D3 F4 36 63 42 74 18 E0 9E AD 1A B4
 5F 98 5B 9A 23 73 FF FB B5 72 F4 86 16 99 52 83
 46 90 C4 9D 7C 51 E4 B5 E2 E3 5D A5 FE 3B E6 2F
 79 2A 64 75 78 18 06 56 ED 0A 7F 7E 8C 6E 59 F9
 6E 9C F6 9D 49 30 35 2F B0 1D A8 51 DA BB A0 7D
 82 6D 08 12 B4 53 3C 3B D8 E9 70 B7 50 C7 81 BC
 34 20 EA 5F 6D 0A 79 08 44 34 FE 80 A5 15 CA B5
 83 CC 93 26 33 0D 06 1E 77 E1 25 96 51 A2 97 C7
 C6 2F 43 37 9D 2F 70 3F 64 45 0A 7E 3B C9 32 BF
 35 C5 E5 70 9D 69 48 D1 C4 84 0D 2C 21 40 A7 14
 21 73 B2 6A 52 6B B6 42 5E BD 13 D6 E5 41 55 D5
 28 57 B8 FB 8A A8 25 20 BD F7 3C 02 64 B6 54 C8
 8A 0A 59 C0 5F 78 EF EA BD E4 5B BD C3 94 26 C5
 62 A2 AE A8 53 02 E3 0C FA 23 46 EE 5E B7 07 95
 4C 11 A9 57 79 9F 54 1C 4C 8B FC E1 65 C3 A1 D1
 79 53 8D 97 B9 24 6D 2D 48 6B 4B B5 F6 D0 13 D3
 D9 FA 72 A8 91 E1 C8 F1 50 EA ED ED EC AA 6D D8
 2D 10 57 C5 26 BE 8B DF 1F 27 97 B3 85 38 3F 42
 66 E6 FA 19 25 28 3E BB F5 D6 76 A3 CB 6E 46 A5
 6F F2 AC 38 AF D1 2F C1 61 F0 96 A0 EB 48 61 87
 4E F6 D1 79 40 A3 8E 1B E3 97 8E ED 94 66 BD 84
 43 8F 92 22 BD FA 1B 21 BD D4 3E 33 D4 C3 9F EF
 44 B8 FE 0D F7 88 ED 84 C9 84 A8 D4 78 90 CC A4
 2D CE 2D E7 42 D1 70 72 1E C1 32 F7 64 AC 90 9D
 AF F3 5B 91 3B C0 94 C2 6C 0E 76 DC 85 85 7C DD
 1F 0E 3F 60 DB 7F 77 40 FA D6 21 B1 B7 FC 85 6F
 9C E8 8F 74 10 94 C0 A9 25 36 42 B8 47 BC CD 2E
 E7 DA 7C 40 AA B1 BA 42 32 71 51 9B 2B AB F2 11
 DE 24 3A B8 93 7C 30 77 BD AA FC AE 9F 48 C1 CF
 EB A5 CD C8 DD FD CD FA 4D 3C BD 65 A4 0B AF 0C
 FC AA 9D 57 53 05 28 DF F9 95 D0 0F 01 B6 8E 61
 D4 E7 39 A8 12 20 85 2C 3B 1B A9 3E 55 CA 3E 6C
 B9 4C A1 55 21 CC 16 F5 61 7E 6B 6E C3 DD 76 68
 54 04 30 13 18 8D 23 75 61 39 3F 7A 33 CC 90 75
 25 B4 A2 F5 5D 8C 83 8F 7F 69 E6 47 45 48 4B 7F
 6F CB E1 3C 8C 31 59 20 C4 A8 D4 5E A2 09 BB 68
 88 BD 52 14 50 8E 16 33 7C B4 D4 C3 B4 06 8A 11
 B6 B1 0B 89 C5 FB 60 5E 49 F1 D5 81 15 01 17 D2
 D1 42 A4 A7 C4 48 A4 B8 49 B7 22 B0 D6 9F FA A5
 4F BC 10 F4 E6 F1 D3 39 44 2E DB 3D B7 2E 15 3D
 74 C5 AB 99 0F 3D 4C D5 DF F8 69 D1 A2 29 86 0E
 AC 71 E7 3B EF 1F 3B BA A8 81 3C F6 B8 2A 7D AA
 11 92 24 78 80 A9 D2 59 6B 2C C0 9D B4 81 B3 AA
 73 0E C0 D7 54 7C BF 70 2F 78 8A 09 0A ED 42 90
 F9 09 84 1F 26 60 93 42 CD 46 07 47 4F 63 D6 39
 E6 11 BB 9D C5 0C A1 60 D2 4F 36 14 88 49 9E 3C
 6D 2B AC 08 1C E3 83 4A 26 4C 8D B4 7C C2 52 B5
 3C BF B3 B7 56 9D A5 A2 FA EA AB 0A 93 EC 6D 95
 70 84 DD AF 68 7E 7B 0F A9 B2 3B 3F 86 2E 7C 0C
 E7 0A C6 33 AB 47 07 61 9B 05 2A 32 8D 60 9D 9F
 B1 CB 8A 9D 1F BA 57 2D EC 9D FB 62 88 B7 12 7A
 B2 C9 C4 EF 9E 85 87 92 6C 01 1C 5E 35 09 BD 24
 31 49 78 43 DA 5C 76 58 FB 7A 9A F6 0C BE D9 7D
 43 67 25 0F 1A 81 5D 46 15 6D 5A 79 DF 5C 33 74
 59 8E D8 D4 22 B2 2E B4 62 EB 14 AA 93 A5 93 07
 4A 1F F0 E4 66 E1 E4 4B 31 EF C1 CB 9A B7 EC AC
 23 F5 EF A3 0D 2F DF D8 98 A5 96 94 3C 99 7B D9
 73 1D A6 6F 58 2A 40 20 00 BA C1 8F 85 D0 27 C1
 49 B9 FE 56 84 23 B8 44 C7 9B 5B 76 10 3E B6 C0
 84 99 75 BF BD B2 A4 70 A8 08 F8 57 58 D2 3A 54
 61 EA 92 7C 40 08 9A 3D 40 9E E9 B6 FE E9 3A 17
 54 16 D0 BD B4 B5 18 EE 9D 07 C6 63 2F 84 0A 1C
 39 FA A1 9E A4 EE 0D 96 6C AC 7D 5E 31 1A 1E D9
 B2 3B DE 6F 68 F4 30 D3 FC FC 46 80 61 8E AF 5D
 F8 C3 6F 35 07 01 D2 F8 14 1E D7 A5 CA 21 DA 0A
 AE DD 20 8D 17 BF E5 5F B1 38 9B 8B 37 26 5A EB
 DE 11 77 A8 E8 63 12 7F B3 D9 A1 B6 14 4B 90 CC
 4D C6 C3 6D D8 C4 71 1D DB 2F FC 57 2B A0 C4 6A
 95 A2 40 D0 C6 35 09 BF F9 D8 EB 49 BC 0E 61 0F
 25 DA FA 50 D0 56 46 34 BE 4D 00 6D 05 66 C4 F7
 1C 41 A5 B8 AA E3 9A 76 71 8C 2C 52 55 01 32 BA
 43 78 17 FA 1D FA 5C 44 E7 86 15 30 AA F0 B1 22
 03 B9 D2 AA 50 11 9B B7 01 23 0E F9 4E FE 19 5A
 B3 EF 02 6D 77 EB 45 B6 D7 18 3A B3 07 BC 5A 24
 13 36 B1 3F CF 0B E2 0E BB 10 67 BC 1D 0C F0 B7
 76 71 16 07 04 2F 59 89 97 0E 1E A5 FA 95 C1 C4
 E7 B1 87 B0 D1 F3 F2 67 04 51 30 DA F3 88 3F 2D
 2F 96 07 6B 88 A4 51 86 C9 F2 DE A9 B7 CB 92 72
 C4 6F C3 B7 A7 C5 FD 57 7F DD 07 EA D7 09 E3 A7
 C2 74 26 BC 05 48 7D DC 0E CD 9C 46 76 22 60 3F
 BC 76 AF 8C 41 B3 D7 98 9E 87 5B 53 10 98 53 12
 75 D9 14 DD 22 16 26 58 B1 04 D6 18 F9 D0 6D 6D
 4F B0 2E CC 1A C5 A4 E1 3B B1 CB 84 07 A1 33 80
 A1 A2 89 2B C8 33 50 7A D1 C7 7B AE 4D 48 E4 5C
 DD CC 6B AC 65 55 00 6C E7 FF 54 7C AE 94 B4 DA
 61 35 1D D7 10 2E 6C 83 89 84 CF CF 6B DE 4D 23
 19 2D CB 1B 51 03 98 66 49 D0 CD 32 54 7C 72 DA
 63 71 70 24 6A 10 F9 0B 5E C7 8A 47 53 FE 9B FC
 7D 10 42 58 78 A8 7A 54 57 23 53 5F 13 C4 FA 70
 0D 27 E2 26 9D 6C 58 38 26 47 24 20 FD 64 17 30
 83 07 6C 8E 72 33 AF DC 61 35 37 41 8A D1 B5 51
 12 5D 28 F4 8E A6 61 37 71 1B BA 22 69 92 B5 82
 CC 34 44 AC 93 A2 AB FF D9 AF 7C 6B 4C 5B 99 9F
 76 24 79 15 BA B3 27 73 2A 44 32 95 B8 6E CF 64
 DD B5 07 D1 AE 4F 38 E5 2F 9A CC 8D 6C 82 95 29
 1A CA 90 14 C9 0F B6 8C 05 F9 28 B7 6E 24 66 2D
 77 60 DF D7 96 57 A3 56 C0 53 EF A9 9B BA 0A E8
 DE FC C7 56 33 71 A1 21 9E 3F AD AD F8 DD A9 25
 7F 31 9E 8A 96 DB C8 C1 F2 75 D6 FD 71 4F 17 DC
 5B 77 F6 8C D5 92 9D 2B 50 2B AB 26 EA 92 F5 BA
 B8 FD 49 CC DE DC F8 74 A6 4A 3F F0 65 B1 7D FF
 0C E3 CF E0 F9 A8 6F C0 2F BA 70 6B 11 EE CB 67
 8C B1 6E 5C B1 D9 3D F3 0C 7D 0A FA 71 4D AF B6
 C0 9D 4C 4B C2 A8 B3 B7 D5 67 AC 62 46 74 41 D6
 34 60 D2 92 9F B9 40 3E B5 61 DF EE 17 A4 8E D3
 9D 3E 55 A6 A3 9E 05 AF 54 54 ED 7E 82 9A FB 1B
 A0 8E 21 18 D7 C1 D1 F7 24 1A 73 4F 49 3C 88 4F
 E9 85 17 25 5F 77 D6 EC A5 7C 08 53 1A 0F D7 46
 59 AE 6A 39 7D 7D A3 1B 93 BB 21 CA FA B5 57 28
 A3 B9 11 65 81 6B 03 9B 4A 6F 8D ED 14 01 BA 04
 16 92 17 F6 50 50 C1 84 39 62 E7 DA 8A A5 A2 77
 26 97 78 BA 58 3F 26 35 7F 89 1F 8B 4C 95 F5 C6
 7A B9 3C CB 74 39 DB AE 46 C4 52 22 E1 72 63 27
 7F D3 CA E5 6C 38 49 58 1E 4A 11 A2 BD 29 B0 E9
 82 40 AE 50 48 9A B7 21 D3 C6 FD AD 6A 72 60 F2
 BA A8 F3 6C E5 30 3A FD 1D 16 7E EC 90 E3 CA A1
 43 BE 45 1F 72 76 1D 5C 04 0F CE A3 E6 0B 6E C7
 AB 62 84 3F A2 21 95 C6 BA E2 DF 67 A8 7D F1 91
 5D E4 40 37 AE DF 9E A1 19 47 3E B9 0E AA 7A 03
 8A 3B 2C 4C 74 B3 5F DC 21 05 04 35 F1 49 8D 40
 CB 68 28 74 E1 D5 A6 1E E8 85 DB B2 6A E0 05 A9
 39 15 B0 71 22 D6 F9 2A B3 F3 80 48 4C 8A D9 CF
 62 5D 52 01 A4 FC 0A 35 95 6C 37 66 24 25 40 8D
 FD 11 A9 C3 AE 13 59 5E 10 7F 9D B5 15 2E 0B C4
 30 32 2C D7 52 4D E2 A0 E8 22 FA 1F 7B 36 E6 3A
 47 93 E9 4B C5 43 08 F5 EE 56 F9 EF C2 AA 77 0E
 23 BD 0E CA 59 3C 6D 96 BB 89 18 BA 1A F3 33 10
 3C D2 DD 7F 5D EB F1 58 3D E2 3D 2A 4A DB E3 2E
 29 B1 81 81 C9 30 64 43 C3 72 50 2F 85 C4 EF 5A
 2A 79 C3 8F AB 2A 82 5B E2 DD CC 9B 00 57 F5 49
 F8 ED 12 50 94 8F 89 CD 3A 7E 36 C1 D3 E7 AE 27
 B7 B9 AF 33 0C E2 71 E9 BC C6 16 86 6E 10 BB 43
 0E B7 A2 98 49 5C 42 05 CE CF A5 B2 83 97 ED 3A
 96 F1 EB E6 D1 B5 1C 2B ED 3E 62 9E 84 76 BE 26
 1F 49 8A 82 96 80 B0 58 3B 34 12 65 13 EB C5 65
 22 F2 47 8B F0 C5 CB AF 31 CE F6 C4 E2 D4 3C 36
 C4 61 02 F7 EA 0D CF 4B D6 1C 6E 31 68 A3 68 1F
 B3 9E FE 17 DF DC B6 40 10 5C 9E ED 6F 01 FC 51
 9A E7 3A E4 39 7E 32 C6 EF AF 40 4E 4B F5 52 5B
 A3 22 5A 06 8E 2E 67 F3 F5 41 B9 7F 99 3D 60 4E
 16 EC 50 79 B9 C1 DC CD 9F CA AA D0 2D 18 B1 D4
 0D B0 15 DB 67 B1 1E B0 E7 8F EB 6D 39 93 25 BF
 57 2B D2 F5 38 30 3E EE 72 23 BB C9 58 98 15 77
 8F AC E4 A7 87 49 D6 AE 93 3E 5A 64 65 C3 7E E2
 E9 2D 8D 55 71 4D E4 43 23 00 ED A1 99 CB 17 3B
 7E 64 47 CF 50 74 E4 A0 76 BA 3D 8F 3F 48 BE 71
 66 1D B5 B2 70 BC BB 00 FA 5F 7A 28 4A 54 0F CA
 F4 FC D1 1F 3A 05 74 C5 00 30 06 8C 98 89 85 E3
 AA 50 F9 A7 A3 8F 07 04 5E FE B3 97 5E BD 93 FD
 57 02 BB CF 71 6F 37 C8 CE 7F 5C 3A 31 86 8E BC
 04 A8 5D C5 3F 98 50 C4 D7 DC 6C 4A FA 04 56 52
 5A E0 01 75 7F D4 30 1E 09 21 B5 E2 63 ED A6 0D
 42 77 DE 4E 5D 4C AB 07 47 B5 AC 8B 8C 5D D6 ED
 89 03 0C 99 23 56 63 2B AE B0 5A CF 17 24 4F DD
 87 C8 E7 C9 12 F4 C1 DF 16 2E 45 66 FE 82 0B FF
 25 9E 72 6A EE F6 26 BB 0A EA 82 F2 0A C3 50 B1
 88 8B 47 E6 22 8C 85 3A 1C 4B D8 44 01 54 0F AB
 7D D3 DB 9F 2E 34 21 64 28 C6 28 F8 3F 08 8B 3B
 57 71 99 DB 25 B7 4A F8 A8 2C C9 2E 63 31 6A 9E
 53 89 21 2C E1 D1 89 C4 CB D7 AF D9 5B B8 E3 81
 DC 08 6B 40 20 E9 48 A6 12 36 5E 4C F0 CE A7 21
 C3 F1 A3 1B 19 5A 83 67 E6 E8 92 9A 6E CC D0 5A
 E7 4B BB A7 D9 9F 8B 9C 2B 11 4D 88 DE 12 4F 65
 87 52 73 A5 4B 5B C9 DF FB FC 12 B0 B7 E0 9A 04
 56 0E C4 9A FE 0A 84 87 12 EB 5E 7D 5A 51 76 00
 50 82 2B 70 7B 28 EA D4 38 28 AF 77 32 73 68 7A
 29 B3 64 E0 1C D4 15 9D 06 6C A7 2C C4 CA 14 67
 52 42 80 15 69 74 54 2C D9 A4 ED DA FE 75 03 18
 F8 A1 9F 1F 42 EC 48 0D 9C 28 24 E4 40 3B CF 82
 18 68 DB 7C 46 5A F2 69 12 CC F9 54 72 F5 AB 9F
 6F 82 D7 22 F4 04 BC 70 7C AF C9 44 E6 AE A3 D0
 0A 91 2D 6F 9E 43 27 59 7D 82 E6 AB 9D 1D 1C B4
 79 5D 1E CD 3E 62 2A 42 43 F8 AE A0 DB 5B BD 34
 16 45 C1 02 26 FD A7 F8 3C 75 55 14 93 2C F4 59
 AE E5 54 3F 96 87 FC C4 80 30 32 C9 3A F8 62 0F
 48 CA BC F7 2B 50 05 4F 10 03 34 C9 46 BD AD 1C
 8B 5D 35 96 1A C3 69 DE 74 D4 CF E4 B2 B8 6C 92
 90 CA 0F 6F 30 1C 84 53 46 BE 41 BD 2F BD 5A ED
 C0 D9 1C E5 67 05 8B B0 49 D1 F0 6B AB 7D 92 96
 20 91 A2 9C 84 90 3E 52 AB 45 56 6F C7 D4 FF E7
 C7 2A 05 74 F4 F3 EA FE BD B0 D5 E6 D9 DD 08 A0
 A6 F8 5D 32 E1 FC BB B7 E3 BB 85 76 BF E1 8E E9
 F2 6C 68 2A 7F 4A 72 59 2F 90 51 A9 E5 09 B2 1A
 64 1B 6E A7 AE 3F FB 10 CF 38 98 9C 4B 51 47 72
 2F 13 BC 2F 2B 56 83 5E EA 66 70 B9 A5 EF BF EC
 E8 0C C4 39 2C EF 0F AA 4B 4F 3E 3F 60 06 43 2D
 B0 99 93 A3 D4 02 11 3B 01 DA 8C 3B E4 13 15 67
 7C CE 22 8A 75 5E 2B B7 CF 0F 2C D3 64 47 38 1C
 0D BF B8 15 F8 FF 6D F0 E4 31 B3 1F D0 D3 CC F1
 21 EF 28 18 D1 20 F5 B6 50 8B 32 6D 0E AE D5 FA
 69 4E C7 A9 19 1A 3C 76 4A 4F DA 2D 16 16 B5 E6
 B8 82 86 87 BA D0 C9 24 90 E7 18 24 29 53 4E 24
 03 9B 75 5B C0 51 0E 23 42 D9 BB D1 3D 35 BF 79
 3E E0 B8 A6 72 EE BD C6 CF 8D 87 80 30 84 A2 C1
 74 FD 5A 92 E3 83 26 A6 98 E0 58 6F 57 A8 1C 58
 D7 01 B0 F4 D1 89 19 E0 FD 20 5E 9A 49 4C A2 54
 20 98 96 98 E3 26 55 99 5D 21 C4 B8 0C 19 A2 31
 55 84 1E B2 4C C6 36 3B 38 24 FC 1E 34 B5 A9 65
 42 34 CF E4 B0 77 0C 93 D7 FF 8B C6 67 97 02 63
 BB 93 F1 F5 B0 EE 08 8D 8F 7E 3D BA 44 17 E3 0B
 98 0A 0A 8F 3D CF B2 5A 10 82 2B 84 78 C1 0C 3D
 91 98 5E 65 7C 64 11 BC 10 48 7D 08 CA DB F9 28
 A0 22 4A 35 4D 58 B1 AA 42 9F 79 0C F9 6F E9 1A
 24 11 F4 71 76 F2 6A 3C 44 63 2E 24 21 77 82 9D
 D1 AE 70 AA 53 F1 44 AE 34 D5 23 33 A2 D7 83 10
 90 39 12 BB CE DB F2 97 6A 04 C5 31 AD DE B6 DA
 1F 30 5E AE 1F 13 6C 06 C4 F7 9A 9D EB 23 16 29
 78 1D B5 AA 78 E2 F9 E1 4E E4 0B 4C 07 58 A5 C1
 80 AA 51 D9 F7 07 A5 C9 9E 05 92 7F 94 6A D8 D2
 E0 1E B8 3F 8C 1F A4 90 AA 1E C1 1D 80 47 76 4D
 16 2C A5 B1 6A 02 2C 1C 05 67 AC 2A F7 E2 8F 58
 ED 01 A7 81 D7 BB 0B EF 49 E6 E6 CB 3F 09 C2 94
 3F 9D 16 49 C7 23 08 3C 1A AA 27 76 DD 87 88 25
 40 3B 52 39 7A B0 8A 17 59 E0 58 08 61 5B 97 85
 EB BB 76 FB 12 3D EF DE E4 32 29 F5 A2 BB C5 7A
 C3 51 77 69 40 51 0B 0B 10 CE 79 4A 59 8E 1C E5
 91 2D C1 71 8A 75 E5 66 2C B7 4C F8 1F 7F 9E E1
 2C 84 44 7B C6 CA 58 B6 E2 C0 39 94 D3 2C A2 4B
 AF E8 74 D8 92 7E 70 90 AA 37 D7 5F 2A BD 6B EE
 C6 E5 0A 35 2F 6C E0 C2 9E 5F B5 50 5D 56 36 0C
 C3 0E 03 9F D7 40 2A AA 5F AA D6 17 87 9C B4 60
 F4 A9 6D C8 1C 48 62 6D DA 3A 56 37 14 B5 B0 77
 18 BE 8F 5D BC B8 33 20 6C D8 72 98 6D 9E F1 CE
 D2 07 D2 F5 B0 CA 30 34 32 07 DF 82 EA C6 88 5D
 F3 3E 33 6E 52 1B 2C 68 68 E1 80 FE FF 4E 66 27
 92 CF 09 CD E9 D1 04 3D 5E 2F E4 C2 13 3B B8 18
 71 05 0B A5 B3 65 B1 3F F6 75 24 88 73 C6 BE 99
 8A 32 CB 72 9C 4C A5 B7 92 31 43 9F FA CC C3 A6
 3C B9 40 54 43 12 86 3C 9D F5 B8 DD A4 35 81 8D
 83 67 5F 8C D9 F6 7E 99 E0 A4 F9 CB 7F 4B 13 E1
 25 15 69 CF 9B 16 90 A0 5E A1 58 7B 51 FA 41 DE
 7D C2 8F 70 D7 7A 6B F5 6F 88 BC 4F 66 FD 78 0A
 13 5C 39 86 17 86 FE AE 59 81 7F 50 AB A8 C0 C2
 0B B0 9C F4 30 11 DA 0B 0D 18 CA BA 31 0C DC 82
 C0 D3 00 3A 0F B5 71 73 95 27 3D 36 37 32 92 E6
 B0 7D B6 50 6D E2 C8 00 39 E8 45 F6 3F EF 8B 55
 4B 2B 79 85 04 F3 0F 41 1F 50 EA C4 7D CC 14 6A
 48 CC 00 54 41 02 5D E1 B0 05 35 BA 43 B7 A1 D5
 36 DA 58 43 77 03 DF F2 36 DE 0E 3C 11 2D 61 8A
 4D 72 A8 02 E4 F3 06 E4 5A C5 5C 4C 7E F6 C3 9A
 6E 0F CD 7E 30 D0 02 FD 64 9D 30 CB 1C 02 35 89
 64 0A F5 7E 2A 16 76 AE F6 1D 72 4E 7A 0C 5E E7
 75 E7 ED 43 AA F0 39 CF AE 52 0F 6B 78 63 42 4B
 51 33 CA C3 C2 24 64 5D DE 4B C8 D9 BC C7 F6 DA
 7D 9C BE D0 CA A0 ED 0C 56 C8 E8 2F 74 49 35 28
 E4 68 A7 7C D4 84 AC 03 6E EE F4 94 CE 6F 03 47
 F9 E9 21 91 81 3C 32 25 C2 C1 09 81 98 0D 01 34
 AF 04 04 C7 16 43 26 9D 24 24 B5 DC B6 CE 99 CC
 63 F7 0B 35 D7 F9 1F 0F A9 36 D8 DA 43 41 CF C3
 84 1C FC 9F 5C B1 17 6B 19 FE 61 F0 76 29 27 9F
 6B 22 02 DE 99 C2 EA F2 FC 55 94 03 6C 09 FC F8
 46 40 75 02 21 61 A6 16 69 8D 55 5D C9 56 2C 0E
 60 21 C0 FC 2C A1 5A AD 73 F4 10 6F 9A 00 D1 E1
 25 5E 7A 53 F0 B0 26 F8 93 F3 5D 99 CA 56 31 62
 F4 88 C8 AA 83 76 32 D0 9D 21 B9 7E 71 99 9D D0
 56 AC 64 C3 50 08 07 4D E8 FF 63 4C 24 6F A7 43
 F3 DD B3 0A 70 6F 74 68 79 1E DB 5D 58 3A 2D 4C
 B7 46 BA 88 31 B1 93 2C BA C4 41 95 16 BB 69 C0
 15 8E A6 18 C8 90 58 D4 6F 20 70 69 17 FA B7 2E
 B6 E6 17 EE 45 47 68 F9 75 13 E6 A9 AC 0D CF 0F
 E2 77 34 A5 21 20 46 43 5B 82 B8 59 A8 C6 84 8E
 2D D4 F3 4B 9E A1 95 0F 30 30 B7 34 C7 36 A3 74
 6C 9A 5F DC 3E F3 14 82 7E 80 D9 1D BE FA 57 7A
 69 10 44 FF B8 3E 40 EE 1D F7 D8 CD 4B 5D CC 6B
 78 0F BF 27 9A 7E E9 EE 84 67 A3 6C 4E 10 79 E2
 63 52 43 26 B8 B6 2B F3 24 77 66 F0 4E F7 61 36
 89 C2 FE B2 B6 36 44 BB 44 5B 9E 1A FF A8 FE 6C
 21 3C ED 16 00 22 89 30 6B AC 53 F8 C0 92 E4 A9
 39 C6 C1 A8 BB E8 80 1E 87 15 8B 12 03 CB F1 65
 22 04 93 F6 BF AF EF 12 39 A6 39 EA C8 8A C0 65
 0D 0D 83 93 D4 38 E2 8A CD F1 F1 6D 6D 0F 4F 05
 C1 A3 16 DB AA 73 D7 8F 72 87 0D 5A 19 B4 50 88
 CA 64 B9 36 D4 89 26 31 C0 4F B1 00 88 A5 17 3C
 F7 CE 6C 37 24 ED BC 88 D7 03 62 32 09 C2 A0 F9
 5F 46 6E 56 06 94 2F 04 02 B5 17 F4 D5 02 D7 25
 7E 3A 6D B4 C7 C2 DE FF E4 6E 8A C6 BD 87 A3 3A
 1A 09 FC B1 CF 22 48 B3 2C 34 6B F1 AE 94 1D 9E
 8D 94 91 7F DD B3 B5 B9 95 CF A3 04 5F 7D F7 A8
 7B 7C 9A 14 7E 6B 87 2E 09 18 EE F4 74 72 8A B2
 43 4C EE 74 F7 52 17 BA 17 2C 74 DA 44 7D 1E 4D
 FF 20 94 82 40 E7 64 EA 6E 3F 15 7A 76 18 63 06
 70 6C 5F 9B E6 DA 14 66 C1 7F E1 B8 12 22 E1 1A
 98 E2 78 A0 99 C3 71 5E 03 55 1B 05 10 2D DC 4A
 1D 8D 82 BA 66 24 4C 97 B7 22 0E E1 23 D1 9C AA
 F4 48 28 57 3D E5 E4 1C 6E F2 CC D5 3E 5B 37 DE
 E3 65 98 A0 2F 2F 06 CC 29 F7 6D 01 3F 6D 13 E7
 98 33 55 27 90 70 FF 9F 21 AA C4 D0 A4 B0 25 D6
 8C 46 4E EC 84 AA 2E 06 1A EB 2B A6 53 7D A9 4B
 01 F3 AA 29 BD CA 28 B3 1F 6C 3C C6 B3 33 C8 19
 07 FB 48 62 29 26 15 8A 9F 2A AC 77 84 D3 B7 77
 0B 61 7A B3 3D 50 E4 8C 41 56 BA BB A6 92 F6 F0
 BB 78 AB 28 20 E4 39 3B A5 B5 2F EE 77 0B 19 0A
 ED BA A2 6C B3 B0 DB F4 96 96 24 CB B8 A0 9A 78
 6B D7 C4 E2 AA 13 F1 07 DC E4 D7 D4 11 8E 22 CF
 2C CA 11 84 1F F1 AD CB D7 BE 70 DA EF E1 7C 61
 DD 92 B0 64 96 40 52 65 5A F3 B6 F4 CD 30 16 49
 E2 E8 96 D4 E7 64 06 F6 02 96 3E B7 5C DD 48 65
 B9 85 CC 18 36 4E 31 95 67 19 A1 E6 50 D8 A4 78
 1F CE 1C 09 50 4D 27 AA 6C EE A8 71 D3 21 BC F2
 8C C7 C8 39 84 98 36 74 92 AE D5 BC 09 B4 1E E3
 E8 7B C1 95 8D 41 C7 8E AF 27 E1 E0 DC 8E 59 8D
 50 51 34 E5 1D 66 09 7F 68 EA 5C C1 8D 55 66 5F
 6C C3 C4 FF F2 4C 77 03 B7 27 A9 AD 5B D9 CD 1F
 B9 95 15 72 63 C2 45 2C 27 CA DA 16 8E BF EC DE
 48 CF BC 75 27 0F E6 A6 6A C9 96 0B 5E A3 D2 BA
 20 B2 DA E2 D1 91 B4 B4 7A 47 47 09 2F 86 7F 66
 12 FE A9 BB 87 85 1C 2E 8D 6B 3C 85 8B 00 1F B4
 38 4A 6E B9 9E 7B A5 97 81 22 E1 A8 5E A5 47 6F
 0B 8E 9B AC 4C 7C CF 84 BA 69 D3 69 D0 60 22 C0
 E6 C7 44 4D 29 CE FD 2B 36 9F 88 44 54 75 EB D4
 BE 26 D3 BC E3 D2 C8 C3 A3 85 0D F7 34 E8 6D EA
 E1 DD E2 2A 1B 2D CD CB BE 8D 95 45 29 18 81 F3
 27 58 60 BE D2 C9 39 6A 5F CC 80 5C E6 F0 52 D7
 D8 2C 07 1D 5B 6D 3B 02 9B 04 B7 B9 04 F5 48 BD
 24 04 11 5F DE 3A 09 DA 44 5D DE E5 A5 A6 69 64
 75 26 8D 08 11 2B E6 87 D9 5D DF 8B E0 AC F5 7F
 64 87 48 09 26 D9 90 BA C8 14 0F 7B CD 60 9F 67
 5D A0 7F 6B 04 63 67 97 DB 43 9A 6B FA E4 5E AD
 A6 5F B7 21 7B 1E D4 4B B4 0A 2B F5 71 3E 48 22
 0D 0C BD E9 D7 BE E7 27 34 B5 33 16 06 44 B6 88
 0B 83 A9 78 E7 25 45 94 E8 A4 1E 40 85 81 9A 15
 53 10 84 7C 47 F4 B0 1A 03 DB 29 3D 15 50 F1 2D
 89 C3 5A 87 64 6B 68 6C 4F 69 26 B0 99 4C 62 10
 7E 5C 50 F6 C3 C0 AF 34 D9 98 4D DF 42 48 79 A6
 C7 2E 59 28 DA D3 48 6D 0F CE 5F 08 3A 74 BC 77
 B9 A6 BF D2 BD CE 13 AB AE E2 0B 20 E0 9D 67 56
 7F D6 5E 1E CC 1A 1A 11 B5 9A 03 C3 42 47 CE 37
 7F BE B3 24 A9 3B D4 44 03 F7 AA A9 D1 92 AB 7D
 76 B3 1E 8C 69 42 5D FC 2F 28 47 66 42 9E 33 B5
 3F 5F 59 A4 A8 3F D9 74 06 64 83 A6 3F 45 1E 78
 FE 4F 80 DF 5C 6A B1 C8 86 2C 15 FF F8 0D 11 DE
 30 93 F6 D8 72 9F E9 FC FD 2C 68 5B 58 81 C8 01
 C2 B8 6D D0 FC 3C 31 E0 20 9C 92 EF 2E BE 69 A9
 77 BB 6F BA 87 88 F3 A1 A2 CE 67 69 90 45 1D D5
 A8 15 A1 43 A2 70 97 57 11 C8 1A 58 66 F8 6E 51
 A7 85 7F 92 0D 65 DE 54 E9 54 C9 A6 35 F9 96 62
 1D 87 CA 51 C8 A5 16 9F CD 3D E7 FF 8B DE 9F FB
 7F 52 7A 86 97 8B F9 39 1A BF 6B 38 B4 89 3A FD
 CE D0 31 8A 94 62 DB 61 FC B4 36 87 7B 14 5A DA
 BD 24 A6 B4 88 3E F5 9E 91 FD 21 41 B4 50 10 5B
 EF 45 61 16 C5 54 99 23 C0 ED E9 2E 6A E4 66 2B
 B8 09 9C 37 59 2E AA D8 55 62 72 37 A3 E0 A7 B5
 61 3B FE A7 44 A9 2F 66 AB C7 7C 57 1B E8 7E 7A
 60 90 23 1F BB 96 9A 95 CD F9 27 14 E1 78 EB C7
 82 25 1D 36 5F 8C 3F 4C 76 8C 2B 7C F8 BF 42 12
 70 6D 96 D6 9C AA 9E 46 57 7C F7 AF B0 F0 71 8B
 1E BE 88 19 C6 B4 C8 70 5D 11 1F C7 91 DC CD 3D
 A2 08 71 E4 3D E2 CE 3E 63 8E 87 A1 58 F0 11 74
 44 2C 64 9B 6B 66 7F 58 24 B2 9C 90 BC 61 9E 9E
 7C 4D E5 0F 4D FB 56 36 30 4B F4 3B E0 F0 70 41
 64 0D 31 65 15 E3 38 B4 6C 6D A6 BD A4 66 A1 F4
 6F 36 B0 9F 67 35 B9 8B 11 47 0D 0A E2 E1 C3 4E
 E1 AE B9 71 6F C1 04 94 86 21 55 0C C5 C0 76 C4
 E1 9A 77 D9 C2 CE F4 76 6B 50 E7 90 FA 55 19 4C
 98 1B 6A 10 D3 DD F4 A3 ED 1A 2C 05 60 FF AF EE
 DA F9 1F 94 73 CE 6E 52 3A 35 24 33 3F 95 FE C6
 C7 9B AA 64 91 33 1E D7 94 7F 1B EC CE AA 8D A5
 DF AA 8D B4 71 39 4B 77 C8 E2 57 89 4C 07 06 43
 9D D8 4A 06 E7 B9 D7 23 87 5C F2 48 E5 22 C3 09
 14 7E 5F AA CE 21 DC D9 6C B7 EB D7 2D 98 95 0A
 C6 E8 ED C9 1B 0A 2A DE 68 80 B7 0A D5 0C DF 44
 0B FB 3A D0 95 8A 40 1B E7 04 CA 85 06 93 B0 D4
 FD E7 40 A8 44 BA 9E 63 76 EC 71 BD 13 BD 27 8E
 14 E6 D4 E5 B7 73 FB B7 D7 83 3D BD 9F 91 56 EA
 BF 9C EC 83 60 D7 45 4A 78 33 36 0C 74 D2 F2 7D
 2F E2 D0 A6 B0 C2 76 5C 2A F8 B7 BB 20 2F 55 F7
 91 E7 69 E0 BB B5 4A 82 D0 F6 0F FF 29 11 E1 08
 8D A3 35 6D 72 CE FB 3E DB 9D 8F 12 4E D0 DF 88
 B0 3F A1 50 A8 FB 5F 76 31 04 41 B8 82 DF 47 21
 A0 C8 DC 22 25 93 D2 AA 79 D7 AB C0 0A 49 C4 64
 FF 5C 83 08 2D B6 F2 E7 6A 1D A2 40 D0 A8 82 D7
 14 50 1C 55 49 2F 53 6A F5 A6 F3 60 A3 9E 0F E2
 C6 67 0E 49 B3 D0 F2 57 7B 09 F5 0D B1 23 18 B4
 62 65 E4 EC 41 D6 C1 4A 91 63 35 D2 10 D8 71 79
 AB 5A BD 25 BF E3 03 84 A5 92 42 6C 7F D5 45 87
 31 57 AC 50 B4 6E 9A FD 11 4B FC CE 4A 12 74 36
 1D B1 0A B7 F7 1C 4F 8E 92 04 B9 BD 58 D4 C6 F3
 8E 77 48 31 44 7A D1 D9 9A 61 89 7E 5C 4B 06 3D
 0A C1 44 4B CB DC A5 A4 9A 35 56 45 0F 4D 14 FD
 88 ED B3 68 80 8A 28 38 41 8D 02 88 E2 5F F2 2B
 E0 7C C4 85 06 FE C8 C7 B9 9E 54 21 CF 34 21 78
 51 C0 21 D6 35 A0 45 A5 70 DE FC 7E 6D 82 E0 20
 C4 BD D3 C3 B8 FB 6D 26 77 55 A1 D3 7E FE 64 40
 AF A6 B3 75 A0 64 46 F9 BA F8 45 99 FA 68 0F C5
 AE B6 CD 1B 39 81 E4 50 F3 BA 4C A7 3C 8B C5 4E
 A2 6F 5D BC A8 AA 8B BD CC B0 23 F1 BD C7 8C 67
 1D 3D 51 21 EA 0A 7F F6 11 04 92 44 81 1E 6E 37
 C0 54 D5 2B B7 1A 6F B0 BC E0 A8 CC D5 04 4D D7
 65 7F C3 5F CE 3D 3B 9A 52 81 71 99 F6 BB E8 B4
 2D 3C DC 29 D3 B4 7D 7E 65 C2 54 B1 C5 1F 6C B7
 3E 12 C3 41 88 E9 F5 28 42 81 8D 77 30 F2 04 8D
 23 D4 FF 87 90 5D E4 0D 46 B9 2A A4 F3 7A 2E 83
 F1 9C C7 DB 33 88 43 87 97 B2 73 5D C6 5A 28 67
 C8 B2 F5 67 18 1C 4A D0 73 C9 86 FD 75 F8 B6 6C
 89 7E 1A F7 57 79 0B 11 34 5E 04 C3 BC F3 96 88
 93 4C 40 5E 29 8D D5 E1 6E D0 77 61 A5 6E BE 6A
 DD 69 F0 FD E8 86 C5 36 CA 7C 37 39 A6 D6 A3 84
 C8 5D F3 AF 66 F8 A4 78 AD C5 95 96 62 A3 38 58
 53 E3 F9 80 22 B7 2F D7 F6 1A 62 9D 19 94 36 3C
 5A F5 28 16 F8 29 61 47 C0 E0 18 CF ED 84 32 3A
 A4 82 2A D2 7D 18 8C 5D AB B5 8F D1 50 3E 31 C9
 38 D6 D9 79 81 5E AF 89 7E 95 1B D2 C2 45 3C 83
 59 C7 E6 65 E7 FD 6F 4C 1F F1 F1 10 8B D9 37 40
 1E 08 47 34 06 4E 3D C0 F6 62 47 D1 54 DA 19 45
 68 3B A8 78 27 E8 57 C5 9E 5B B6 F6 19 19 84 08
 88 DC E6 54 7D 57 93 76 3C 84 67 68 74 5C A0 B6
 07 B0 6D 78 7F FE B1 E2 7F C8 95 A6 A0 33 12 40
 39 17 A4 AA 0E 3C 37 56 A0 65 47 58 50 D9 D1 FF
 82 94 E2 6E B0 14 44 35 AD C8 F2 8F DC 79 8F 0A
 C2 DB 99 D1 1D 83 AE 69 63 B5 31 B3 CF 20 01 39
 84 AD C0 7A 94 F1 5B BF E6 19 BE 4D EB 04 28 5A
 9F 56 D3 2F 7D D6 D0 8B A1 37 59 73 6E 94 29 D0
 B1 54 0D 60 C7 2C B1 78 73 69 A7 C2 04 3A 5A 08
 D1 32 6D 60 D4 98 99 7F 17 0A 72 FD ED 65 8B 56
 89 DF FE E4 A6 3D E8 FE 95 1C 55 69 A7 E0 50 8E
 2A B9 A7 2D 43 91 8E F4 C3 12 DA D9 42 10 14 67
 33 1C 80 34 05 FA 3F 1D F0 97 2D FA 5A 99 94 F7
 7A 58 17 AE C6 89 7C 7E 36 8D EB B4 EB D3 5A E9
 12 35 CC B9 A5 14 43 B2 E9 B0 84 29 BA 40 FF 75
 19 EE A8 45 FB A6 55 34 55 7F 73 9E FC 9D 04 2A
 7A C9 27 CC B4 50 2E 36 4F FF 48 F8 79 73 72 EB
 1B 16 95 A7 DA DC C2 A2 76 D3 35 35 B2 03 73 8E
 61 96 4D D4 87 B0 CA 75 F6 6F 9F 02 C0 3C 46 7C
 9E 17 32 5A B4 F9 4A A0 D9 D1 A4 1A 46 B7 89 29
 55 4D 32 3E 85 16 A0 8E FB 5B EC 43 36 7A 6D B0
 EF A9 5B C6 51 A3 33 A5 74 2D 77 D5 6E EB 51 35
 6F 21 A0 C6 EB 01 A0 4D 6E 48 A5 11 21 98 A7 C9
 F4 26 2C 66 F1 C9 60 38 90 EE 06 21 CC 36 3C 39
 72 C4 34 49 32 A0 BE 74 58 BD 0C E9 76 00 57 7B
 2C FD 03 CF CC D3 E9 C1 C9 EE BD D2 49 39 67 99
 FE FD DF F5 72 C8 AF 2A C0 10 03 5B C1 DF 15 EF
 7C 24 FA 27 54 76 5C CE 05 DF FF A8 D5 CC 4F 84
 40 9B 4C 0A FF 9E 72 DA 6B 07 43 B7 37 BB 13 06
 42 62 91 29 9E 15 4D D2 26 2F 78 6C 4D 0A AC 16
 94 F2 FD 57 84 78 04 1C EA 0C 6A 6B 67 4C F1 DE
 56 FF 32 AB 9D C6 6F 4D 6B 41 CE A8 96 06 DD 29
 29 ED 22 C2 10 D5 5A 18 C8 29 93 73 76 BC 26 81
 BD 1F 6B 78 B6 AB 7A F6 47 81 C1 17 E2 2C D5 70
 A0 A6 1F 7D 03 20 8E A0 9C 23 C2 BE DC BF FA BA
 24 EF 65 E1 D7 26 99 33 F6 34 BA 58 7F DD 04 5C
 D4 DB 4D 88 87 FD FC 62 F4 54 81 8D 1D 46 95 2E
 3A 37 0E B2 2B 97 FE 52 79 50 18 2D E3 02 C2 55
 96 17 B8 C4 E1 17 A2 1B 1E D5 39 AF C8 E0 86 E3
 11 61 F2 98 A8 B5 0C 1F 7A BE 38 A9 67 6D 9C 97
 E0 E8 7E 89 95 CD 5E 74 79 0E F4 98 FF 86 C9 AC
 A9 FE 49 19 D8 1E CD 9B 4C 97 7B 77 04 89 5C 8F
 94 8E 40 14 9B 08 B6 B0 48 90 CB A4 2E 5C 6E B9
 D8 B2 DA 88 FA B6 EE 6A 18 04 CF 02 C6 BB F0 10
 97 D2 B3 02 FF 33 8D CA A5 86 9E 8B FE 2C F5 CF
 FF DF E3 9E 82 A8 FA D6 B1 D5 06 0B A9 A4 87 DC
 00 12 92 0F 50 8B 22 DA F4 38 00 D6 E0 37 D3 3B
 53 4C F3 F0 56 C2 0E 89 FE AC B3 38 3E 53 A8 C9
 E3 D9 00 7D E2 FC 0F 1A 66 35 A6 3C 70 0C 7D BD
 06 AD FA 82 E5 2C E4 D6 49 4E 1E 7F 5E 04 F0 BD
 97 CC BC 2C 8B 93 76 42 7A 6B 60 E4 F1 91 EA 54
 0B 22 DC A1 04 4A F8 78 5C B7 B2 BC FB 76 63 04
 19 EC DC A7 EE E8 1E 71 6E 8A 57 D5 09 67 51 CC
 56 2D 4A 44 15 4A 74 A1 8B CE E6 A3 CD 50 F9 AB
 D2 7E 88 DA 5C 42 44 3F F9 11 F6 D2 6D 7B 9D D6
 E3 C0 3D 57 53 9E 08 DB 96 7B 35 61 A3 D5 C2 FB
 FB 6F 14 65 39 02 59 C0 A0 A3 C2 FF 5E 54 16 E2
 D2 EC B7 3B 22 30 96 76 60 A6 52 BE FA C4 B4 F0
 61 F3 08 FA 7D F8 F0 44 A2 1A 70 F4 F2 6B DC 81
 0E 8A E8 FE C5 FF A2 B7 67 64 57 F2 C6 0F B8 BF
 13 19 0A 45 E8 CA 42 C9 62 2C 4C CB B6 04 D8 77
 8B A7 38 A5 9C 0A FF 00 83 9F E0 11 75 CD B3 00
 B3 4D 26 1A E6 29 50 2D 48 89 28 96 29 EF 31 C6
 41 AB B9 4F 12 79 2D 82 B5 88 6A DB BC AA 5D A0
 34 51 5C 12 82 B7 07 1E 37 C0 C3 AC 1A EA 3B 3A
 A3 CC 6F 8C 80 BC CF 31 D7 25 AF B1 70 30 46 F4
 C4 DF C3 AE B0 B6 EA 33 CD 26 A4 2E C0 51 B7 3B
 14 2A 4B FE C0 31 F2 84 DA B0 32 08 3B 66 FF B7
 0D 78 33 32 C9 96 36 CD 24 B2 43 AC 13 39 59 B3
 AB BC 22 1B FC 55 85 1B 54 65 65 CF 43 D4 23 6F
 6F CC EE 7D B5 12 FA 27 35 02 D0 13 46 63 FD CD
 C8 6D A7 D5 04 37 79 A8 52 92 28 A8 5A 24 24 C1
 C8 4C 26 CE FF 7A D5 D5 85 0B 12 ED E7 B9 48 4D
 EA E2 56 A8 B5 88 71 66 99 C4 B8 DF B9 CE E5 CA
 B0 B6 CE FB 09 F3 5C 21 46 32 85 A9 CC 65 3F 03
 E1 28 6D BB D5 E9 B3 CB 04 B1 B3 6E 59 8B AA B1
 D9 FB BA 68 6D F8 AA A4 C8 67 9C 23 E0 5E 0C EC
 62 7B 2A CB 77 C4 1A BE 54 90 B6 C5 A5 A0 6A 80
 2D D8 7A 8B 90 B5 4E 12 F5 80 88 1F CE AD 16 25
 51 1B 1C EB 15 89 1D 62 6B D2 36 7D 78 CF 71 85
 F4 83 77 50 F5 4E 55 99 02 BC 6A 3F FF 54 6C 0B
 36 C6 23 59 EE EA 2C 40 5D D2 18 A5 AF 10 0C 8B
 E7 B2 76 BB 3A 7F A4 D1 10 AE 23 E4 83 38 07 1F
 D2 20 3C 22 FB CF 94 89 0D 41 62 AD DC 91 6C B8
 28 95 CF 6A 2A CD 94 7A 75 94 7D 4C 69 F4 1C 6C
 FA 3A 03 92 52 78 39 75 63 F5 3B 31 1B A4 B0 2F
 52 5C 30 1E ED 11 11 A7 7A 48 7A 3D 22 AB 5E 72
 09 B1 62 6C 66 0F AF 64 58 6E 33 BA D3 03 E6 CB
 0F 26 22 CC 21 78 32 4B A2 7E 62 A0 F7 F1 FB 2D
 B0 A2 9B 81 69 24 8F 85 D4 D6 6D 7F 3D 4B A0 93
 FF AE 0F E8 02 8D DA 7A D6 8C 28 62 4C C9 7D DC
 AF AD C7 25 34 8F D8 00 8C F3 B3 07 E6 EF 3F B8
 5D 23 F9 BF BE 4C 38 8E 4E 94 42 F0 EB 95 97 1E
 92 BC 8E C1 BE 63 8F 70 FD CE CB 9A E5 96 D3 27
 EC D2 B7 B3 6E 05 6A D6 E1 1A F8 C4 4F 64 36 4A
 CA A9 8F 22 45 F9 65 78 AF 4B 78 B8 44 0D 4A BA
 7F 3D A6 32 8F 9F 86 46 0B C8 D5 8B F0 0D B6 8E
 05 1A 01 0A CF 6D 00 D9 1C B0 C5 62 02 42 8A B7
 12 3D 83 A1 3C FC 3C 18 80 49 6D 4B 54 C9 1E 42
 DB 8F AD 02 4B 14 0F 04 14 31 34 93 3D F5 C4 01
 8F 39 4D 42 49 B3 54 05 C4 55 E6 09 45 EA B5 9E
 F7 09 B7 33 7F 7A F1 36 A9 5E AC DB B4 63 7E 5A
 A2 C0 03 96 91 F1 4C E8 D8 ED A0 68 A8 30 76 FC
 6F 9D F6 91 40 33 D7 63 B2 51 8E 95 2B B5 A8 57
 28 AD CB 56 E2 03 B5 2D 58 3A 48 13 45 A3 D8 67
 DD 3F BB F8 49 95 6A 66 92 7D 92 41 25 51 A2 75
 BD 51 BD D0 5A E2 6B 0F 09 69 09 11 AB BB 9B C4
 08 B2 C7 94 2D 27 01 88 83 69 42 07 10 31 AF D2
 D5 B7 62 E5 23 80 99 1A 66 A9 FE 39 29 F5 9C FB
 90 B9 A1 A5 79 8B E3 AC DC 7D 3B 9D 05 5E AE 4F
 86 1D 0A 3D 56 3F 71 94 5C 3E 04 90 97 8A EE 45
 DB 55 77 60 7D E7 CC 70 B3 2E AD 34 2F C7 5E 88
 77 F1 D6 63 A7 FC 2E B4 FF 97 7F 6A BD F2 69 49
 75 E3 5E 6E 1C 39 E4 09 E4 FD 97 65 04 9D 9B 5D
 05 4B 83 D9 B0 BD 34 D0 35 BB 8D 02 65 14 C6 8A
 C4 52 D0 B0 F4 8C 5E C4 74 87 19 43 88 D1 DC 6A
 E6 42 FD 4D 97 4B C6 5F D4 2F 23 4F 3E 7C 1A EC
 53 D8 33 CD 2E 0E 41 66 FE 14 1A F3 E3 64 9A F7
 BA 93 1C 96 D7 53 A6 94 9D 60 05 96 29 A9 65 95
 CD 9B 26 3D 86 A3 C3 64 6C C4 B4 33 88 18 DF 3F
 59 D3 01 A5 84 FA C0 8A DD 99 07 93 CA 91 9B 0F
 82 CA 5B 24 21 FF 1F CD 95 B8 E3 EC F8 61 E3 2E
 AF 86 A6 F9 A9 73 60 E4 17 A2 F0 42 C4 67 F1 4D
 CD 42 C6 07 36 92 67 59 1B D2 8A 8A 63 EE F9 0F
 95 0D EF D6 EC 48 FC 2A 15 29 FB 28 35 D5 7B 6B
 7A BE FF 47 A9 61 9E 00 DE D0 A2 81 86 FC 7D 36
 73 46 22 2B 24 83 2C FC 48 62 F8 65 4C F2 10 48
 BC DA 10 73 F7 93 78 4C 6B 09 23 8E 86 76 31 19
 3F FC 52 81 65 E7 54 86 A6 77 CF 80 05 80 F8 6B
 F9 2D 73 40 FD E1 F0 DD 54 5D 4F 97 2A 35 E0 80
 15 DA D3 BE C5 B6 E2 F1 16 FC AD DD 9C CA 66 06
 9B D0 57 65 AC 57 94 1E 13 90 FC 46 CA 84 0A 5E
 EE C8 6B 14 37 A6 BB 4A E3 4C 48 CF D8 8B 48 73
 60 24 73 0E 7E D2 1B CF 16 AE 4B 4B 6D FD 33 7E
 C8 B8 3C 28 93 AD 5E 94 9A 13 B9 22 12 93 9F 4E
 24 31 48 A4 73 8E A6 4F 41 DC 07 2A 46 A4 4C 50
 53 34 1B D5 B4 E0 49 0C 88 39 9F 42 CD 8D C5 36
 8D E7 8D 6D 0C B0 14 0C C4 3D 78 DE DF E6 C6 10
 A9 7C AF EF 9D 8F 4A 63 24 39 C8 01 F3 0F 4A 52
 6C E2 FB A5 31 85 46 37 E8 49 7A 46 89 FE 53 B4
 5E BE 65 53 F4 F5 26 C0 51 DD 8F F7 C9 59 52 AF
 F6 34 D0 1B 87 1B 24 50 50 25 44 F8 9F 7F 46 01
 14 A0 DA B1 EF BB 6A EA 9B 35 F0 FF AC C3 3D 08
 F1 7B 22 53 10 D4 9E 02 EE 89 4E 85 03 41 12 8E
 18 BA A2 84 26 CE FB 05 19 B1 E5 73 43 70 BF D7
 D8 A9 CB ED 86 DC 79 94 CB 50 3A 9E 46 C8 4E EF
 A3 C1 82 19 24 11 71 9E 2D A4 FA 8A 5E 34 12 08
 33 A5 2F C8 72 5C B9 C1 E1 C1 48 2B E2 3A 5F 3E
 FF A6 91 3C B8 9F 8A E0 B6 F3 AE D9 D8 D5 79 81
 17 9C A8 B5 4E 4C 31 12 59 17 8D B6 B3 DD F8 FF
 CB ED 7F FA 51 04 2A ED 42 7C F3 A0 5A 40 E6 D6
 C5 CD 91 B9 4E 64 CF 85 47 CF 66 20 B5 BE 31 9C
 B8 62 C0 3B 27 82 C1 57 68 40 26 6E BD AD 49 C6
 61 05 D5 2F 01 35 6C EA CC 5F A8 56 BC FB A6 DB
 FA 15 6F 66 A0 E3 81 E7 43 64 45 72 F3 E1 86 C1
 3D A4 61 56 67 EC 07 80 33 BE 5D B4 B6 29 7B 34
 1D 91 6E A9 8E F4 1D 53 4B 4F 0C 05 84 70 6E BD
 70 82 42 18 A5 9A D6 80 83 FA 19 73 BE 9E 8F 27
 1D DB FC 34 AB BA 24 F2 F2 B6 79 F9 D3 C0 9E 1B
 B2 81 F4 2B 01 7F 74 33 5A 01 FF 5D 51 FA 27 1E
 FD 60 03 14 D8 E9 3C DF E4 3E 6F 2D 6E DD 07 CE
 55 05 8B 63 68 23 1F B9 7B 24 82 6C 66 98 0E CA
 C8 22 31 ED F0 C3 B3 5E FC 0C 03 0B 01 B8 A6 6D
 8B D2 41 7A DA 16 24 EA F8 6E 9C 48 A0 6A 57 69
 43 EE F0 68 77 B6 29 9D 4E 4B DD E1 BC 02 33 07
 00 38 CF EE F3 7E C6 B8 A8 34 36 27 E4 58 A5 C4
 AE D2 B7 6F E5 BD 7F 2E 7F 57 DB C9 5B C5 06 E3
 81 11 9D 60 23 5B E5 18 66 8F FC 77 15 68 3B C5
 D2 47 55 2D 64 E7 F7 24 98 5F 08 29 12 36 67 D3
 F2 D7 C4 D3 1B 92 ED CD 39 6B DC 4C 6D 48 20 94
 D4 8D F7 DF 2E D0 7D F8 B7 8A D6 6C 85 AD 62 9A
 ED 32 97 B8 5A D3 8F C4 32 A0 10 90 09 A2 84 5A
 20 4F CC 51 18 2A BD 61 AC F7 F7 8B D2 AA F0 10
 21 10 CD CA 07 5E 25 E3 7B 42 1E DD 84 3E 2B 27
 C9 9D 50 8B 10 60 0F D1 A1 94 AB 3A 8B EA B9 54
 F6 53 C4 5C DA 80 97 99 AA C3 A5 4B D3 74 8B 77
 69 2F E2 39 E9 1C B9 BE 92 6F A1 76 09 12 58 90
 3C 2A D0 68 AA B6 33 DB 50 86 70 FB 7B D5 95 F4
 07 16 53 66 6C F1 84 6F CE 33 2F 72 65 02 D0 FE
 04 B1 70 7A 87 56 F2 95 6D AE B8 F5 AE C6 FB 7C
 CE 5E C1 1F 05 A1 83 5F D2 90 D4 09 CC 46 BC 8B
 D4 D7 B3 50 2E F7 52 94 DC B2 A1 94 6B 50 1D E6
 54 80 F4 90 4F E8 58 92 5D 86 60 BE 79 C2 4C E7
 0C 07 5D 4F 3A 83 A3 B8 CE 19 03 8D BC FF 33 D6
 7E 25 93 42 9F 0F F3 1E 4F EB 8E BB 4E 90 40 03
 D2 89 79 09 9C 12 13 19 4C 69 A1 D1 2C 42 6E 8D
 81 B2 CC 96 25 24 BC B0 92 65 0E 0E FA 02 7D 9A
 6D CB 89 0F EE 11 A0 F8 44 9B CD 49 C2 22 C9 7C
 A9 7F B5 17 18 A8 A7 B5 F4 A0 87 8A 98 3F AA 0F
 C9 F1 6D E4 83 5D CC 6C FA 0D 98 67 1C FE 54 C0
 D2 BF 28 44 5D 27 5D 3E 12 35 D2 05 B8 E5 7A 53
 B4 FF B3 B2 BF 99 B8 59 4B AC 45 E6 74 16 E9 F3
 55 2D 4B 1F 74 84 EC 26 CB 4C E3 90 C5 AA 84 43
 F0 67 EA CF 15 E0 43 CA CD AA A0 B6 CF F7 B7 61
 76 7B 9B 12 D0 D7 77 25 80 35 A5 09 1B F4 0B 16
 D9 60 44 65 26 1B D5 55 C8 F7 A4 D7 CE CD 9C C7
 7B 68 08 89 F1 CB 9D E0 D4 E4 27 3D 76 71 C6 D6
 A3 E5 CB FD 43 FC DB B9 3C F0 3C D4 2E 64 03 77
 A7 C1 70 D4 58 7B DC 36 A6 35 B6 72 E8 47 1C 23
 85 73 81 68 CA 08 B9 4D 43 84 93 92 3C 9B 44 1B
 29 36 DC 9A 6E 01 A1 D1 1F 4C 15 E4 BD 40 76 6C
 F2 89 C2 B1 0B 4A 53 05 95 C2 C8 EC 1A 07 C1 FB
 0E 0D 1E B2 FD 56 44 42 93 B9 59 6F E3 A7 11 63
 32 76 E1 50 B0 A4 B5 F3 25 AC B7 FC D9 04 86 BC
 0F 46 AE 63 5A 2B 2D CE D0 67 7A 62 DA 8C 43 3F
 CD 3E A8 BF 1C 35 3B 12 2F 9D 90 3C A7 00 C2 22
 CE 0B 8E C9 28 28 D4 92 61 2F 0E 08 DA 75 02 9E
 8C 2A 07 A0 FC DE F3 B6 85 0B 30 F1 F7 95 4E 46
 24 D3 B8 8C 85 1B 18 B9 CE D7 C9 27 45 8C 3D D6
 9B 84 61 F8 8C 05 74 1C FD E3 BC AA AE DB B8 40
 10 94 F9 06 B7 24 40 DF 6D 74 77 21 3A DE A3 A0
 D4 F3 8D 70 F8 21 F1 5A C2 C8 54 2C CC 5F 7D 9E
 85 CC 84 8B 36 51 14 A1 87 2F 95 82 6B A4 C8 9C
 DE 94 A0 08 52 27 BC 48 74 1C DB 31 8F E4 E4 74
 BB F4 85 92 DC 53 AA A8 9A 89 20 0D DA 84 3B 57
 EE 9A 6B 06 17 C1 7E A6 67 79 E0 40 1A 93 82 D8
 D0 C5 6F 50 40 6C DD CD 0A DD AB 10 48 E7 C1 F6
 F0 08 1A 45 30 F7 B8 68 94 6F 40 A5 5F 38 33 1A
 7F 67 F2 44 10 8C 82 D1 23 F2 8B 46 95 60 43 29
 0D 02 63 F0 24 E1 5A A6 A5 A8 DE C7 34 95 3E 52
 4A AB F4 C6 7E 75 28 93 AE F8 9B A8 A8 5B 0C 47
 CA 6A CB 4F E1 D6 02 F2 EE 66 5B AC 54 50 1E 8A
 A9 ED CE 73 87 0E 86 40 EE 54 B9 0E B3 C3 D9 11
 76 B4 ED C7 FA 3E C2 07 10 2E 8A CC E0 6C 8E 71
 AF 49 4D A8 53 48 98 16 B3 AE AB EC 02 65 0C 27
 8C BB 3E B0 F8 B7 31 32 F0 59 A9 5C B5 50 76 40
 FC 81 02 63 3B 9F 2D E1 68 50 FD A6 86 3D 6D 49
 C3 33 F1 2D 65 65 E4 76 A4 D7 7C 0B 20 45 F2 08
 C9 9C 09 89 18 A7 87 D4 51 99 63 F4 38 2E 58 F7
 0E 6E B4 05 16 7C E5 9D 0A A0 CD 54 B3 E7 33 E1
 0E C8 73 EF F1 E3 73 B4 75 14 23 89 99 0D 37 F9
 B9 81 A7 F5 65 CA 37 76 EA C5 5E 3A 53 5A 7E 9A
 FD FB BC 64 6E 25 67 B8 59 98 C5 21 43 E4 3A AA
 02 61 C1 29 A0 2E 5B 7B 36 A5 89 A9 7C 7C B8 8F
 5A 66 35 6F B5 16 27 D3 62 F6 AC 50 AD CA 17 28
 A6 96 27 61 C2 B6 05 1C 08 7B 26 B5 E8 FD D8 5B
 2B C6 63 12 1A BC 2C AA 59 DE CA 3D 4C 6C EA 82
 AF 20 24 67 27 F2 47 0B 57 C1 5A D3 E5 55 74 86
 52 14 C7 67 DD B6 E0 85 B2 99 3D FE DC 79 08 96
 AB D1 5B 6B 37 24 AC 12 EB 6D D7 57 18 31 BF 0C
 12 AF D3 7B D5 22 A9 1B CB 72 68 E6 30 59 C5 4D
 F9 78 8A F0 57 14 77 7E F5 AA B3 9E C3 7C 3B A0
 6F 6C C3 80 73 49 13 B1 F3 16 24 0A F6 08 FB D1
 98 0C 8D B3 DB 73 94 50 C1 86 87 2A DE B4 53 21
 E2 6A E0 7C A6 B3 8F EF B8 EC 7F C5 89 36 62 0A
 11 CB EC DD 4F 3B 15 39 81 28 F1 2F BF E6 73 C0
 CC 27 3E 17 82 A1 47 E7 FC 30 FF 91 45 4E 20 23
 70 B3 41 63 8A 17 80 65 30 28 A6 29 29 03 E0 C2
 2D 4B 95 A2 A3 10 75 72 C4 89 4E 98 F5 A9 A5 64
 16 F2 99 30 00 58 FE 1B A2 B6 0A 77 27 75 AB AB
 8F 69 53 14 DA E5 25 E7 0B BE 29 50 34 0B EE 67
 73 A6 A5 B5 0F 41 48 4E A6 BC 81 63 67 05 E3 61
 E4 2A FB 2B BA A8 A8 B2 3E E2 65 6A C3 9E 96 68
 F9 1F 8B EA F5 9F 96 74 42 37 88 87 64 6D 7D 27
 4C 83 F6 D8 45 E1 42 7C 8F 3B F9 37 AF EF 2D 47
 97 F5 78 B7 10 E5 F0 90 3A 94 3C 1F 4D C6 75 D1
 C5 AC 1A DA A7 97 1F B3 62 52 72 B3 60 6F 73 B4
 CE 94 3B E5 54 C7 EB 20 76 56 0F A7 EA B0 52 04
 B3 1C 65 F7 50 BB 53 4E 8E EA 3A 98 32 FE 21 D6
 74 0B C5 A7 42 8A FC 67 A2 64 2A 59 82 54 C8 D6
 08 3E C5 70 B9 CB 23 75 D6 7F 47 A8 80 30 72 63
 C1 C5 39 63 BE EC 71 7C 8E AB 33 8E 0D 87 EB 9A
 66 CC 40 F6 39 3A 8F 3A 70 33 BF 41 67 28 F9 F2
 11 3F C1 0C 69 13 A8 15 15 95 F4 AD E8 06 71 85
 AE 88 E6 61 71 7D A6 3A 48 5E FC 36 07 31 30 88
 CD 9B C7 BD 00 00 0B 95 65 EF C8 27 3D A8 99 FD
 26 BA EE 09 AA C3 92 9C 27 B0 D3 C3 70 8F F8 64
 E2 52 4B A6 B0 6B 0B 58 CF F2 89 6A CE 9B 1B 7C
 73 B7 57 C2 FC 2E 7C F8 80 9B 35 32 CC 17 A9 F1
 0A 81 42 1D 4A 6E 9B 54 A5 58 FD 67 9D 20 80 92
 03 08 F8 D0 28 35 1F DD 30 BB 74 D6 34 4C D6 1C
 18 6E 90 F0 E7 C4 DA D0 31 06 13 15 81 02 A0 8F
 23 9F 08 67 BA 65 59 4B BE 93 6B B4 E3 81 20 12
 D1 B4 1A 8F 2B 12 01 00 BB B2 9F A9 7C A4 5A 60
 3F 19 24 51 17 61 0D 07 F8 2A FF 6E B7 DC A2 75
 C4 C7 8F A8 39 4A DD E0 4A C4 74 74 AE E1 9F 68
 92 93 08 28 42 FE 73 B9 4E C0 88 EB 33 D8 B9 30
 B0 A8 D9 4C 79 91 5F FF 16 05 41 52 DF 9E A6 81
 B3 E7 2C 58 BB A3 B1 36 E3 3C 89 9A C8 07 12 2F
 8C 29 60 0F 73 FE 41 E4 FC 70 D5 D0 32 89 89 FE
 00 B3 BC 43 EC F9 93 4B 2A 2B 1F 6E 4E B0 FC 90
 1B F2 4F 7A 12 7B 37 6E 2B 4C 46 01 F0 20 F2 B5
 4C CD FF 22 59 04 EE 48 E0 F3 8C 1F 1E A5 47 2B
 8E D0 5B 1E B1 DC B3 8C DF DB 5A 3F 15 C0 31 64
 0C 88 D1 F5 54 25 BC 70 6E BF 05 97 CA 1B 75 0D
 2A F6 39 48 B9 EB 38 5E D1 40 65 E4 5F 75 93 E8
 E5 8D 96 59 C9 B1 F0 E5 B8 C2 E8 F0 B0 46 B7 AD
 15 53 B8 83 67 77 1F 25 9F C7 AC 1E 4E 12 8B F9
 85 7E 73 11 BC CC 9C 4C B0 C6 42 D4 54 38 67 00
 8F 05 FA A9 5F 89 E4 AF 96 E7 4C 2A 28 8B 05 5B
 4D B7 D1 58 DD 5E 9E 76 37 CA 8B D4 84 0A 45 1E
 55 7D 91 CD 2D AE 01 9A 50 8D 3A E2 FF 1D C5 3D
 F1 51 5E FE 74 9A EB 44 58 36 42 4D 46 C8 C1 B0
 CB 53 1D B8 60 63 54 CC C7 26 E3 B5 38 6A 9D CB
 3D CB E8 92 1E B7 C0 6C 84 FE 6B 76 6F 4E 43 C3
 7A 11 AC 7E F2 C0 79 A0 9D C2 08 24 1F 3B A1 D3
 C6 0B FE 73 D6 6F ED 15 7D 5F 4E 83 BD 92 F5 FE
 89 C7 99 5A 68 FA 74 C4 23 6D 83 C7 D4 EA 27 07
 5C D7 EA C8 A9 F9 29 08 FB AB 10 95 2B FD AE AC
 BC 37 1B 0A 4B BD C7 58 93 0C BE BF 99 C9 AA 1E
 C1 F8 0A 64 9C 14 19 30 8D 66 71 BF 90 B7 3B 5D
 9B 36 33 A4 73 8B 11 9B ED 19 52 96 CD 6C B1 03
 2D CA 90 7D 0B 4D C5 32 C5 68 69 31 EB B8 65 27
 C5 65 D4 88 5A 3E D8 07 AB 4B 6E 0B 07 BE 55 B4
 F7 C3 00 0A EC 92 BC 24 A7 B3 F9 E3 D7 41 08 E9
 E9 C3 6B 6F 27 08 52 7A 44 7B 98 8D 2F 20 59 65
 8E F1 6F 8D 1C 27 DC 1F 45 BB 18 CE 0A BF 6C 4A
 A8 12 AA EA D3 36 21 74 64 9E 95 DB 6A 50 71 CF
 9E 55 21 D0 67 ED AF 16 34 EB 63 62 1E AA 9B 61
 7D F2 3A BB 10 99 AA DA AB A9 3C B3 C6 B4 E9 7C
 91 6D 7C 9C 68 0B BB 80 A0 7B 52 EB 8F D4 B5 29
 16 38 B6 2A 5B 87 52 F8 B4 00 A8 03 8B 38 7B 1F
 4D 0F 9D 30 71 DF 03 9B BE 63 B3 6E 78 BE D7 96
 5A A6 1D C5 0E 59 C7 86 14 32 B7 41 BF AC 38 F1
 92 22 4E EF C8 15 B2 AF 7A BC D5 3D 99 ED B8 2F
 64 F7 54 93 28 34 CA 9C 66 99 DF CE 2E FF 33 39
 99 4F 1D 63 D6 1D 7A 5B 15 44 BE 92 5E 76 8B 59
 B7 2B 23 A9 AB 60 05 50 F8 A8 D6 BE E9 AC 44 38
 4B 15 4E 63 81 02 C6 A7 C0 F6 A4 12 B2 C8 39 E1
 1A 3D 3D 77 FD 84 C7 AD 02 42 36 B4 2A 6B 5F 10
 B3 C1 9D 24 FF AD D0 92 01 59 BB 65 CB 9B 64 19
 FA D5 39 CD 2B E9 B3 D1 58 9F 09 04 0E 57 27 BD
 64 12 73 B5 79 66 D8 14 0E 2C 07 D6 CA 64 8A 71
 77 A9 20 00 A7 8F 2D 87 CA 81 E4 4B F0 CC C7 53
 DF D8 A0 9B 73 22 CE 9D 8C D8 78 B6 27 CD BF 3E
 5F B1 A4 05 C0 07 24 F0 F5 8D C9 75 CE 46 7E B3
 06 25 20 E4 B7 C2 05 B2 AB 5D B9 A0 3A D2 62 B3
 77 E8 FD 7B 33 2E 0D DE 3A FE 9A F3 CF 8F 71 FE
 1B 7E 62 B4 47 56 AF 0F 0F 4C 0A F8 01 28 1C 13
 2E B3 7C 95 A1 18 8F F2 D8 4D B3 9A 9A 12 F8 68
 9E 5C 6B 4B 43 81 6B B5 F2 37 12 0A DF BD 57 BB
 A5 84 68 49 7E 38 35 D4 01 AF B7 24 AF CB D6 B6
 5C A5 E6 35 FC 44 AD 15 83 B4 90 71 FC BD 7A 42
 18 C9 A9 29 DA D9 5B 19 47 F5 F8 97 50 6A 19 DE
 06 77 E9 A1 20 D0 1A 4F 3F 7D CD 3B FF 84 F8 4D
 51 22 87 FB 06 DF 24 64 8E 20 61 6F 20 67 D1 CF
 98 EB E1 6B 69 58 C5 E7 7B 8A 52 03 DE 4B 8E FC
 7E DF 7F 01 E6 09 A1 A4 48 44 EA CB C4 CF D0 A0
 BB C9 80 12 35 2A 12 65 B7 9B F7 2B AD 3B C5 86
 7A C0 A7 0B 96 9D 47 23 A4 21 FE 93 A0 15 73 17
 B0 8E A9 5A 5A 5D C5 F0 48 0F 38 30 AC EC 28 FE
 85 4F AB A0 F9 14 06 EC E0 B2 48 60 E3 59 53 9F
 BD BB D8 70 F7 00 C0 64 AE C6 25 DF 69 64 E4 05
 8C DB A5 07 6E D1 7D 27 12 95 BD BD E9 A7 1E BC
 C8 A6 5B 9B 0D 7C 7A 94 01 E8 6F 6D 9C C7 5F 2F
 43 72 34 76 15 BA DE CA 76 B4 8F 52 2E AF 42 EE
 FF 35 D6 5B B4 2C E4 5D 3F 3C DF 0A 0F E1 D8 7E
 BC 62 EF 76 84 30 D3 C3 20 1D 27 E2 C1 8E CE E1
 BE C1 ED 4C F5 35 CB 3A 14 2D 96 3D E7 92 BA D2
 0D 9B A1 D7 78 7D AA F0 12 93 E8 F3 95 EE 1B B3
 F8 C5 F8 42 5D A3 83 C5 C1 6D 74 F7 08 CA ED 5B
 17 FD 99 2C 81 7A 60 0D 40 A4 42 2D FD 9F 78 7B
 C9 68 A2 62 C1 44 A8 4B 14 BD 3B 5C CA 9A D9 3E
 AA 39 7B D6 1B 3E B6 BE 1B 2B CC 2B 6D 5F EA EB
 D5 2E 20 C1 AB 27 97 BB CF 4D D7 CB 52 7C 24 98
 90 DD CA BF 87 3E EE 89 62 A6 04 80 C8 42 4B 92
 4D 44 58 CD 3B 34 D0 4F 8F 48 8F 02 26 74 83 DC
 B9 B5 18 CE AA 77 6E 17 64 76 B9 AB 42 9C 2F 88
 6E 06 DA 51 FD B8 57 D5 32 4F 9C 6E 84 43 F8 D6
 DF F6 B1 61 F3 F0 8E C0 B7 E1 AB A7 0D 55 CA 20
 B3 4A 5E A9 AC 82 3F A1 CF 5A 81 91 EF 2D 1F 8F
 29 BF DD B6 4B D5 CA D9 60 98 3E 13 E8 27 B4 93
 16 67 00 5F FC 6C D0 5A A4 B2 6E 4D 8E B5 46 3C
 37 8C FE F7 75 CB 6B 91 AE 01 7C B9 40 E6 D6 6F
 8C 5E 1D E8 53 44 AA 25 4B A5 B0 67 9E A4 74 4C
 C5 AE 55 43 1F F2 A9 E3 9D 4E BF 43 1F A5 A3 AF
 64 40 23 E0 36 01 D0 F2 70 BC 76 C0 87 71 77 48
 AE 6C E4 5E 93 58 A8 C7 21 EE 73 A5 27 1B B5 50
 CF FF 45 73 9D 24 F8 D9 0A 5E 43 DF 30 E6 EC EF
 3B A5 5E 55 77 3B 1E 37 92 96 DE B2 3B 72 13 CD
 0E 12 28 E2 EE CD F3 51 18 F9 AD 6F D6 93 00 E7
 92 B3 21 9D 15 90 7C 0B F9 FC 4C 23 9A 07 AD DD
 28 3E AD B2 EC 7B 41 01 E6 04 69 76 B4 DB FC 29
 20 1E C5 A3 24 53 01 EF 09 2F 25 61 4B FB 35 37
 2F 4B 24 EC EE 6E 0D F2 AC 66 16 76 B4 CD F5 59
 55 21 E8 55 10 C0 AA AF C8 13 F4 C7 60 E5 C1 6D
 2C 70 C5 06 8F 0D 20 25 DD 78 D4 17 81 DB A3 40
 1B 9C 71 EE C6 47 3F 60 D2 DA 77 13 45 45 59 EA
 CA AB 84 DA 4D 93 22 29 8D 09 AD E9 19 D6 78 01
 8C 9B B1 9D CA F7 76 E8 D6 B5 5A 79 85 E3 5C EF
 E4 36 B9 70 9F E9 E3 94 89 80 A7 16 7C E9 F5 39
 C7 46 C5 D4 E4 83 26 7E A5 50 FD 4E 57 FA BB 22
 64 75 ED A6 BC 11 D0 54 D7 86 B6 16 C1 ED 29 05
 FB 11 BD 7C 1D C9 20 25 70 80 90 AF C0 E1 D2 0D
 B0 3B 18 C2 A7 E8 EA 67 EB 6D 94 77 78 66 96 19
 EC 36 88 35 D3 E9 01 DC 8D 00 83 E8 84 29 F5 90
 F0 74 FD 1E 7E A4 AB C6 DF 41 A5 E9 AD 8A F2 6F
 D0 16 38 BE BC 3E 53 68 BF C8 23 45 60 D4 DE 4A
 03 B0 F0 DC 86 0A E5 56 CE 22 D5 9A C1 09 71 BC
 53 7B 67 8D B1 5C 51 6C 8C 1A ED 46 AD 82 0C F7
 67 10 B4 D1 CD D0 23 6A C0 AC D3 93 FD 5E 7F 5E
 60 22 32 3C C8 D4 B1 85 65 87 AC DE 34 10 74 98
 29 CC 6E F2 B7 0B EA 24 13 B8 80 30 8F 77 4B 84
 E3 D8 03 09 24 9B F0 DB 36 2C F9 AF B9 4F DC 4D
 4D 9D F3 CA 29 37 67 EA 14 2C 27 6E 2A C1 E2 79
 4B 87 0A 1C 10 62 B7 4E D1 7E 26 90 FB 9C 13 DD
 7E 7A DA 39 1C B4 CA A9 73 5E 7E 30 F9 82 7E 0A
 96 8C 05 FE 19 6A 2F F4 9E 46 01 66 6A DC 6D D6
 C0 C3 D4 D1 69 8C 01 F9 62 80 FB 8A AC 9A 76 75
 BD DC AE 3B 5A 8E 4F DC BD 10 B8 66 6B E5 84 8F
 72 5A E8 78 C0 36 48 84 78 AB BC AA 2F 35 F2 A8
 7F 5C AD 05 BF 99 ED C6 74 BA 01 E4 46 DE 12 F9
 3B 67 21 88 6D AF 0C D5 83 F2 06 0F FA 90 82 76
 F7 EB 31 21 77 F8 7C CE A0 AA 57 24 AA F6 E7 E7
 A1 70 BE 60 00 24 0C 97 BF 9D DD 86 ED F9 5D EA
 7B 84 7A D6 70 2C 20 64 83 13 18 85 1A 68 7D 94
 50 EE 9D 9A E1 7E 71 73 AD 37 3F AA 61 E3 24 8F
 FA 10 BA 40 39 C0 42 BB 54 6B 47 B6 B5 FC 50 DB
 84 8D 0B 42 7C 0F 81 59 36 AB FE 4D B9 49 83 C9
 A4 10 9D 72 CD AB 5B 9E 42 77 F7 7A 0C CB E6 9C
 86 5A 2A EA 2A 99 3F AF E7 87 32 97 7D 69 C7 35
 B5 77 D5 23 EF 3B 0C 44 D0 83 46 E9 3D 85 9B DA
 5C 4D A2 BF AD 57 4C 29 BC 13 73 C0 77 BF 12 AF
 98 6F 6E 93 99 98 61 21 05 95 CB 5F D1 D1 67 AB
 D9 D7 1C B2 29 E8 BE 3F DA AF DF 76 13 26 E6 3A
 65 0D AE D1 99 F4 F2 82 8B 98 0A 58 40 9F A8 02
 20 DD C9 F9 16 1A A0 47 DA E1 01 6B B4 46 50 96
 48 1C 36 82 C1 39 13 F6 3D E5 A5 44 6F EC 8E 66
 EB 62 64 DF DA D4 78 F4 C1 FC 25 BE A9 04 44 91
 25 32 7C C2 7F CF D0 36 B7 78 BB 45 C0 79 6D BB
 80 58 7C 2E 12 CE 60 F9 B4 BD 18 C4 E2 68 8C 5E
 BA 57 C3 2F A4 41 CA 87 2C 57 BC C5 9C B3 37 78
 A6 59 56 BF 17 7C CD E8 13 67 8A CB 22 9A D9 13
 92 34 7D 19 79 35 19 15 15 B4 7A 89 AC C1 E2 6C
 CA 92 0F 78 72 B9 B5 AB EC 6F 77 89 A0 79 30 69
 35 B1 5C E3 CE 57 0D 6A DF 3C BC 8C D6 DD FF 16
 41 27 96 4B 61 85 16 F6 10 CB 38 F6 D0 9C 11 21
 84 81 54 3E A7 09 A3 6A 9D A6 AE 6E C5 D0 55 FE
 51 5F 00 67 25 B2 B7 C2 45 AF 6C EC 99 7C B2 FA
 BB 38 BE 3D E0 7D B3 AA 94 51 84 DE 5C 27 90 69
 FB 0D EA F3 E5 14 EC 32 86 8C 8D C6 15 6E DE 49
 A0 60 C4 D4 04 CF 8F 28 B1 A0 98 B1 26 E9 6F 76
 49 B3 77 06 D9 07 CC FF EC C5 C6 89 55 F4 80 5E
 23 3D AE 77 D1 ED EA A8 51 D4 6E 6F 59 2F 02 1B
 04 00 B4 B7 48 C4 47 92 FF B1 24 54 9B 9F C0 A8
 C1 62 8D 86 02 B1 ED CF B4 E3 D8 56 93 13 BA 68
 83 D3 1B C5 5F 06 32 9E AD DE BE 37 13 30 45 47
 94 6E BD 03 79 76 46 F8 27 B6 06 8E 44 CF 92 44
 1D 1B 93 11 DA 85 B2 AC 84 D5 76 D1 A0 BA F7 F8
 2F EF BE C8 7A 58 8E 95 19 AB F2 87 ED 6D 84 CF
 A3 D8 02 5B A9 DC F9 A7 74 FB EB 3B 8A 2F 24 6F
 B7 EE FA 14 53 FF 36 51 3C E2 86 9B 5A 66 DD 27
 DA 75 A2 06 3F 37 BE D0 63 43 96 B0 2E 3E 4C 2E
 BD 21 A1 AA 60 16 C2 93 69 65 E2 BD DE 09 C5 10
 D8 4F C9 E8 32 54 A3 86 FD 1A F1 D9 2B 8C F1 B7
 97 85 BB F9 DF AE EB DE 16 CA 0B D6 5E 40 42 A3
 97 61 5F BA 37 C1 0C 2A C6 39 CD 5E 7F 71 07 8D
 BE 1A 51 51 D5 E0 87 8D A0 18 F2 75 3F 31 59 23
 42 8F CA D7 D4 31 74 3E 5F E8 65 84 EC 42 89 E3
 AD 3D BC 9F 69 96 8E D5 AF 83 88 A8 67 6E 15 17
 97 5D 70 9C B9 D4 4E E3 8C 23 B6 F9 5E C4 EB BA
 E9 E5 E5 0A D2 69 D5 59 BB B6 00 F3 AF AB 06 40
 CB 13 08 ED 11 08 CF 05 F6 3E EA 73 1F 04 31 56
 2C 0F EA 55 E5 B0 12 5D 06 28 05 D3 BC 09 1A B6
 AA 3D 56 5F 51 F5 8E 85 F0 FD 12 CF 84 27 32 10
 C9 9F 18 4C 09 F1 F5 EC 83 3B AD 66 A2 AD E2 FF
 8B C0 32 B6 0D E1 66 84 7D 45 F3 75 06 9D 54 05
 F0 5A 2A 33 7E C6 41 C2 ED 71 82 3C FD 78 78 E4
 02 0B D2 D4 4B 56 25 57 B6 67 39 1F 0E 8C 5C 90
 42 B3 88 DB 61 F2 D5 59 D8 0F 87 6C 38 C1 EC A9
 A0 D2 A4 DD 30 31 18 98 5D 61 74 A4 F1 11 E1 34
 40 BE 9B 28 E2 CE 2E DF 7C 8C 0B 4A 17 F2 A3 01
 4C AF B3 AA 0D 26 95 3A 1C 5F D4 D2 E3 5F E1 77
 E3 39 64 8D 22 31 26 DD A9 93 19 32 63 27 BE 65
 E8 60 86 8F BB EC B6 4D CD 40 8B E9 0B C1 46 D8
 47 46 D9 DC F9 38 1C 70 25 CA AA D5 4A FA 88 2E
 EE F9 A6 E3 07 1E 78 A0 3C 60 34 5D F1 FF C9 33
 44 0F 59 5F F9 36 69 F2 DD FC F8 A0 C1 D2 BF 1D
 2B 8F EB BC 84 33 71 BC 66 F1 A0 10 F5 2A FC E3
 4B 23 4B 76 38 D0 FB C0 02 0C D4 96 35 4C 12 B2
 16 7C 8B 13 16 48 11 F0 A8 D0 AD 49 DF 03 FE D4
 3B F2 C5 92 2C B3 BD 80 BD 26 E0 E5 4A 90 30 7D
 85 91 7D 79 08 77 AA 20 0A F3 81 24 A7 AD 17 15
 90 DF 51 21 C6 72 D2 A3 80 5A 04 C5 A0 77 6D 25
 5B 91 A4 51 3D 5F 38 58 53 88 D4 77 1D 58 1D B0
 68 12 97 19 69 11 4C CE A2 B0 4B 90 C2 4B 93 68
 A3 80 95 C5 B0 12 83 63 C7 6C 65 76 2E 41 E5 EE
 E4 FB 0A 4F 20 4D DC 7B A4 0E 97 79 10 B1 E3 B4
 4A 81 7B DF 55 A7 BA 19 41 A8 7B 55 11 BA 2D D5
 FD 64 5E 93 BA 63 1A E2 16 8F CC BD 22 9E 5B D8
 07 67 1F 29 06 1F 66 1E 67 48 6D 8B 45 90 7C 59
 E2 BF 0D E4 8E 1E 21 86 77 57 FE 87 B9 52 9F 03
 33 40 B0 66 1C 67 C4 3B BE BE 80 AF B9 6A B6 25
 85 A3 C4 5C 9B 4A 23 17 D5 94 AA BE FB 17 E7 DA
 F6 AD 25 A9 07 5F AE 39 90 06 D0 06 AC 95 E4 F1
 60 D3 F9 4A A6 8B D0 07 B7 90 AF 2D 90 46 B5 FD
 81 FB 0D DB 1D 19 A0 F0 C2 64 DA A8 93 08 8B 34
 A6 1E 00 6A 5A 6E D4 1A 31 C5 78 91 3C 0B 43 28
 86 10 80 E0 3F AA 13 BB EC 2E 21 3C 18 EF EB 74
 8A 53 8B 19 33 3A 5F FF E3 96 FA 66 EB 6A A3 4E
 04 8E 08 E1 EA AB 95 26 94 A5 91 F3 03 42 6B 28
 83 2D C5 7B F7 05 51 72 E5 C6 B3 E6 53 C5 24 1F
 89 19 78 45 F9 39 CE DB 5F BE 88 FA BD DD 33 F9
 93 93 F8 2D E3 B6 B1 53 6A 67 1E ED 1A A8 14 29
 67 7C C2 4C 98 C0 59 72 71 D8 35 70 64 45 59 30
 DA B2 06 9D 63 4E 42 FC F7 66 22 68 1F FB D3 58
 B6 3D 4C DA 93 AF 05 0F 9F D7 7B 97 70 FD D6 7B
 B2 65 DC 24 4F 6B 70 F4 72 85 F4 7E EB F6 EA DD
 93 D8 CA 62 26 08 93 BF 56 68 21 8A E5 6B 9C F2
 9A 2C 14 23 F7 AB D5 9F 95 53 1A 92 D5 F4 37 2F
 E9 78 C4 70 95 38 DA 65 26 FB 7E 97 6A 1C 5D CE
 D1 6A AB 59 25 C7 A4 62 2E 64 70 27 02 DC DE 0B
 C1 C2 EF C1 35 67 5A F6 E4 D3 13 F0 F6 EC 04 02
 C1 C1 8C 99 00 89 02 B7 92 B6 60 BA D1 D4 78 2A
 81 7E 65 45 DF D9 7B 27 7E B6 23 2D DE 7F 91 EF
 D9 4C 15 E1 5C DD 79 BE 43 37 73 C1 BA 05 B8 B3
 72 23 60 11 79 81 9A DB 89 EB B6 F0 99 A0 D0 08
 34 A8 45 FA BB 43 DD 8B 64 EA 18 D3 83 90 5D A0
 2B 75 FC 87 C2 31 AD DB 7D 06 F2 C2 C4 39 6D 1C
 89 C2 81 CD 67 3A 22 1F AC E6 C7 E9 47 11 7C 9F
 44 B2 CE F7 59 D6 87 DC 79 00 11 24 44 A3 7B F2
 18 96 02 C1 2D A0 92 17 65 EA 00 F5 6C 02 9A 8F
 52 10 C9 BD C3 65 78 83 E1 A9 21 06 DD BE AB E4
 1E 70 AC A7 F9 80 D4 77 92 D5 F9 D4 3C A2 E3 FC
 27 13 C6 5E E2 3F D8 EB DE F6 0E AD CD FC E9 5B
 20 7B A5 60 F1 23 07 A7 B8 CA 3C F4 FE 7A 8C ED
 C7 B1 3B DA 24 A4 46 61 63 38 87 E8 B0 52 BD E2
 37 3F 55 F7 45 3F 35 88 74 DC EE 03 28 9A 26 11
 4D 0D 84 ED C3 95 6D 7E 1F 4B 8B 76 9A 8C 4A 32
 0A CA 82 60 03 4F DC DA B2 D5 24 94 3F 78 82 F4
 D5 C2 80 96 2F 95 6B 46 1A E8 CB A4 D8 0A 62 49
 BE 1A 4C 33 FE 21 30 AD 97 2B BB F7 6C D0 C8 98
 2D 97 04 7A 0F 4D 77 07 01 B4 70 CF 81 C2 63 38
 61 C4 8C 0D 05 4B B9 75 C4 B6 79 29 F2 5C 2D 6D
 C0 45 99 02 DA 9C 85 86 27 5E E9 B1 ED C4 E4 0E
 00 3D 36 46 79 CE F2 64 53 E0 F2 EF 9F 38 72 16
 12 C4 B9 3A 07 7E 8D 15 67 76 D3 FE 75 E2 47 97
 69 9B ED 3A 00 4C CE 1D 82 FD B4 05 06 80 4C E3
 B2 F1 D0 19 A6 8F 77 1D CA 5B 73 26 20 96 37 E3
 54 09 FA 22 70 13 EB E9 5C 24 F2 6A 7C 82 CB 33
 66 B1 9C ED C0 65 9D 08 89 9F 1C E3 B0 0E D2 C8
 73 71 E9 36 9E 6A FC 84 BD FC 74 10 D7 0F B9 BE
 3D 80 EE 8D 59 E9 D9 60 58 40 79 7A 22 CA 39 41
 51 0E 33 F8 54 6E F9 F9 65 84 F9 21 27 7D F3 8E
 DE 49 90 0A 5A 42 0D AA D0 5D 38 70 3E 65 DB 3D
 15 78 EF AE FB A1 67 64 92 79 1E 52 B9 D8 2B 7D
 61 A4 DA 7C 6B FB 8E D3 13 7A FF 12 0B 52 6F 98
 2D 8A DC 1D 1C 23 B9 E4 30 6A 14 80 08 EE 62 35
 82 73 1F 13 3D D6 EC B1 46 FE 5E 5C D9 9E 10 E9
 83 19 28 EB DC 8A D0 6A F0 3A E0 31 9E 14 CA 07
 79 E4 5D DC C6 93 00 7C EC 9E E0 86 11 A1 6C CB
 68 64 75 B6 8C 3D 86 D8 49 7C FC AA BB 4A AB C7
 E1 67 18 3C 1E 44 70 6B B8 DE BB 42 FE FC EA D3
 8B A6 61 4F 09 F6 12 F3 80 88 46 C3 A0 4E 46 1B
 92 A3 07 28 BC A0 AA 4D C2 22 29 5C 19 40 96 0B
 B1 1C CA 7B 1B 90 C3 52 9F 80 0D 2B 49 37 76 29
 1D 1A 88 AE 15 84 07 25 41 DC C3 A7 AB 7A 5B D8
 8F B6 4A 03 61 9A 1E B3 D8 7A 64 8C B5 13 BA 35
 A6 57 FB 87 3A 67 4D D0 BC 7A 20 D3 B9 F2 81 89
 30 66 9C DF 2C 9B E9 C2 D6 EF 48 8A EA 8B 96 29
 01 4F A2 68 B9 80 AC C3 63 A9 4D 70 C3 68 74 B1
 2B 6A 99 62 56 91 04 B3 64 E4 8A 8C D2 30 77 53
 52 6A 25 2E 5E D5 95 6D 6C 93 CD 04 B5 92 20 84
 47 D3 6D 9C 5A 24 B7 93 A9 89 96 67 7D 0D DA 66
 99 48 D2 DE 08 D5 A5 8E E7 BE 9D 59 B8 85 B8 C5
 FE 38 10 86 26 8E D7 D7 05 CC DE 6B 88 DF 80 92
 7E 1D 4B 76 A6 4F 2A 2B 80 15 F9 2F D8 61 BB FF
 96 BA 09 D8 C9 0D 5E 55 E0 FA A2 44 58 EB 97 11
 AD 79 C0 C3 66 44 73 90 32 88 99 78 E4 5F B1 68
 B8 F8 13 BD 85 30 9F 0C F5 21 F3 F0 F8 E2 50 CE
 30 71 8F CE E1 F3 A4 30 1A EA 69 40 A0 7A 37 47
 BA 6E 4C 97 21 26 57 89 81 76 17 5F D6 48 76 4E
 72 75 A8 C8 63 C8 2D 08 90 73 18 E9 BB 7F 71 4E
 DE FA F7 24 FE F1 71 85 02 76 BE A8 C6 C1 E4 E4
 4F 11 CA E7 1F D4 E9 81 80 DD 97 40 A0 2A E8 06
 7A 67 7E B0 FD A3 05 91 BA FE 30 41 EE 34 CB 8E
 42 20 B6 1B 33 52 46 BC F1 1F B3 09 84 2C 8D EC
 9A CF 74 85 D3 1E 18 00 46 30 F0 AF 4F F1 C8 D8
 2B 88 3C 3F 78 1F 41 86 F2 D4 A0 AF A4 78 1F CA
 4E 09 6B 2D 96 53 D2 40 40 01 44 43 65 F4 D0 48
 39 07 92 62 53 59 9F 62 B2 14 85 48 C6 D5 E5 77
 DD AA 65 52 8A 4B 2A 21 EE 06 D0 58 B5 1A C6 68
 BF 16 8C AD 5A EB 73 E2 7C C2 13 77 0C 28 10 9C
 27 27 0A DB 3F 6A 65 6E C3 55 A2 F3 91 54 2F 96
 48 3F 7C 35 A9 74 2D 33 A5 05 13 85 8E E9 09 3A
 BC 0E 13 C2 65 7B 0F 1E 5C A8 AD 71 35 8A 51 59
 18 C8 67 C7 65 ED 9B 21 F9 0E 3B A3 82 CA 43 30
 48 42 59 C0 0A ED 8E EC 96 21 BE 80 68 F9 D2 EB
 31 63 F7 43 1A 7E C5 B5 D8 DC 29 0A 49 28 F6 0E
 E0 FB 65 D5 32 D0 66 0A A6 33 F2 90 7E 2D 6F A3
 C6 73 5A 67 A2 E6 AD EA 95 5E 49 D3 97 6B C4 B7
 26 B5 70 E4 4F 11 F0 B7 6D 4A CD 33 84 C8 CA 6B
 92 5A 67 AA DF 6C 05 A3 A5 87 A8 47 28 B8 EB BD
 1B 23 DA 1F 72 DB 53 21 80 CC F2 92 A2 61 9E CE
 39 05 D8 23 5C D4 B2 A8 F0 7B 1B D8 3B C7 33 02
 78 4B 9E 93 49 D2 9D 5F E1 AF 7F 27 83 C1 D7 BF
 4B 05 9F BD 98 C7 D3 EC ED C8 2F 2A BE DF C7 A1
 46 93 F4 66 97 15 43 7F 68 BE 8F C0 45 55 8D 6A
 8D 9E 39 F7 6F 13 60 78 17 BB F3 56 02 39 79 8E
 71 CA 41 28 1D 9D 71 D5 74 B0 EF 09 DD 1E 07 3A
 18 51 9F 02 6E 1F 2D C8 6A 4A 63 8D A0 DB EB F6
 FC 55 27 48 22 1E 2A 69 7D FA F0 75 81 A7 B9 83
 66 97 1C BD 5C 59 38 4E E3 5F 7F F1 EC 87 15 66
 D7 0F 6B 8C B0 00 24 84 E5 F9 24 D0 79 D6 CD 02
 AC 38 F6 F7 64 65 5C 06 FA 51 C2 7D 15 FF DE A6
 57 97 C8 D6 A0 24 57 6F B1 D2 70 3B 58 61 F1 06
 75 02 67 63 6A 32 99 E0 5F 31 98 66 84 9F DE 1D
 E2 73 AC 45 DB BC AF 6A 7D 66 D6 B7 24 29 95 3E
 77 7E F4 91 97 A0 A3 83 F9 88 E6 B4 B3 33 18 F3
 53 F8 64 88 DE 43 90 CB F6 F8 9F 7E 37 63 66 0F
 F7 55 AA A0 5C 1E 91 4F D3 4B AA 16 8D C2 94 F4
 E0 A2 0E 81 30 D9 C9 80 FA 7D CF 26 AA 19 7C CF
 2C FB FA 52 FA C7 25 87 B3 1A D8 18 6B 0C 60 28
 0B B5 C3 9C 28 9A D2 09 3E E9 96 B8 54 5A A9 EE
 C4 2D A1 E9 AB 5F BD 36 2D 3E F2 45 AE 4A 2F DA
 ED B8 0F 15 F4 2A 42 F0 6B F0 B7 95 65 97 51 F7
 74 1B AD 80 77 24 12 3C 33 86 52 0C 25 5A 3D 1A
 02 2E 29 A1 4C B2 91 CB 33 4F 0F B1 95 EE 13 75
 5B A2 7B 4E 08 36 2D B0 34 80 72 44 1F 98 A8 B3
 B9 29 79 1D 3D 12 B5 4C 00 21 16 BF D7 17 61 0C
 A7 ED 4E 55 A2 24 6D CA F8 3C 5D 6A F3 70 AE B5
 46 53 DD B4 DD 10 8D 1A F7 03 85 81 8B 31 16 53
 44 FF AA A0 4D BF E8 51 AF 97 28 82 D0 A4 C9 24
 34 52 FD CA 0A 05 8A 05 D0 7F B1 21 44 A7 20 99
 47 94 7F 56 E8 03 85 C3 59 10 FD EE 13 67 58 DE
 20 56 A2 67 48 F7 C3 A2 92 C8 13 F5 4D 7C D4 0C
 1E FD B5 08 93 92 01 55 19 04 A5 9D 0D 13 48 40
 E5 21 04 FC 06 D0 73 4D 31 C6 4D 53 73 D5 58 26
 71 41 BF A3 B1 14 9E 84 EB 60 36 4C 53 37 ED 81
 5A 4F 22 68 5F F2 82 F6 BD 96 1E D1 1D DA AD 11
 FC 1C E7 2B E4 BF 87 43 57 75 65 A4 1B 55 4D 47
 7A 51 B9 65 F6 38 26 10 1F 3D 92 F5 8A 01 48 0B
 34 FE 8A 13 BE B1 73 FA 13 B1 52 9C 2B A2 C0 3E
 E4 0D E5 A3 E1 76 12 FE 00 5A 2C 91 E4 76 63 1A
 60 7C 35 81 DF 86 C3 86 B5 8B AE E7 CB E0 BA 4E
 73 DE 5F 4A 4B 25 E6 62 83 79 16 94 D3 55 A8 65
 28 BB 94 BC 06 02 F0 22 DB DF A3 2E BE 33 E0 DD
 83 15 8A 61 A4 EA 41 EA B1 89 19 40 2A C0 B0 AF
 D7 AD F3 4E 83 A2 C8 E8 4D EF BB 35 4D FB 79 1A
 DA 3A CA BD 3F 85 2A 7E 5D F7 63 64 4C FF 97 21
 3E 34 C4 60 02 83 68 D5 33 95 FB 2E 45 B4 AF 7E
 91 D9 DF E2 3F BF 16 8B 69 63 DA 22 2D DA C3 36
 FA FB 5B DD 64 81 DA 1F D1 1C 7E AA 0C C0 65 E7
 50 33 22 AA A7 3D ED 1A 69 42 10 28 DE 23 DB F2
 3E 1F AC 48 98 88 58 E2 86 C0 4A B5 14 11 92 76
 53 78 E5 C7 D3 6E A1 B7 C0 1F F0 30 22 EF A3 70
 96 B0 1B 6F BE 4C D5 81 E7 C6 AC 48 08 D4 6F 7C
 87 5E 3F 55 A9 11 6A D7 E2 93 AF 18 6B 12 23 C1
 B5 E4 42 47 CD 07 B2 C5 1F 6A 3A 62 99 B4 80 A1
 E7 A1 7F F8 AF 60 F0 DF 21 9E 3D 9F D0 B9 68 4F
 60 4A 54 2C FA 74 FC E1 70 14 53 11 32 46 A0 E2
 F3 91 2A 75 E0 B0 F0 6D 1F 9D 35 D1 BF 97 1D F0
 E2 84 C0 22 74 4A 38 13 6E 98 3C 0F 50 F3 2B FF
 CA E3 A7 85 D6 3F 68 83 5E D7 32 91 D5 3C 01 C4
 FC B1 4D 69 D4 BD D5 D0 FF B8 07 B9 0D 4A D1 85
 BD 35 3A 74 AB 6D 81 DA 1A 3D 6C 5E 1E 98 3B 22
 4F 1F 9C 26 B8 5E C3 CB 0A B9 17 DB 73 E0 B6 3A
 15 70 1D 0D 38 03 BC 19 82 C8 70 A2 97 D5 78 06
 2A ED 0A 96 45 09 C0 A1 EB AA FF 7A 84 C0 5E 0B
 FD 21 D1 3C 5A 0C B8 E4 44 8D 19 61 97 2B 5A 3F
 58 C9 FA 1F B2 B8 D2 7E AD F1 40 63 F8 60 99 DC
 B3 4C 30 BA 67 8B 8D A4 E0 8E BD F6 C1 3C 87 01
 21 DA 9B 45 04 68 7A 9A 94 F0 DE C2 CC 59 08 05
 0C 21 EA 6D DF 69 4B 80 30 BA 2C E4 F4 52 BC 20
 2E 32 35 BB CE 1D C9 3E F8 AF 15 05 F7 97 C0 43
 7E 42 94 3E F9 73 2D 4A 61 D3 58 95 0A 68 99 5E
 49 7E 1B A1 60 22 91 A4 6D EA 7F 75 0A F8 7A F9
 0D F1 A5 94 72 BF 57 F2 B9 48 E2 B7 D2 E5 3A 4C
 A6 9A 58 8E 7B B2 B8 E4 C4 5E BE 20 ED A6 89 F4
 95 F9 93 B5 D2 5B 8C B8 9C CC C1 A3 4F 60 8E 6B
 9F 63 A6 C5 4F F9 6C E0 D8 6E 7D 62 B7 86 AB 3C
 68 75 92 64 95 D2 8C 64 A7 5E A8 39 60 AA 0B 93
 B9 3D 0E 0A 37 4C CB A6 67 D8 89 84 ED 6B BB 44
 5A A1 C6 F8 14 8B 3C 2B BE E8 C7 E8 8F B9 95 8A
 42 64 ED F1 60 48 A1 2E 0C 0D 53 20 B9 FC EE 1B
 00 FE 3B 27 6D 51 07 47 62 7A 8A BE 07 C0 E6 A5
 86 88 C2 58 FB E9 CC BD F0 A9 B5 8E 18 F0 A9 7C
 2A C6 D5 94 79 12 2C AD B8 06 7C FC 48 B1 C8 E8
 1E 59 CB 7E 3C 22 DE 3E AB 32 F8 CE 9B C6 E9 91
 B0 F6 65 D7 C2 18 1A DB 49 DF 55 AE D2 95 F7 93
 15 B9 66 5F DF 16 2A 61 BF 8B 3A 86 72 4F 78 98
 A9 17 AF 9B 62 F1 10 96 B3 54 4B 37 55 7F 67 AF
 7F 40 D2 ED 3B C9 5B 28 72 90 AE F9 BB C2 DE 4D
 D8 5B 8F AD C1 2A 1F ED E4 DC 38 15 9F 22 E4 3D
 E5 46 F9 97 E3 01 39 ED C9 63 BA 89 D2 F1 CA 12
 55 BA BD 24 4A 3A A5 D5 96 25 8E 85 A4 BF 96 22
 8E 59 4F C3 29 CC 5C F5 88 3F 0A 68 81 04 4E 8C
 67 0C B0 9C E1 60 A5 9F 3A E8 F4 97 74 76 A8 B3
 66 54 0A BA C4 63 11 03 EC 9F ED 43 17 CA 5E A1
 F6 FC 88 DC 5B FF 96 C7 63 64 66 82 F5 BA 2A 51
 AE E9 42 58 B2 82 75 17 4A D8 DE E9 68 06 29 37
 81 7C 76 EB BF 28 E2 C8 FD BF DF C5 21 71 12 5B
 CA 52 0D 94 92 BA 53 3D 0C 2D 96 76 5B F3 0B B1
 44 CC C2 A8 63 5F 38 4B 9F C7 B1 7C 0F 66 57 8B
 82 18 6A 5D 07 47 67 F2 35 CE 18 E2 F4 E7 EC 3F
 94 EC CF B3 11 7C 48 28 33 03 A1 22 76 A9 45 B2
 23 62 D5 91 2E F4 CB F5 3B F8 C7 A3 2A AE 29 40
 6E FD 18 05 1F AC 3C 02 E3 C6 D0 73 5A A8 23 50
 00 02 B5 6B 69 83 63 EF F8 1B B3 73 7F DF 94 D5
 38 80 88 D4 AD 5D 4F FB 32 6F CD 99 E4 00 76 5C
 4F 97 A6 2B 45 A3 95 83 3A B4 D1 9F 5F 71 D2 0C
 0D 69 83 12 98 3C A3 74 E9 9C A1 58 C3 64 EC 44
 08 B1 15 61 4B C4 76 45 8A 83 08 DA AF 51 6D E4
 A9 96 FA 98 E7 9E D0 A9 06 E4 28 31 72 9D 11 19
 D7 07 85 19 ED 7A D2 B7 F7 DD C9 7A FD 93 1C B8
 6F 8A AA 2D B8 38 1C 7F C2 F9 F7 FA FE D3 B6 86
 B7 6A 13 2D 9B F7 5A 3D 07 07 B4 F6 30 47 C5 BE
 E1 E0 FE 47 C6 C7 30 1B DF 9C BE D5 87 09 20 25
 52 B9 B7 0B CC 9B 0B 13 DE 59 31 4E 74 8D 91 F1
 70 09 57 40 23 5C EF EB 90 63 55 23 DA AF BE B3
 F2 B0 B1 8C 68 20 FB 38 93 A6 AD 39 A5 1A 02 AE
 BF 8D D5 AD AA DC 5B DF 5D CF 44 F9 48 A0 BC 32
 99 6B 57 F4 44 0E 80 63 3B AC 58 C5 DC 4A 7A C6
 F5 61 D3 54 4E FE D2 6E C8 79 64 09 31 28 B4 47
 73 4B C7 07 89 2A 86 C5 4C 58 57 D9 D5 3D 67 11
 E1 86 88 53 AF 7E B7 72 8A 8F 82 4D 0D 16 66 05
 3A 12 F4 5D 23 28 7A 5E 21 7A 77 2A 7A 3A A8 F4
 96 C0 C7 C7 51 CC 59 4A 30 F8 6A D4 6C 21 57 5A
 FE D8 ED 21 DE BA 2A C1 16 B6 44 68 05 FB 62 BD
 78 D5 44 16 32 57 72 48 76 0E 09 F4 DE 9D 21 BE
 1B 4C 4B B3 7A E2 D3 4D 35 A6 B3 C2 BD 0F 8E 8C
 BE CC 1E 47 67 8F 72 01 6B 28 D9 A2 19 1B 8A EC
 68 DC DC A3 7C 66 CB FF 9D 56 9C F9 84 A8 63 DF
 5F A9 FC 2B 5A 93 BE 64 E7 D7 8A 28 4F EB 65 BE
 11 08 AD A8 A9 F6 A6 3E C4 74 0E 32 FF E6 7D 92
 E6 98 6F AD CF 8E 33 4C 9C 74 BB 51 65 8D 3F CE
 77 2D 5F 36 8C CD 1F 62 81 80 57 4E 5B D7 A3 D1
 B0 D2 EF BD 09 62 E3 41 34 33 15 4C 04 74 86 D5
 6C EE 04 21 B2 D5 B4 EE 9A 96 9C A1 F3 B3 A4 1C
 8A FA F7 FC 18 5E 88 3E D6 CD 98 BE 5C 48 8A A6
 D8 46 45 A4 DF F4 CC BB BD 97 73 5B AB 81 AB B9
 C1 AF 1E 4E 6B 53 DB 38 6F DF C4 2D 2A F8 F4 DD
 CA 9A 2E 1E D9 DC 87 E5 E9 AC EE 74 4C B3 7D 16
 4D 9E A0 A4 9B ED A1 00 92 98 89 0D 92 59 EF 62
 61 4A 3A 48 F5 8D EF CC 65 A0 C9 F0 A8 1B 5D F8
 94 B8 84 F6 AD 6D 17 40 98 8A 05 F1 34 AD DE 30
 A8 D0 D8 B2 7A 7E 4E 7E 00 9C 7B 51 84 88 B7 57
 0F E6 37 60 9F 77 57 C5 F6 BA 37 44 AE A0 4F 0E
 AE FE A7 8C E6 47 96 F9 C5 F5 73 E7 A9 A7 34 04
 03 3B 48 87 AF 21 29 AC B5 B6 58 09 55 B9 96 E7
 23 D5 C5 D9 97 FC 26 8E 87 FF BF 8D 09 1B A1 32
 54 9F D6 81 34 55 71 C4 19 AE FD 8D 61 01 A4 AD
 57 67 C0 97 85 55 EF DE 1B 5B 26 8C EF 08 2C 37
 7F DE 2E 2A 41 9C 53 C7 82 A5 16 CF 50 0F E0 C3
 59 0B A9 1B 76 2D FA 5F 1A 08 F3 34 FA DF 5D BB
 7A 2F 49 51 53 A2 73 16 7B A8 EC 26 19 09 66 2B
 97 0F D4 2B 3D 03 18 C2 18 44 A9 CF B7 8C 1C 5F
 D8 39 9F C4 96 FC B5 AB DE 36 52 5B 7D FA 32 DA
 03 49 AC 62 7F 8C 5E 52 CF F9 8E 25 4F CD 6D 4C
 9B F5 5D FD 06 43 70 63 6F 76 2B 5A 27 3A 18 E0
 04 79 FA 4D D4 F5 B9 77 4A 01 4A A3 95 20 23 D0
 2A 9F B9 14 98 89 8F 1F FE 13 2E 3E C0 73 ED 0E
 3B D6 BA 12 19 F0 27 39 78 33 3D 75 B9 6A 70 D3
 0C E4 6F AA 49 A5 E6 11 D9 6C 88 D9 1E 30 B8 F4
 91 E4 4D 79 BE 35 ED 51 53 6E 63 92 50 17 F3 97
 90 3D 5A 5D 0A 8B 64 92 59 BE 3F B9 67 3C 71 1B
 0C F7 64 11 36 5E D8 29 4E 69 F6 DD 63 18 C8 98
 75 2C 0C 17 DE 3F 17 DC 6A 69 AA B0 2C E1 C9 1E
 8A 14 3A 71 1C 13 B7 E6 DA 89 CF CF 4C 3B DA 77
 D9 B8 AA E9 F3 62 07 36 28 A2 85 13 C2 04 DD 3F
 BE C6 99 27 2F AA 72 E7 5E E9 DE CE 2F 13 55 C6
 C7 72 A1 9A FA FC E4 E8 55 19 5F FD 86 A3 FD BA
 FD 41 AF FD 2C 9E 0C EF 6B AC F1 63 96 8E C0 41
 F9 60 1F CD 54 EE 2B E5 B4 AE E6 C2 5F B5 9C E7
 9E 7B 40 92 EC B6 79 35 7E B4 44 93 FA 24 DF 67
 C7 D4 2B 29 1D 97 AA 4F 6A 1C 44 46 D0 BF E4 59
 36 29 96 E3 E2 DE 27 4C 03 2F A1 81 41 71 E1 18
 34 CB 16 18 AF 70 00 99 48 D1 89 01 AD 9C 70 3F
 41 02 A3 1A D9 9A B2 93 B5 AC D9 4C 17 80 83 45
 86 05 46 8E 34 64 31 AF 9B 1D 57 B7 B2 82 D2 79
 20 64 E4 E0 AA 00 CD BB 75 B1 C4 B0 03 3E F7 AE
 5B E2 55 AF F0 5B 93 72 0A ED 5F A2 2C 6F F6 63
 53 B1 08 A6 71 4F 86 D1 A7 D0 5A 6F 94 9C D9 11
 00 9F 88 B5 9E EA 65 D5 08 BA F9 F4 CB AC 15 2D
 AA DB DB 63 3C 19 63 12 91 0C B3 2A 37 9E 40 6E
 A9 49 AC 9F BB 53 B2 E8 78 C1 2B E2 3C 0D 96 8D
 91 DE 7B 49 95 3D 61 47 04 C2 51 46 4A 29 11 CD
 BB 4B 11 D2 76 12 2D C0 41 B1 E6 C8 1A 5C E8 F5
 42 C1 41 1A FB 69 24 A7 FA 1C 39 6A 95 9B 30 6C
 65 E0 08 89 D0 EE CC 22 0C 0D 40 DD D1 7F 7C 7F
 8A EE 62 E0 FB 56 68 81 8A CF D6 D3 35 64 69 80
 9A 15 04 11 C6 84 0F BC BA 74 68 75 37 06 21 56
 58 70 F8 90 47 1D 21 16 7C E2 DE 05 B0 30 9F 7B
 F7 E0 D5 6E 10 B4 80 BF 6C 8C D9 6F 04 A3 45 93
 2D 3B ED 64 E8 C9 51 D8 3D A1 F2 8E 82 D4 6D 35
 28 53 C7 31 7E 4E 09 33 0C 83 93 9F 13 1F 59 E9
 5C 27 18 F8 F2 84 6E 30 F2 71 FE 71 EB 9A E6 C5
 DE C2 86 2C 66 7B 48 EE 94 53 01 9D 90 4F B5 22
 B2 CA 68 0F E1 64 18 10 B8 47 43 7A 1D 95 94 E0
 C1 6C 98 34 69 D6 F1 62 2B 12 FF 50 5A 03 03 05
 02 06 DE C5 F8 80 24 09 29 39 BD 5A FC 47 BE B1
 05 44 0E FD D1 92 95 09 C1 6B 00 E7 F8 5A BC B5
 F6 06 0D F7 2A 71 46 91 13 97 0D B7 FC CE 1A 76
 67 4F 61 EF CE B1 62 36 86 0C A7 58 D7 1A 16 0A
 05 DD 54 30 C5 8F 4E F3 DD 24 C4 63 09 F3 60 7B
 9F 0C DF F5 99 F1 4F 4D 5F 60 CF 0B 27 92 D3 4A
 53 86 13 A4 C5 0D 32 21 7A C5 ED B6 C1 10 1E E6
 BB E7 88 0E C9 F9 AB CF 6A 02 8F FD 28 31 45 76
 79 0C A4 CB 2A DE AE F0 96 04 47 03 B7 3B 37 C1
 AB 5D 5E F0 14 75 D5 86 D5 E6 65 FC 96 94 FF 44
 74 B8 E4 B8 E7 CB B2 59 2F A5 36 DA EA 1E 1E EB
 CB A1 3C A5 9B CD 98 9A 5A 12 1F 72 B3 F5 81 8B
 96 6E 77 58 57 88 29 F2 19 5A FC D8 E5 81 F8 ED
 6F 77 93 A5 E6 69 58 82 56 24 29 37 62 0D 59 1A
 49 D6 23 28 2A D7 AA A5 92 47 24 56 6B C8 1B A8
 38 E1 1E AD 14 59 81 54 87 A7 58 1E 6D B7 D7 84
 B9 AA 94 3C 8D A7 19 5F 0F 61 C0 1B BA DC 35 7C
 91 BF E7 81 CF 87 47 42 22 E1 09 9C 23 15 BB 99
 0B 35 23 FB A6 64 1C F6 E2 86 27 B2 24 2A 4E 00
 9C CB D3 D2 CC 7A 64 14 99 D1 20 30 01 81 07 6F
 E7 B8 6E 25 CA 9C E4 43 1F AC 3C 92 32 F8 C6 DB
 F0 23 18 A5 23 7D 90 FF C0 A4 0A 1B 04 8C 3C 3F
 A1 90 40 DA 5C 5D 6E 1E 9D 72 5B 97 C1 90 E8 EC
 EE ED D6 7D C7 27 A7 64 E9 DA 70 A6 EA AC 94 E1
 66 5D 8B 83 D6 5E D6 B6 D5 C5 25 97 85 61 F7 BB
 CB 2A C3 90 B3 E1 3A EE 13 77 BB 47 75 55 9A C2
 FF C9 C5 98 BF 72 75 D4 F5 D4 68 35 27 E9 E8 E5
 4D 3B 93 DB 74 22 D1 D0 8B 48 75 E4 48 17 9A BA
 C9 4A A3 B2 F7 8D E2 E7 22 D7 B1 35 25 D4 B1 80
 CC 59 FF 5C 12 5D D6 96 8B D2 79 8C B8 C7 47 1A
 CA B4 58 03 1F 2F 1E 5C DA A2 9A F7 C4 CB DE BA
 C0 64 DC 2C 47 E8 2A 1A 3F E0 8D 70 50 B2 A7 55
 DC C3 D9 75 97 2E 95 34 26 0F 2C 8A 2A E7 EB AC
 3A 1C 2C EE C7 B5 5F 34 79 00 79 8E 13 B6 3D 91
 10 D5 DC 3B B3 C8 0E 09 BC 9A FA 0B 34 C7 31 55
 77 9D DD 4C 29 46 3D 99 49 F3 DA 2E F5 F2 F5 0C
 81 57 1F E3 CF D0 C9 44 3D FB 3E 78 C7 70 1F 40
 EC 20 D9 D2 58 7E 25 4A 87 F0 B8 04 29 20 70 B7
 94 5C 43 88 8B 1A 4E 34 30 A6 9E C5 92 8A 1A F5
 E8 2C E3 95 8A 6A 14 26 42 4A 87 5C 8C 3A B6 CE
 8A E3 4F 83 7B 3C FE CF E5 73 6B CB FF 21 F6 B2
 CE 8C C3 4A 8D 7D A2 9C 21 DF 1C 52 06 96 27 3F
 7A CD D0 15 D1 50 69 C9 4B 63 A6 67 1E D8 49 1C
 50 B7 D7 CD 6C 2C EE 7E 82 8F AB 9C 2B B1 56 68
 79 69 AF FD 21 33 73 AE 69 F6 60 D6 EA 2C 34 E5
 74 5E 3D 2D 83 25 41 BB B6 AC 02 49 D4 1C F7 48
 E8 A0 50 61 A3 50 D6 EC 10 A7 26 72 4C B9 DF 2D
 56 60 ED DC F4 4D 42 8A 1B DF C1 0B 8B E2 93 50
 23 82 0F C6 84 07 ED AA 66 76 13 01 2C 74 ED 9E
 13 6F 0D 6E 36 31 ED 80 93 82 CD B6 A0 BE 07 17
 BA 91 37 D5 5F D0 32 3C 20 9A 36 FC 32 67 65 46
 52 A6 D0 11 D3 3A 31 D0 EC 99 09 2B 6A 99 C2 4E
 A1 4D B1 EF 49 79 1B 96 FF A7 76 B0 CD 7E 97 1A
 44 2D FC 7B FA B7 4B E7 81 B6 15 E2 B2 B3 83 49
 FF F2 2E 6F 31 D2 67 2D AE 9A 47 92 84 A9 3E 06
 BB 7E B1 5A 5B ED 11 77 71 88 0F F7 4E FB 8C 16
 70 AF 56 40 3D 05 77 CA 8C 26 5E F4 4E 31 8E 53
 59 2A 6D EC 61 DD D3 70 1A DC 60 96 49 C7 77 E3
 48 D9 E0 5B 5E 21 BF A1 57 91 7B 8B 78 CE 11 1A
 FA D0 2C F1 22 92 8B C1 7C 7E C1 68 F0 8D 13 90
 E4 E8 C3 A8 95 15 63 9E CB A7 41 91 87 3D 6E 69
 E3 76 CA A3 CF 21 19 AF 36 EF 9A 97 B2 0E 24 73
 FB A8 83 21 AE 71 DE 1A A7 34 8C 93 FA 71 19 C8
 E2 19 F7 C7 B9 2A 22 B4 16 15 B2 03 88 EC 23 BC
 EB F1 CD 85 01 50 EF 69 DB DC 4B 2E AC B8 DA A0
 6D A2 86 51 FF 8E 3B E0 1B 66 7A 11 3D 9B 76 74
 9D 7E 71 28 B3 D5 B1 A9 1D 65 9C B3 55 7A B5 F3
 2D 3E CB 9C 4F F0 D8 02 B4 37 52 E5 E7 D9 78 D8
 50 14 08 F7 0E 14 C0 E1 E8 12 58 A0 4B CE 36 49
 ED 0C EF E4 25 0D 1B A3 2C EC FE 1B C6 A5 E2 2F
 5F E0 FE F7 3F E1 E6 B3 A8 9C 18 FA E9 C1 25 B5
 F6 C4 1D 59 50 31 B8 21 1D 5E A3 EA 1E 25 AC 3A
 B7 4C 0D EC 64 3C 03 0E 4D 01 6E 3E 5C 45 65 21
 91 69 A5 FC 9A 1E 99 B3 0E F2 F3 0F A2 26 5E C8
 B1 71 FF 31 29 70 CF 6D CD 3D 64 79 D9 C0 0C 52
 5E DF B2 92 F3 24 38 A5 B6 06 BA A7 94 C5 C3 67
 F5 58 F5 81 C6 99 FD 73 EB 94 66 EE F9 AB 26 F2
 DA 9D 9C 8F 41 A7 F7 A1 FE 0D B0 BD 66 B4 9D 8A
 88 D3 1D EC A2 83 35 47 E5 C5 EF D0 C0 10 E9 0D
 7C 6E E8 1F AA 04 52 49 4D F7 9C 3F D3 E8 E5 DF
 41 26 C6 70 AA 5B C1 04 3F 79 C2 5D DF 3A C2 17
 A0 7C ED CA AC 9D 06 A0 D6 A1 54 1E 4E 1B FA 8B
 D8 CE 42 30 93 1A 57 A9 74 0A 93 1F 6B 6D 54 EB
 A6 90 81 22 BA D2 BF 59 FB 69 E5 78 44 D2 B2 32
 71 D3 9A DF 05 49 A1 0F C8 65 F7 C2 5C 26 52 70
 D4 FD 09 05 FD D3 38 7B C5 A7 3E 2F 88 D2 7D E9
 D3 C4 98 09 8D 0C 96 99 8E 9F BD 39 92 B8 FC A8
 A3 C3 6C F6 97 11 25 13 D8 4B BE 98 F3 CB 40 3A
 A6 11 E6 8D BA F3 8C E4 98 6F 6A 7C 7C AB FE B7
 E7 4F 8F 4D A0 6E 37 F1 FC D6 9F EF AB 19 EF 49
 E8 AA 47 45 8B C8 93 E5 BB D5 F7 9B 3D F1 28 FE
 AA 03 29 01 4D 07 82 78 EC 26 B2 83 AC B9 F6 9F
 53 E4 62 A9 8D 98 6F 49 74 2A 9D 23 B2 1E 3D 3D
 10 04 3F BD 9D 11 3E D4 1A AA 51 24 80 EE 82 7E
 98 26 DA EF FB 6A 10 D2 EE 8A 35 55 B2 69 AB 86
 7F C1 28 E5 7D 0E CB B1 2B 90 1A 35 82 F2 4A 69
 1D 1A 44 06 2F 55 65 C0 24 1F E3 20 00 DB BF AE
 83 24 F8 4B 17 93 42 F3 95 D1 A7 AD BD 2C 48 6C
 7F 1B 43 34 67 A4 94 D4 EB 61 A6 31 0B C6 9A 2B
 8F 87 42 E8 2B DA 1A 1E 06 2F D7 56 77 B2 D2 7D
 F2 48 A4 9F 6E 39 17 A8 94 25 A1 44 F7 BA 65 3C
 69 B8 E1 5E 10 C1 52 91 1F 7A C3 11 EB 8C 55 76
 7B 84 07 11 E0 6E 8B A2 8B EF AB 10 D5 62 73 57
 E9 F8 AB 97 7A EC 5E DC 6A 9C 27 82 B4 41 CF 51
 0E C0 B0 3A 42 DE 70 74 09 AF B3 18 C2 F2 6D 98
 FC 7D BA 3C A6 35 C0 C6 A2 CD 5B A0 B1 27 76 27
 D4 43 73 39 D5 51 24 FC 28 90 C6 26 E6 1C 3F FA
 B0 64 1B A2 14 13 71 EF 72 85 11 16 23 8C 9C 15
 9E 5D 86 5E A5 73 D5 17 BC 70 A7 DA 65 49 4D 53
 C9 BA DA C5 4A 3D 60 0B F9 E9 98 F7 15 31 8F F7
 0F F9 9C 14 87 53 C1 50 54 F5 D3 4B AC 1A E6 32
 E8 D2 F0 66 E7 48 4F 66 8E 8C FB 86 0C 88 B7 34
 DE A6 AB B0 F6 6C B9 09 FF 5D A5 79 5E E5 98 E7
 45 4B 49 2C 1A 6D FD C6 E4 B2 90 C5 45 0B 0F C5
 28 DA FE 28 B0 B0 0E 01 1C 8B 78 38 0C 16 A0 AF
 EB 30 CF 4F F4 15 00 12 5B 5B 1C 57 FA F0 CD 86
 E7 96 87 1D D9 2A 20 2C 52 DA 27 2D 25 EC DD 69
 B4 D9 BF EA FB A2 FC 27 F7 1E EE 7D 33 85 88 19
 F3 83 CE 9C B5 21 82 EE 9F 2D 20 EF 07 5A F1 AC
 53 53 67 E9 14 BD 1A 44 06 D8 9D D4 09 58 E3 15
 6C 0D BE 7D FF 36 A9 9A 08 DA 17 02 76 83 85 43
 6D EC AF 4B B8 56 42 80 FB 99 58 D5 5D B3 9B 0C
 1B 20 68 90 9A 27 5B B2 7C 0D B7 3B 0A A8 F9 2E
 89 CB DD FF 09 BA C2 86 E9 B5 52 61 D3 99 E0 13
 06 75 30 1F 46 47 EE 8E 40 64 DE DF BE 93 93 C4
 3A B2 01 09 6A 73 70 F7 59 F8 19 5E 31 C3 D3 D1
 F9 3A AA 9C 18 A0 D3 FD 16 47 D6 8E 37 1E B1 83
 E5 74 9B 9C ED 88 BA 37 3D 4E CC 08 3C FB C7 B7
 6F CC 35 71 04 83 47 21 18 D7 BE B5 1C B1 06 20
 F2 ED F8 55 1E BB 7D BE 42 2B 08 44 3E 1E AF 56
 C9 44 16 B4 D0 46 05 BB 49 8A D3 10 BD D3 F8 1E
 37 08 B2 34 99 CD 4D 3D A2 C5 C7 32 26 92 71 4F
 A6 3D 49 20 97 A5 22 7F AC 20 63 85 3D 88 CD 34
 7B 8D DA 7E 81 6C 4E 62 71 71 2F E7 01 59 B3 18
 76 4E 05 A5 C4 D7 6D 5A E3 B8 41 9B 63 81 49 6B
 80 6E B1 64 7C 4B 61 F6 32 A6 93 9C 7D E3 8B A5
 E9 B2 D8 14 1F 65 FE C6 92 C4 B9 7B 74 8F 45 A0
 5D 30 9C F3 A4 6B EF 1F 03 D6 E0 C9 4F 57 A2 6C
 27 4E 63 93 1F 59 10 71 32 E5 8B 50 86 7D F0 D8
 85 24 2F 67 9A A9 83 6D 37 7E FB 62 3A E8 82 2B
 0F 36 3A D6 E5 33 95 EB 5B 7C 8E 3E F0 F8 DA 06
 03 39 ED A0 87 5E 74 D5 49 58 F9 E9 0C 39 BB 6B
 1B 8D 2F 29 9A D6 56 66 35 6B F4 B3 91 EC BD 03
 0F 54 F1 22 66 AA 3C 18 FE 10 DE 9A 91 0C E4 4C
 E7 66 D2 92 C4 9F A6 F5 28 EE A5 C9 74 42 C6 D6
 31 5D F3 D0 54 01 AC 5F A9 B8 F6 75 CD A1 BA 05
 6A 4C 52 EB 81 E6 C8 92 32 D0 4B 08 3D 24 29 E4
 4C 4B 55 5D 7B 02 B9 75 F6 7A 84 12 79 1C E9 EB
 07 BA 95 12 B4 59 43 CF 21 B3 22 93 84 FB B5 91
 B5 66 7B BD F4 B0 8A 48 5E 29 8B 84 5C 91 A1 99
 86 5D F4 22 08 17 33 E9 49 9C BC 50 4E DE 3C 82
 93 D0 FB 35 A7 85 C3 04 0C E9 B9 6E 14 73 0B 36
 1B 49 3D 5A 0D 66 2D CC 77 FE 14 03 5E 11 1A C3
 AD D5 59 57 6F E4 6E A5 CC 53 9C DB 00 56 77 BE
 B3 94 ED 63 9E 95 D3 79 F6 F2 E1 85 7D 9D 98 E6
 88 14 0E D4 9B AE 05 33 39 3D 08 3D 85 BD C0 47
 1F 92 39 6E 7A E7 E9 A8 8B 23 56 29 15 0B B0 30
 F8 BD 2A 91 5B 6C F7 2A A7 57 31 98 04 2C 2F 87
 A3 E2 AF 48 B3 CD 7F 91 BC D8 A8 D9 BD 27 84 D3
 0D 93 4F BF 30 3B 4B 16 42 C0 95 AF F6 38 63 D7
 70 3E F7 45 5A 9E 2A BF 44 0D CF 6A AB 10 56 03
 56 95 90 69 10 CA 00 17 9D 61 64 EA 16 FA 71 46
 94 C4 29 CF 77 A5 FA FD 48 D2 BA C9 38 EF E2 F7
 BC 39 64 5A DB 69 1C A7 72 74 D1 4A 16 2D 96 CC
 F2 46 B0 C4 AA BE 3B 82 AB 55 25 7D FA 63 41 B3
 11 9C 9D 68 CA F2 38 F3 B1 C4 62 1D E2 5A 4B 31
 6E 62 22 2E 56 00 A2 11 0C F5 81 94 10 C9 49 F7
 C4 6D 44 69 4F 4A 58 1C F3 31 B9 4B 11 AD 51 35
 C2 68 A1 DD 9C 02 01 BC 40 B0 22 55 60 46 4A 08
 0B 8B B4 D8 69 43 AE B8 E7 82 C6 1B 91 07 BB C9
 BC 68 DB 98 1C 8B 4D 49 B8 F2 E2 28 5B 68 1B 2A
 67 DF E2 F8 38 83 F8 63 B7 AF 4F C0 0A 72 5A 5C
 84 BE D9 2A 4A 5F 5F A8 02 C5 88 14 83 E9 09 08
 E6 57 AA 09 76 3E 8E F8 56 79 FC DE 1C 27 79 C5
 AE 42 7E E7 3E EB 46 A4 5D 56 2E 77 3C 46 9F 19
 2F 05 9A 08 80 AB E7 C9 DE F8 D7 82 0F C4 63 00
 3D 5C E9 A8 D2 EA 2F DC 64 8C F5 F4 3B 3B FC 16
 33 32 E3 4C 43 84 EC 0E 73 B2 BE A9 8E 59 8A 6C
 F7 36 AF F2 68 17 86 7B AF 3E 62 DC 8A 08 B8 AC
 E9 47 68 61 98 C0 31 81 F6 4F 62 45 1D 96 F2 4A
 DB 93 E8 64 2B 6E FD 56 D7 9D 10 B1 D2 CA 4F B5
 68 21 12 5D 6D 93 3F 6E B6 2A 10 E6 EF DE 68 01
 CD A4 FE E8 79 C4 B1 A9 D4 C3 CD D6 D0 97 15 EF
 FD AE 22 77 48 76 E3 F5 5E 91 53 C4 32 57 C4 23
 12 A7 BB D2 9B EE 8A 4B 6E 1D A0 35 BA 9E 89 7A
 29 09 9F 57 36 D8 F6 AF 15 6D F7 8D 4A 8D 16 0D
 98 34 48 3B 24 D1 A5 91 D2 E7 2F F5 63 75 A3 AF
 6E 6F 5A D8 61 7C 67 85 1B 38 4E 59 89 E8 2D 44
 98 7C B5 3A 41 CA FC 0D 8E DF 69 61 82 F4 07 9F
 4B 14 BF B3 5E 7B 7C 55 26 26 6E A6 37 54 07 9C
 F9 AF DE 70 BE 9A FE 74 72 1C F5 99 19 2B D5 5B
 8F F0 4F 85 AD AA 4B 39 58 3D 20 8D 75 2C 2E 89
 73 64 C0 C9 21 DC 7C 19 D1 51 1F F8 0F 16 FE C5
 CE 1E A0 9C D8 64 29 34 C5 6D B4 AB 9D A5 22 77
 E2 B7 31 32 62 6D E8 54 95 5D 43 E2 96 C5 E0 9A
 3B 6E E0 0B 3A 32 2C F2 26 03 7B 3B 05 89 30 D7
 63 43 60 78 9D A6 9E 76 47 D3 E2 AE A1 A7 58 20
 73 0C 26 17 6E 7E 4A C6 B0 9F E8 80 A3 E1 AC 8E
 35 25 23 17 68 7D DB D1 9C BA 44 8A 17 2E CF 93
 8A 31 A9 C4 33 64 72 CF 9E EC 58 FE 80 7A 65 75
 A8 5D 50 6F 07 C0 D3 A2 79 D8 FC 25 EB D0 FD CB
 44 C5 95 44 D9 DF 31 29 2D 67 CD 05 DD E2 19 11
 E8 B3 70 1E F9 53 98 B1 BC B5 54 5F 0F CE 53 8A
 7A 43 FB 95 33 63 62 53 BA 3C 28 F0 3F C3 5C 50
 E9 9B 78 7E 55 99 CF 50 3F 47 9B 64 86 37 5D 97
 BA 41 9F FB D7 CC C9 4B 7F F7 6F FF 82 9D C5 DD
 02 52 8F C0 B8 EF 81 5E 23 32 EE 7C D6 E1 62 37
 B4 0A 2B B7 F1 52 77 A4 D4 11 81 3C 05 D8 CB 91
 EF B4 13 6E 42 58 79 BC 8D B8 65 4E 5A 3D F1 FE
 F4 C0 60 CE E3 05 1E 88 C2 36 67 A1 26 DB 14 B6
 CF C9 3A DE 9F 97 46 02 36 10 71 DC D1 CD 25 04
 E3 E8 A6 D6 1F E8 76 28 A5 B1 10 2F 46 FA D6 E1
 F7 4E 52 D9 90 91 58 94 13 71 8F A0 16 36 E3 21
 A9 A3 44 D4 BA 77 40 2B 6F 5B 27 CC 49 E8 B6 C1
 72 FB D2 79 E7 85 5C D3 15 45 2B AA 21 F3 BA AE
 A3 74 9B 7B F6 59 1B 15 4A FB 6C B8 CA DC D7 1F
 72 7B 27 C0 8C DA 5D 07 84 92 B2 F5 DA 2A A7 37
 8A A3 A4 5E 86 BB 63 9A 42 64 E1 48 09 51 3A 46
 64 E2 33 AF CF 64 0D 2A F1 AA 57 5F BB D6 BE 7E
 C2 99 57 5D 7D 5F 02 D2 32 BA EA D1 6B 29 94 52
 9E BC 22 4A EC 53 34 47 FD 89 D3 4C B3 2E BC 14
 17 8C 57 09 AB EA 43 8E 0F 71 E7 BC 96 85 BC 40
 55 77 6C 9D A8 E5 3A 02 1B AF 61 25 D3 CD DD 42
 33 11 E6 AB E3 FC 12 28 23 F8 19 2A A7 3D 90 58
 9B F2 31 3B 3A D2 0F E8 E7 12 64 A6 D9 73 8A A3
 59 4F AA 58 1C D5 1C 75 33 59 E7 08 91 9F E9 EA
 21 06 1D 1F 47 44 59 0A C0 F2 96 98 38 87 74 E3
 E6 9B 3E 0A 40 39 57 34 D7 0D 03 A5 09 3B EA E6
 0F B1 88 8B C2 2F E5 E9 81 1A B8 B3 74 AB E1 E9
 05 1A C0 0F 82 08 12 E9 6D 6A 79 3A F9 E0 FA 53
 0C 4C 5F 55 4D 04 D4 2E EE 94 90 36 05 40 32 24
 08 EB 37 60 9B 25 9D C5 75 95 AB 5D 9F 6D 46 85
 4D FF B8 B3 1D 84 0F 22 03 A3 43 80 2B 84 D1 E4
 D5 AD 63 A9 B5 87 3A CC 61 F7 D4 03 30 59 8B 46
 D0 08 1F E6 19 0E C6 8E E1 0F 26 D9 16 E8 DF D4
 D7 3E 15 B9 68 83 A6 86 93 13 A1 87 DF 9A 15 02
 ED AB A7 EE 1C 0F F5 3C 49 96 86 D3 E0 6A 82 A1
 B0 6C 11 36 96 6A 9B C6 C1 75 54 52 09 F0 6A 36
 A6 AF 6C B3 E8 DF 6E 6A 35 F1 40 83 45 A0 B1 3C
 3D 51 0C 84 14 DF 30 80 39 56 C4 B2 D1 62 C3 5C
 92 2C 23 AC E2 D0 13 8F E2 EE 50 2F AE A7 1D 69
 BB 6F 2D 03 E0 95 55 D0 68 EC 4B A8 EA 03 E5 BB
 DE 67 91 5C 19 D8 94 54 E6 33 06 C6 8E 45 28 FE
 F1 E8 D8 2D BF 5C CB 82 05 3A C2 DA 5D 99 5D 82
 F8 6F FF 1C 78 30 E6 15 67 44 B9 6B 07 67 88 2B
 DB C6 79 01 E0 D7 9F 43 10 A3 FC 6E 92 E9 10 2B
 88 E7 17 5E 83 6B 88 2A 87 64 64 FE 3E B0 9A 8F
 50 24 86 B3 05 8E B4 C8 A6 5B D4 88 F0 CA 7B F5
 E6 41 D4 9B 44 EB 3D 45 DA 38 00 D4 28 7C 04 73
 A8 78 22 43 98 A9 EB B7 0F D2 53 0F 47 0F 65 D3
 61 43 FF 9C 9A 67 CF 7E 60 85 FA 8A 18 88 4F 87
 87 DA 32 18 54 64 41 F3 2B 3D AB 17 F8 D1 3E DA
 63 9E 5C F7 77 59 45 64 D3 96 65 AA B8 85 C2 76
 3D 00 B4 F2 EB 6D A4 BD CA BA 2D E3 A0 72 0F 8F
 6E 93 2D DC 10 9F 20 D0 67 3C 7B EB DE 0E 4C ED
 73 FB 55 D3 CF 38 30 F2 5E 7A 93 C6 5B 5A A3 46
 86 D1 8A D8 13 6C 03 E0 E9 7D 66 42 71 ED 28 D4
 93 DC 3D 64 98 38 45 12 E6 27 66 18 F8 CD 28 EF
 D7 F2 84 B2 03 9D 57 7D 51 0C AE E2 F1 94 1F B9
 8F 14 55 27 30 08 FF 9B 14 E8 44 08 8C F1 D7 55
 B3 D3 19 E1 75 F8 3B 7D E5 04 3A 9A AD E9 79 38
 48 62 09 F2 F1 0E 2D F8 DA 90 41 77 5C B1 FB 5C
 C2 C7 E7 3E EE 6C DF C9 14 60 79 39 4F 7C 4F FD
 4B 5D A0 55 E5 12 31 E1 C2 48 97 85 FE 20 8A 07
 41 E2 5B D8 64 3E C1 AF 94 E1 F3 C9 3D E8 17 E0
 03 20 70 15 98 D7 3D 30 61 4E 97 49 47 FD BC 93
 A4 73 F6 78 E8 A5 13 F3 72 EF E8 BC 23 62 E8 B9
 7E 89 9F 19 11 38 36 0F 63 74 4D 23 4A 74 60 D9
 5C F0 AF CC 7F 99 4E C3 E9 CE 64 B6 23 AE 3C B6
 56 F0 3B C5 2A 6B 85 10 9C 12 6C ED BD 57 C3 E9
 80 7C D7 B3 93 B2 96 01 3C E8 A4 99 C7 52 A3 51
 F9 71 9D 9F 50 80 21 6C E2 1A E0 BB AD F9 5C 8B
 96 AF F1 CA BF 03 2C 8D 8A 07 EF 05 75 FB A0 E3
 9A 9B 86 34 0A FC 25 60 85 A0 68 02 94 01 2E 99
 8C 77 02 8D 90 00 4E ED 82 3D 7F D4 AF 9B 9B 3B
 16 F9 EA 45 A0 88 23 65 23 81 D4 4D A1 9A 91 9D
 42 3B 7A B8 67 BF B2 57 78 E7 01 DB AA FE FF 6C
 ED 0E 07 41 14 52 5A D1 C3 97 44 BF 07 78 04 4F
 D1 62 E1 5C B2 DA 62 0C 6D 85 6D 3F 41 84 8E EA
 8C 24 5F 90 BE 88 84 EB 39 16 45 E5 3C 07 D7 30
 9B 71 7B F0 9C 4D 7F 3A 15 FB E6 C7 89 E1 C2 F1
 DE 54 77 43 72 4D DE 25 72 55 38 00 B8 20 28 CA
 6E 19 F4 5C 28 00 E9 5B C3 2B 86 6F 25 BA 33 37
 6A 61 08 1B B7 36 DC B0 24 D4 DD 02 39 8B 76 27
 B9 9B 0F 84 3E FA 81 20 7F E2 8B 66 03 D3 5F 4C
 25 FD 5C 20 A7 F4 98 C7 83 33 BB 0A A2 6E 04 28
 FC E3 76 10 92 18 63 D4 F7 7C 89 FC 9F FD 63 82
 44 5E E4 81 BF BF 4E ED 68 45 61 92 FB 3D C3 DB
 14 B7 DF 4F CB 28 4D F0 CB 8B B5 50 57 96 8B 15
 86 53 F2 74 57 5F 00 69 9B 63 EF 7D 1D 30 B0 B2
 44 43 99 AC 2C 2B 2F E6 BA 38 6E 56 21 F9 8D 5B
 83 D9 69 23 6A 78 4C 08 05 4B 66 BA 05 80 59 02
 9E A2 0A 01 F3 2A ED 7C 2A 38 B2 4D B5 B3 83 39
 04 B4 C2 47 2E D4 E4 2D 92 78 CE 0E C4 B4 8D C0
 EA 02 6D 93 EB D4 E0 42 9C BF 37 C4 2D 6C C9 EB
 D6 E2 59 B3 42 E7 4B 3A A8 9C B6 97 8F 54 0B F2
 B3 CA 23 15 5F FC 26 CD 2A EB 02 61 6C 54 9B 8C
 BD F6 6F 9F D2 41 51 BD 75 43 AF 04 E4 65 3A 2C
 97 C7 DC 97 61 EB 17 99 1B FC D8 B2 B8 E2 CC D5
 6A 49 00 93 81 D9 03 33 DB 8E F4 9D DC E4 94 B1
 C2 4D 76 70 5D FF CC CF E5 D2 92 0B C7 B8 BA 2F
 45 EF 45 51 88 50 EE 9D 59 4C B6 31 E6 0A 83 CF
 A0 87 76 06 CA 2D 1F 09 09 F2 1F 1E CB F5 89 04
 B4 12 2A 1D B7 88 85 61 59 B7 1F D5 EC E2 2A B8
 07 AC FA 27 1D 82 DF 5C 8A FE D3 9D B9 04 C2 E2
 8D 3C 52 43 6B 50 AA AE 58 E4 DF 79 E4 81 AF 43
 50 B5 A9 9C 42 28 86 7E 11 41 61 A0 23 85 09 F8
 EC DF 8E 72 57 37 48 D2 04 7D 39 FC 4A A3 D6 91
 B4 C2 01 43 9A 8C 4B 10 81 CD EB 7B D8 94 38 49
 05 09 1E 8C 2F 99 2B EA 38 99 1F DC A5 2B 27 20
 0A 69 C6 B4 EB 47 29 51 A1 86 14 42 97 AD 5D 55
 25 F8 DF C5 C2 07 6D A0 14 AB 35 9D 0A B3 3E 6D
 E6 7D 86 55 DB F6 9B 20 7F 3C 48 4B F5 49 B0 F2
 F5 AC 61 01 00 3F B5 EC C4 A6 7E 99 6F 48 0B 5F
 25 2D 33 4F 06 5C C3 33 54 E3 12 38 69 30 FA 45
 57 6C CE 18 A5 8D 60 08 C2 EC AB 9E DE 93 33 2A
 9E 4E 2B 9C FA 39 14 9A A2 D0 7A 5D 65 73 0C 15
 A3 40 6F 8D 4B 8E 4B 9B AC F3 6F AB A8 43 4F B8
 E0 BA 58 F9 47 A6 5C CC C8 0D D1 92 E0 A2 82 5A
 5D 8E F8 59 D9 04 76 A9 0F D5 33 3B D2 FF DF E0
 46 9C D6 92 14 31 DD F2 E3 64 82 92 B5 9C 21 DF
 0E 2F C0 38 E1 5A 3F 15 F3 5B D4 BC 8B A0 BA 72
 13 71 D9 7C F5 71 81 3D D2 A5 D6 F1 F4 19 9A 6F
 5C 0C FB 78 EB F9 E5 5C AA C1 85 72 BD AE BF 79
 C7 56 35 34 6B C5 FF 31 FB 8D 0F FB 98 81 52 EF
 56 39 F7 38 90 A2 6E 9F DD 3E 83 36 05 12 B3 C6
 C8 5D C1 F7 08 A0 8E C0 5C 08 AA 7A 49 ED 49 7A
 27 42 CE 14 A8 48 A0 2E 97 49 81 B0 7A A8 BF 84
 8D 02 93 D2 3C 63 7D 3C E8 1D D6 EB 83 D0 CC F0
 C8 D7 79 73 AD 5C 8F 21 87 A2 6E 93 58 4D A9 10
 79 84 2B B3 46 92 FB A4 B9 80 F4 C5 DC 61 00 A8
 6F 9E A1 1B 70 9A 4B 6B 70 13 9F 4C 75 A1 C4 EA
 2F A4 DD C0 81 02 15 5E B2 35 32 72 FE 25 88 3C
 CA E5 59 FB C6 D0 48 10 A2 56 49 90 2A 4A C2 5C
 7C 4E 62 4F 1D 65 1A 87 BB 8A 9F EF A2 80 1A 27
 01 78 27 A4 CD 58 6C F9 A7 9C 6C 17 92 8F F0 0A
 F0 8F BF 4E 28 3D 57 85 4F 10 AE BB 0A 48 2C A9
 7A 47 80 4C 66 51 5B A8 F1 BB 71 CB 80 49 1C 5D
 8B 4C 08 1F A8 57 7F 31 8D AA C8 F1 70 C2 D8 39
 0C 77 5D 98 AC 2B C7 34 64 FD E5 FA D5 96 87 8D
 61 9D A2 40 37 AA 56 7E 41 F5 7A B5 CF 4D 5D F1
 14 2C D0 80 49 1E D9 81 28 49 CB 66 93 85 8B CF
 A3 77 FB 70 20 CB 01 D9 F9 B9 F7 54 95 CC 8B BD
 1D 28 6E 28 02 1F 7D 5B 0C E2 96 39 33 F4 EF 1B
 A9 98 D5 A5 69 CE 1B 7C 5D AE 51 79 1B 2E F3 45
 2D E4 8F 53 0E 08 21 FF 68 68 C1 AE 7D 50 D5 15
 EE 24 49 74 69 C7 83 99 94 65 DF 2C A2 19 BB BA
 B5 40 9F 6D A9 80 1F FD 5A 2E 25 93 2F F6 92 9B
 04 38 36 9E FD 83 ED BA AA F5 52 D0 8F 49 B8 00
 C2 EE D0 98 93 CA 7E 00 6D CF D2 E6 79 9C B5 26
 F5 EC C9 F0 4B E7 24 42 44 AE B0 C8 D7 64 FE CB
 D7 CA 80 91 77 93 98 C4 4E 32 F5 90 01 D3 77 97
 CE A4 06 E8 3E 7F 79 E9 C6 5F A8 39 51 7C 14 D7
 BF 02 78 37 B9 37 8F C3 68 BE BF 63 B4 D8 F7 FA
 6F 7C F5 8D FF CA 9D 15 5A 59 5F C0 9A 08 60 9C
 13 C4 6B 4E 5D A7 EC 4D 9E 96 46 B7 BE 8D BD A4
 59 DE E8 28 B4 59 DD 79 21 51 F0 8C 8B C9 B9 8C
 3E BF D1 54 E9 01 39 B0 02 9D C7 30 F7 07 3E 0C
 04 0C FA A1 35 77 80 84 9B 87 53 D9 8E 88 07 EB
 D2 55 85 5F 56 9A F3 3C 5C FA 0C 9A 26 DB 17 4B
 E9 F6 CD B7 49 D9 C8 94 A3 C3 2E 90 2A C6 23 7F
 69 0C B7 25 B5 78 2A 6F 78 56 DA 5E FA A9 6D 85
 CD 5C 7B C5 70 83 2B C2 5B D7 D6 D1 B8 F9 4B 7B
 CB D5 AE 40 CF 3A 9A D0 A8 35 4B B1 79 37 69 93
 DF 3D 65 41 BD 3E DF 77 C1 CA 1F E5 39 16 70 45
 83 50 AC D2 D7 68 40 FF 41 C0 6F 85 6F 8C 62 66
 F9 6D C7 8E 73 F7 3E 44 61 E1 D2 DD B8 9E F9 31
 4C EA 66 BB 38 D2 12 24 CA D6 F1 7E 68 CA 52 FE
 08 F8 36 D4 60 A8 1A F9 8C 33 18 BD 26 AF 84 55
 3D 9F A8 33 3B 8A 91 76 7B C9 4D A4 7F B2 86 B0
 DC 11 54 FC B4 C6 F9 2B AF 30 B3 56 D7 1F 71 A4
 15 7F 05 B5 A0 70 FD 0E 4E C2 DA 89 42 2B 29 D2
 55 5A C9 30 E6 D8 E1 39 C8 8E 97 0C B7 8D BD 25
 35 7A 8C 4F 56 6E AB 5A 6C E2 74 C2 BC 42 55 06
 B4 E1 D2 27 2E 57 B3 94 76 72 17 8B 89 1A 84 B6
 FA 8A E7 14 09 32 7D F9 B3 3C 80 9E 51 15 75 4F
 95 D4 42 01 EA CF 7A 5E 0E 31 F7 F2 39 DD DA 13
 98 DB 7F 8C EA D6 0A FB 9F FF 3C 03 AE F1 0F 4F
 C2 B8 C1 87 3D F0 F7 14 22 13 7E 25 4D 57 7E D3
 40 C2 D7 8C F4 E6 76 B8 01 18 C5 33 3B B2 AE 81
 DC BD 84 FD ED F4 0D A5 E6 56 DE E0 6A 82 59 C6
 8F 9B 37 78 93 F1 97 ED 57 88 FC D1 0A 22 17 D9
 42 FB C1 41 0D 55 0F 81 7C A9 11 3C 02 BD B6 2A
 EC E6 D7 49 A3 AE 91 33 0A 91 50 20 58 7E 16 DB
 0C F4 45 26 77 76 34 41 4C 0B 15 A7 4E 31 65 14
 39 CE 3C E6 A4 1B 0E 72 DE 1D 79 4C ED 1B EB A0
 3B E8 4D 57 AC 90 41 00 EF 0D FD DE F0 15 F3 04
 21 A4 24 DE D5 02 0C 16 57 ED 15 8B 0F 51 69 2B
 19 A3 92 D0 85 E8 6B 29 56 E5 BF C6 C1 1C B8 FE
 3F B5 9F 91 C1 F8 7E 7C B5 2D A1 70 68 59 64 E6
 3F 24 0A 59 F0 CB 75 A0 3C 1C 5E DE A1 E1 F3 77
 25 C4 76 DF 17 01 0B 26 54 D9 D7 E8 53 7F 13 AA
 9B C2 DF 3C 26 D4 23 AD 51 CA 3A 25 1A 98 65 78
 DD 07 7C 15 5B 81 8E A1 EA 48 39 59 D7 F9 E3 2D
 12 17 D9 D6 DF 37 63 60 B8 68 E4 A1 53 FE DF 46
 E4 4C 3F 80 4E B5 F6 34 4D 60 39 69 6D 1A C1 DD
 9F 71 7B 4B 8C BC A1 27 F6 24 CB E6 26 28 D5 BE
 38 D2 36 12 EF 58 01 CE A0 C8 BF A6 CC 34 21 EF
 AB 4D 5B 4B 2B 05 9E C8 E9 04 7D 40 E4 3F 45 73
 AE E4 E6 34 F9 13 A3 69 6A 05 E0 C0 37 98 D3 75
 3C 40 6D 07 52 13 BF 12 7C 4C 9D 4D 90 75 F4 1F
 86 29 2F AA FB D4 37 87 C3 35 2E 99 AA 7C B5 C0
 89 93 D6 37 DE 87 79 97 AE A6 00 E5 9F 53 BE 45
 01 E9 E9 1D CE 6F 21 31 3A 30 D0 C0 23 1C D3 F5
 9D 16 0C B9 06 47 BC D7 55 B6 88 1D E1 06 94 65
 A0 A8 B1 8F 64 F5 BA 83 18 E1 E8 97 80 D6 5D 89
 41 C2 DC 71 B6 33 5B 44 A7 C8 1D 42 CD BF 1F ED
 A2 9F 5D 52 24 90 E9 5F 61 68 ED 5C E6 10 4B 6B
 97 17 F4 45 8F 22 E8 80 2D BB F9 95 15 EB 5A 35
 7B 1B 5F 5A 13 41 6D A8 D9 79 7C A9 49 FE A2 DD
 5B 21 14 75 F6 DE 82 47 42 36 E2 07 7E FD D8 ED
 8D DC E9 E4 8E 75 A3 49 63 42 12 04 A8 63 2D 54
 2F F2 E5 FC 26 DF BA 49 F6 B5 9A 37 80 D9 5C 82
 13 D9 C6 85 CD 0B ED D1 FF 5A 2C 6F EA 23 23 2B
 76 07 A4 40 5F 14 F7 16 43 85 09 8A 79 A5 29 93
 CA 77 02 F5 1C AD 5D FD 89 7C 02 DA 52 33 2F 6B
 0E 80 D0 8D 51 D7 52 1D 09 27 75 1A 30 B1 29 11
 9E 69 BC C4 73 39 A6 66 62 7A 7F D2 60 31 B9 86
 36 1B 10 C7 44 CC 50 B2 EB F5 B4 BC F3 FF 43 D3
 99 52 AF CD 23 CF 9C 42 A7 8C 28 9A 83 9C 4E 8D
 8D E0 42 99 70 CA 07 88 78 EB 92 25 BF C8 8B 76
 EC C6 98 67 F0 5E 01 F2 73 39 A5 92 02 44 5C 05
 5E 75 7A 13 06 AC 09 F9 DA 11 28 BB 11 74 88 AA
 35 82 61 3A 31 B9 EB 67 DB 76 35 EA E0 43 B8 D7
 14 B9 81 3A 89 74 F1 2C 99 53 4A AB F7 55 7A 03
 5C 15 35 15 E3 91 07 BB A7 97 72 E5 B0 73 B6 6D
 AC 6F 41 74 56 17 25 DD 3A A7 8A 50 B7 C9 14 57
 15 E0 E9 C0 5E 68 58 FD 6C 16 62 AF F4 57 47 8B
 56 7D 89 DA AF E1 4E DD D5 04 CB 20 60 F0 D4 68
 5B 9E EB 5C B6 20 A9 4F F2 5F 6C 72 FD 62 DD DD
 E6 4D 76 AA D0 8C B3 8B 5D CD 1D 91 F6 39 14 95
 3C 93 2F 52 C4 8E 39 28 6C 4C 0D 2F 85 A6 33 E8
 B6 0A AA EA DD EF C3 C2 15 22 FE 43 3B 24 EA 52
 A6 3F FE 90 02 FE 36 47 76 61 2B 3D 66 0C 91 7B
 20 31 15 6B 38 09 C9 0B CA 44 34 74 E7 C8 FF D0
 57 13 BE E1 F0 47 D6 38 7A E0 3B D4 0B 7F 7E 6B
 17 2C 03 F9 6E 4D FE FB B3 99 50 B9 2D D1 0E E4
 0D 03 16 7D 81 57 CF 29 74 51 57 56 9D B4 92 01
 98 81 79 64 AF F6 B6 93 C8 EF 46 80 28 5F 37 01
 99 AD 5F 50 0F 4D F8 D3 10 33 71 E2 20 DD D8 01
 7F 8D 8F F2 DD 63 05 BA D1 6D 74 98 EB 0E 62 AD
 C6 0F C0 BE 63 E2 9E 74 15 53 BD 5C 01 AA 35 4E
 03 E0 0B 8F DC A4 92 BC 69 CC 8F 47 7A AF 0A 55
 D2 BD EF F7 C8 FB 97 21 73 35 CF 95 A5 EC D5 04
 6D FB B2 10 62 7E F4 EB C5 20 03 3C 9B DA EC C2
 98 FC 36 2C C3 CA 27 89 F0 AC 56 9F A6 EE 99 00
 8F 99 15 9A 6C 91 8A BB FF C3 00 4C 71 F2 FB 38
 4D 1D BC 9C 9F B0 CC CD 03 CC F6 34 9B D7 79 8E
 1F 37 F0 42 D5 89 EE 74 AD DC 09 E2 48 F2 36 25
 33 32 F2 FC 54 69 BF 58 AE 28 92 1A 00 35 C6 7C
 10 19 FA 44 1F 51 FD 26 FF B9 CF B7 BF 5F FE BB
 08 17 D8 24 0D C0 B8 D4 05 A2 27 27 AA 21 08 1C
 C0 15 70 38 65 E3 17 E8 73 9C A7 BE BB 97 67 FD
 4F F8 23 31 FE 8A BF 94 DD 51 F7 8A 9D 9F EC C0
 DA 73 1D 12 8F 74 FD F3 08 14 43 A4 D0 52 BF 14
 5A 33 81 81 A4 E3 5B 95 05 79 E0 E2 A3 9A 2F 0D
 8F DA 51 F6 4B D7 A0 CC 4E 1B 8B A4 AD 36 75 14
 8D D9 F2 7F 63 7C 91 EC 84 D7 4D FF A5 26 33 B3
 BD B7 F8 8F 3C F6 D6 90 64 2B 95 33 43 84 F8 31
 D4 C8 AF 9B B7 34 1E B1 C4 43 B4 D8 67 2B A9 2C
 4B AF 00 8E BD 45 46 C4 C5 9E DE F2 3A 6E DF 18
 27 C3 49 02 3B 76 AC 32 4F 41 31 57 C3 91 54 8C
 40 E9 BE 2D A6 CF 95 A7 42 79 45 6F 37 F5 3D CE
 BA EC 21 87 7C 10 67 76 99 42 F7 65 8C 65 2A 6B
 24 CD 84 7C 7A DC 8B A7 0D 38 3F 3B 74 90 29 A8
 4C 15 E0 21 53 E7 B5 27 8F 02 49 F2 74 F5 D0 03
 34 2F 16 23 68 F5 45 8C 9F A6 C2 93 CF F3 9D 69
 AF 09 AA 7B F6 A7 AF 52 D8 ED 87 14 18 9C 17 E2
 42 98 19 C4 AF B0 29 61 65 92 D2 47 0D D4 60 1B
 5B C7 65 F9 79 47 CE FA DF E7 41 D3 49 95 4C 6C
 FF 86 F6 F5 77 40 8A 5A A4 BB 55 0E 2D 7A 80 5D
 40 22 62 AF BF 52 D1 5E 7F 09 E5 D3 83 C8 83 D6
 B7 BD 3E 8A E7 C4 2A AC 6D 57 0E 83 73 8E C0 7E
 70 E5 A7 4F BB 94 2E E1 10 7E BB 47 9C 43 40 F7
 7A 63 F2 D4 DB 7C 7F 99 CF 46 42 2D BF 07 E3 20
 8A F3 CD 4F D6 C7 E4 D7 26 C3 EB E1 C2 C2 6D A1
 62 25 33 34 43 65 A2 C5 13 A0 82 54 7E A2 45 1E
 08 2D F7 1B 99 D6 0D B3 B6 90 A5 BA 84 C2 C4 01
 64 F4 19 1D 3F 1F FF 32 69 6E 43 60 83 6B AA F3
 1C F5 98 D3 59 84 9F 34 24 51 B1 E2 CC 68 C7 30
 C6 98 6A 41 4F 57 05 DC 4C 0F 0E 19 5B 68 A6 51
 2E 82 73 FE DC 63 99 A2 92 52 B0 B8 7E CD D6 55
 A0 F2 4E B2 29 60 3C 9A CC 67 DF 8A 8A 27 C2 09
 FB 7C D4 0B 21 3C 28 AC 79 B9 95 86 7B 7B 89 9F
 A2 BE 6A 86 1F 23 96 D0 86 43 06 99 F6 DD 78 BD
 2B 35 FE B1 A7 D5 97 47 59 C8 1A ED 26 E2 93 6C
 8C 24 A7 52 95 EE 29 74 6C 01 5A CE 9E 58 4F 7F
 13 31 67 38 0E 7B 0E E8 65 96 E8 12 5B 62 96 E2
 09 4A 0B 19 65 43 D2 43 2F 7C CD C6 39 CC A9 4E
 B7 1B FE B7 E9 A2 61 03 A5 8C 3F 2C 2A 75 B3 E1
 A4 B8 E9 69 D3 0E 47 52 60 A0 65 55 6D 99 43 99
 B9 40 EA AF 10 B8 62 47 4F 5E 08 C2 06 FC BA 53
 35 E2 10 CC 5E E6 12 9B 80 0D 68 E2 74 A0 EB 62
 09 A1 25 96 E5 3E 4F 1A 70 58 DE 8B D9 BD A5 96
 60 64 9F 1E 85 CE 29 F5 EA 67 24 A4 DD 2A AE D0
 80 F3 83 41 0B 20 22 5E BB 19 01 7D 4D 46 03 AB
 B7 CD A0 3B 50 73 39 2A 85 76 34 AE 39 E1 ED 44
 2D 7B 7A 37 FB A0 7E A9 7E 05 66 73 DD 04 D2 34
 AD 57 0A 51 0F E1 31 6E C5 B3 B7 75 8F 69 49 65
 10 0C 38 6E 6E FE 89 FA C8 96 AF 2A 0C 07 33 68
 47 E6 8E 56 23 37 90 DC 48 E1 A7 A5 C1 33 58 35
 92 B2 E9 0F 90 57 75 E6 95 92 7B 6F 48 94 E5 4C
 6F D1 CE 4B 5F B1 85 E4 46 BA 3E 61 18 A3 CA 2C
 61 03 AE E1 BB 7F 39 8D A6 B0 0B BE F9 72 FB D8
 FE 0D E1 F6 C7 9A 8B 0E 51 B3 84 D2 85 19 1A 0D
 D5 47 68 38 13 C9 0A 6F 26 0D B4 42 FE 00 62 C8
 3E 21 2A EA 36 6D 06 45 2B 41 90 33 79 B6 AA D3
 08 41 C8 A6 96 EE 18 1C AC 26 2D 7B E5 DE 86 D0
 5E C4 E3 11 4F 7B 5F F9 B6 8C FF 64 9F E0 25 92
 84 34 7B 0F F4 C0 AE 90 D5 52 3A D3 F9 FF 62 8D
 F2 08 1F 5F E0 4D A0 10 76 BA 1C EC 40 25 9F 21
 FB 90 49 6D D7 6C 2B 46 53 77 13 F0 24 84 62 4B
 2C 53 30 9B 80 B8 A4 6E 36 FA B6 FB BF 71 D9 41
 B3 02 98 51 B1 7B 22 67 2A E0 89 BC 3F 18 7C 42
 B5 50 66 CC 1F CE 6B BB C8 B7 B9 62 E6 F4 BF D5
 B7 4B 72 78 E5 3F AE E0 B6 1F 3D 2E DC A7 62 CB
 E7 0A 86 93 30 D7 D9 DA FB 0C 5C 04 46 6F 26 F0
 10 EB 40 9C 18 C1 7E 7D 7E A0 4F 41 1E EF F4 0B
 AF 8E 8D A4 C1 4A 93 63 A0 C1 8F 39 DD 17 B9 AB
 6B 49 57 1A 3D 9B 6D 13 D0 4A 0C 9E DE 38 A3 FA
 C5 98 75 CB 84 B5 11 F3 30 73 05 8D 83 43 DF DF
 C1 F8 53 39 EA A3 58 C5 F7 E8 3F C2 F7 5C 06 0C
 46 0A B7 1F 3F D5 8A A0 43 61 E5 FC EB 63 E8 5F
 3E 4D 4D E5 FD 2C EF 99 F7 12 99 10 B2 DF A7 B6
 B6 03 B2 C5 03 B3 D7 21 C5 AA 68 3F 3F BF D9 13
 83 6D 91 7F 19 78 EC CA E7 49 1B A9 3F 22 84 79
 C9 E7 A0 68 84 43 FB 7E BB 05 86 EC 41 61 9C 47
 3B A7 AB B7 A0 5E BA B1 5C 06 B5 69 70 9A 68 33
 AC 7D 9E 13 EC BF 18 D6 2E D2 62 71 47 C7 F2 7B
 41 13 AB D0 4B 7E 09 87 BD F6 44 82 43 66 03 7F
 A4 2A 69 40 E6 32 54 59 B0 B9 DE 28 D2 18 28 32
 44 93 C8 25 E9 D0 61 29 82 4F 93 62 EC F0 DA FD
 F2 78 2F 01 D6 8F AB 6D B8 E6 DB B0 B8 0B 89 10
 DA A3 F8 7B 19 E1 9A 02 3D C0 EA C5 F7 8D 37 08
 15 09 E9 04 56 A4 EB 2E 01 94 40 F8 3D 97 14 CC
 D1 F4 0B 3C 3B 69 7A FB 86 92 CC 26 3C F6 CF 7E
 72 D6 D4 97 17 E1 5B F2 91 14 80 D3 C7 C3 67 E6
 D1 E8 B5 89 DA 08 54 4A 9F F5 7F EF 2B C2 57 68
 43 1C F6 FD 1F FB 70 47 F6 A1 9D 5B 41 1C F9 55
 3A AA F0 0F 7B 35 33 AF 10 06 E1 5F CD 52 74 12
 E8 EC 0C 15 38 CD D4 E6 59 CB 0F 6C F8 99 D7 02
 81 62 3F 1C 59 22 44 1E 37 9F 1C A6 29 B5 B6 BF
 96 8C 0B 69 6F 76 FC 57 64 33 95 C5 A4 BF 49 20
 20 75 68 E6 8A C7 E3 A5 45 82 C2 72 27 2F 6C 64
 0E 52 77 25 19 AF 45 4D 4E 55 9E 02 E2 13 CC 1A
 14 F0 F5 86 4E CB AB EE 49 0C 6F F1 43 B1 FC 3C
 78 89 8A 15 07 D8 4A B3 4F D7 39 BB B2 0B EB 96
 37 35 40 61 DC A5 04 41 43 20 2D 84 26 5A 4C 7D
 98 47 3B 06 B2 03 40 42 70 E4 23 81 F3 4B F4 40
 07 8C 39 09 3C 9E 5D 01 04 C1 8F 74 DB EE 06 0B
 46 48 0D 44 70 46 61 A5 CD F9 73 15 C3 37 3F 33
 DE 9C B6 32 4B 58 B9 40 83 56 FE C5 B5 6B 65 DE
 C4 5D 34 23 7B 67 E3 9C 65 AD 79 A2 C0 4D D7 DF
 76 84 17 4D 20 00 E2 77 91 D5 90 22 3B CD 94 07
 83 AA 38 0A 65 8A 56 65 C6 E8 B3 2C 94 0E 37 19
 BD 90 37 D9 25 AE 51 2E 69 DB 3B 43 6E C0 72 A4
 23 8D B0 E1 9D 0D 37 AE 66 64 FA E8 C6 78 51 3B
 0D BF 51 4B 1D C0 C3 98 79 54 74 83 17 9C 77 A3
 EA BA C6 C6 EF 31 6C CB EF D8 CD F1 70 E6 60 47
 A7 2E B6 87 A2 E2 71 66 AE 21 0A DE 9D 09 7C F0
 B9 E9 9B 7F D6 2C 18 69 84 72 EE A8 1D 88 63 41
 23 90 BD 0E B3 50 5C 6D BB 8E 91 14 49 45 13 1C
 2C 22 80 08 DC 35 44 77 BF C5 6D 3B 13 CF A6 2A
 3C 5D C2 32 87 17 17 A4 28 4A 7B F9 C5 EB A2 0E
 F1 62 7B 47 1A AA 1C 51 F7 D6 89 C7 87 AF 0A 05
 7C B9 AF D4 C9 78 8E 1A 2C 38 75 8B 34 CA AA C6
 0B BA 9E A2 9B 9D 9C 8B 10 4F 5E D6 36 92 54 82
 35 7D 40 11 8F B3 E6 6B 8B B6 9A 53 B5 0E A2 26
 79 E3 1A 6F 1A 78 69 3A 0D A6 42 69 3D D4 0F A7
 DC 9D 65 5D 97 CA 68 0C 13 56 DA ED CE BD 54 55
 70 78 C7 E9 42 C1 5E E0 25 47 C1 74 BA 87 DB FB
 7C CE 44 D2 E7 86 83 50 64 61 66 63 48 74 00 A2
 16 8C 56 93 79 57 E7 CA 8D A5 D0 56 49 EB A1 E3
 54 A1 7C 16 1E BA B3 AA 02 72 F9 69 C3 D6 5D 41
 BF 6C E1 5F 3B 3D 60 BC C2 31 29 EA BD FD 29 19
 78 F3 75 BD E4 17 C3 D6 47 3C B4 39 56 0A 41 9A
 24 FD 83 7F A5 85 F2 9F FD 02 7C B4 FB 3D 9C 0A
 3F 0D 93 B9 D3 50 43 B3 10 69 9F AC 3F 03 3E E8
 B7 FF 4A 56 51 FE D0 E7 BC 27 C2 A0 91 F2 C9 DC
 C7 B6 51 74 49 2C BB A1 E3 61 ED 59 0C 9B 6F A7
 F9 5B A7 EC ED 6F F2 87 60 50 D7 44 2E 1F C7 41
 2A 43 5F FA A6 9D 8C 0E 55 94 59 CD 15 F4 D7 3E
 40 E3 DD 7D FD 86 B6 FF 42 0C 4A B6 2B 08 19 3C
 28 CE 06 A9 58 92 59 E3 D1 40 25 29 B7 2F 89 76
 F1 27 E8 CC 1C CF D8 D5 A8 97 78 8B DE D5 FF B4
 1E 07 C4 AC 56 0C 0F 96 5B CA C1 FD B5 6F 4A 63
 E7 EC 58 90 19 F8 BC D4 8B 96 C2 17 4D 9E 0A CB
 4D 6B 84 33 66 F7 6E 68 9F 97 F5 68 59 92 CA 47
 41 9C 1F E5 C8 27 E5 12 F1 78 6E DB F7 91 1A E3
 E6 55 ED 40 14 97 1E CF 2B FD D8 89 DD C7 2E 55
 F4 29 42 D6 D4 69 47 59 74 E9 5A 39 9F 2E 66 09
 E7 30 44 7B 33 DC 7A 7F 36 38 05 7A 48 69 E1 09
 0D 94 C2 80 4F F6 3A AE C9 05 A5 E2 10 E2 2D 3F
 4E 80 A9 B9 D3 1C 5B 59 E3 0E EC 0D FC 17 F5 F9
 3D 43 1B 69 A5 64 F9 FD 66 90 E8 09 32 C8 8B D2
 C7 47 AD 82 86 A0 62 B5 73 E1 09 85 F4 3A 6A BB
 04 87 B2 F0 D5 29 37 49 EC 23 0A 6E DF 0A 6D 5F
 F4 0D E8 77 AF AA 2E B8 D6 A6 13 C0 CC 8D 2C 70
 2E C9 B5 69 DF 20 E4 9D B8 4C FD 92 FC 71 2D 4D
 92 CF 47 28 14 6A ED 65 E9 FA D4 1D D3 81 C2 5C
 B4 88 29 49 D8 06 B9 46 A1 93 45 ED 94 0C A9 D1
 6C A4 5C C1 9C 4F 01 F5 A2 88 44 83 C3 0A E2 0A
 57 01 38 5E D9 30 A7 1B EF 42 B9 74 F0 80 65 7C
 00 7D 9B F4 E1 58 7E EF A1 1E F9 E7 9F 98 C0 48
 AA 37 11 B7 EB C0 44 2C 4B C1 52 7E 98 77 9F FC
 36 83 B4 D9 E1 FE 2F 0C 0B 40 17 FE 5A 96 A5 0C
 D6 50 AD 72 37 E6 96 F3 C7 B8 17 63 06 60 C9 92
 49 01 B7 BD 96 F7 5C 6F E7 42 9C 79 98 03 A5 C7
 B6 85 08 28 49 68 BA 8D 0B 3E C7 8B DE 1F D2 35
 E8 04 BF 09 A2 13 C1 FB 80 05 D3 FC 20 0B 78 55
 73 40 B4 F0 F7 07 2B B2 40 E2 2C 4B D5 03 B7 40
 48 1C 25 D0 2E BC 09 0F B1 4B A1 03 0B 81 50 6D
 B2 5C 31 BE 0F 78 00 D8 73 FD 2F 61 C5 22 BE 91
 E8 B4 1D B7 48 15 7D 3A A2 99 50 A8 78 41 12 AF
 BC 06 1A 64 F3 E2 48 99 E8 6F 91 F9 F5 03 4B 01
 CB 60 D9 CC 42 24 4A 83 39 91 10 AA 65 01 52 5D
 04 46 10 F7 97 A9 48 F3 C9 27 CE 6F 33 54 54 A9
 24 04 20 5E D3 0E 10 39 DA BF F8 9C B5 2C 85 B7
 BE 75 5D 92 B9 BA C5 03 12 78 88 08 E4 57 D3 C6
 C5 38 45 6A 3C A2 26 0C 85 A0 D2 3C D4 EA CA F0
 E4 E2 2B 88 99 11 C1 6A CB 7F F4 36 89 3F E7 50
 5A FA CE 62 52 D6 6C D8 7B 49 99 52 2E 8E 1C B5
 AA 01 EF FD 4D 77 3F CB C0 5B 5A 08 7C A0 B6 2B
 AA C3 2D 2D 99 4A 44 7A 78 3A 47 A8 F5 F7 F4 D4
 F5 7D B1 FB 29 E4 CD 95 DF 4E 09 DB 35 40 F3 84
 BC 56 B4 85 7D C2 D3 0E 98 C8 CC 7A 71 88 0E C4
 83 57 93 F1 64 C4 72 0F 1D C0 3A 26 E4 36 6F 0C
 45 01 5E 30 71 D2 CB 3E 9B D5 3E 5F BC F4 47 4E
 5B B3 D5 86 1A 95 82 E5 DD C9 8E F1 31 AC 79 DD
 9F 09 DA 00 86 3A 26 C5 17 76 63 2E 99 C7 0C 95
 2E 51 C5 10 4A 77 42 1D 9B EE 67 F0 C2 86 32 54
 79 CF 3D C4 21 B1 AE 35 4C FF 12 2B 45 DE E7 92
 92 3E 6D 0A 39 A9 5C 14 4B 8D DC 24 73 11 6D AB
 D4 EE DF 9F 0F 83 B6 84 FA BE AB B7 39 93 9F F0
 6E 5C 6B EA 06 A3 AE 29 81 47 26 62 2F D6 A1 82
 73 90 22 0A 4D 14 0D 27 21 41 EE 0E 1D 25 28 C1
 92 84 C0 E7 85 93 21 FB E1 85 F4 AB DA 03 F6 14
 A2 C6 C0 0E 6F 37 07 33 28 F1 6F 11 5E 76 0C E3
 BE 9C CB 10 CD D9 E3 40 D5 CA 62 BF 1A DB 31 AE
 24 81 3D 21 E5 5A 38 CC DF 3B B0 C0 0F C5 AF D8
 7E 7C 60 1B 0F AE 5F 6C A9 BA E6 C0 B8 86 E9 F8
 FA 6B FE 79 9E 1F 1C E6 79 2D 33 46 4C E5 61 D1
 96 B2 20 18 5D 63 C1 F8 32 B1 65 EA 5F 82 7B 0D
 D4 72 1D 5E 1B 71 00 84 A5 EE D6 68 8B 02 14 80
 A8 AA 3E 0B AA F6 6A E2 35 CD D5 F6 25 8A C1 1C
 82 8F 31 1F 50 8A B8 46 DB 0A AC 3E 3E 9A E9 FF
 1B 75 A5 1E 81 47 1B 4B 00 E8 0A 08 E2 C2 B5 46
 ED 5C 65 CB 26 13 96 0D E6 B5 9E F6 71 3E 46 8C
 90 42 20 64 23 38 E0 5A AA 69 0F 39 B4 8B 31 10
 65 14 A1 BF 4A C0 87 70 38 06 D1 EA 55 6C D0 EA
 44 50 A0 F4 DE 20 1C 00 8F ED 21 F1 AB 47 DA BC
 8C 96 CC 7A 4D 7A 24 CA 67 4E 2B B9 CC F0 C7 90
 AB 7D AB D1 98 4D 5E AE 88 54 0E 88 81 53 BC E7
 8C F3 1E EA EF C1 22 06 DB 5D 5B BB AD 5B E8 40
 94 14 6C 37 53 60 AA 18 08 FE 00 7D F9 DF D6 DC
 81 41 FB 15 A0 B2 41 33 C0 4B FE BC 73 4C 3A 0E
 F6 89 01 71 1F 60 C6 34 B4 A9 B4 36 2F C8 41 56
 24 C6 B7 1D D1 47 80 7F 23 95 29 19 B4 28 0A 82
 11 C9 63 1D 39 80 7B 30 63 2B 47 EA BA 03 F9 89
 38 EC 43 38 A7 14 CF 47 96 0F 79 D9 3B 1C B3 6E
 01 36 CE 33 56 E1 D3 FE 16 24 D8 B9 14 E5 75 25
 C2 82 A2 76 E3 0C FC D1 9A 98 23 A6 BE 49 42 9C
 AA 89 FB 81 DC C3 EE 6D E2 70 EC FF 30 38 FD EB
 97 6F 51 04 E4 CD D1 44 BC 6E AC 3B D6 5D A2 D0
 69 A7 87 80 A5 E9 61 46 33 C1 83 20 3E B0 E1 D4
 70 35 EA 32 1E A2 74 3A B4 5A 47 DE 17 5A 44 84
 9A F4 2D 6E BF 0D 2B E3 0F 5B FE A5 AD EA AD 57
 2A F5 D9 33 92 D3 1D 91 70 5D 0D 68 29 09 6B 00
 B9 3C 9E 3B 20 AA E9 5C D9 C1 96 FC 08 00 90 96
 29 03 DC 7E DC EE 60 56 FC 9E 30 28 E6 8C DB 45
 D2 02 35 78 D7 FD BB DB FA 4A F6 0F 30 DA 21 88
 9B DB 88 49 0B A6 70 30 BC 84 06 02 70 9C 47 9C
 AB A7 C8 69 BF B1 1B 97 7C AD A5 B2 1E 24 29 3A
 9C 15 8A 45 FB 5B 60 54 BF FA 4B 71 B4 63 22 3D
 7C 36 B5 32 20 56 E5 0B 18 F2 61 79 74 BB 17 90
 C4 C7 53 B9 00 D6 C0 C9 5B A5 F3 85 C4 9B 08 94
 5F 7A A6 3D E6 14 73 7F BB CC 6F B7 85 D2 0A CC
 59 06 BF 58 D6 CA C2 D6 E0 55 98 97 7B 2F 76 28
 D7 85 7A D8 99 5F 5D 5D A7 61 91 B8 80 92 D5 16
 4B 21 06 F6 77 F9 5D 5E 8F E0 36 95 40 C6 32 12
 8B E7 ED 90 22 FB E5 50 F5 A8 DB 77 12 CD B3 F9
 A7 FB CD 57 B5 74 C4 01 CE C5 A1 67 20 7F B9 10
 2C EB D6 E5 42 7A F9 79 E9 D1 DF 4E 81 C6 56 95
 F1 D5 DC 45 AF FA B5 E2 4F DA 8B 4F F5 E6 BA B0
 09 0F 29 86 66 A2 07 10 78 90 F3 DF 92 83 09 4A
 FB EC 20 08 E6 E8 E9 95 39 57 1A 75 ED 35 9A 8A
 9A 03 92 92 AA 9B 99 80 81 0C CE 5B 84 9C D8 F2
 01 5D 42 12 57 23 FB 83 26 4C AB 68 66 9E 9E 3F
 3C 6F 02 8D 29 4B 0B B2 6D 00 14 B7 13 B0 5D C8
 13 E5 CF 5C 02 D1 2C DB B6 22 B9 6B 7A BE DF 94
 08 A2 E9 D1 B1 1F 1C 36 0A 42 7E D6 D7 C2 10 41
 7B C5 BF B2 CB 71 63 AD D3 DA A2 87 C6 BD 95 6A
 79 F2 75 F9 5C 96 46 7F D8 FB 5C BD 7C C5 BA 23
 B3 21 91 74 2A D1 69 B2 F7 3B 73 32 4C F4 C5 F1
 B9 AD 20 E2 9C F9 A8 D5 08 F4 E9 D6 E7 80 61 5C
 7E C3 31 1C C8 34 31 4E 9F 12 E9 B5 52 6C 90 BB
 8F 77 A5 81 54 A0 BB E4 3A 87 FC 0A 97 71 A7 D0
 67 4A 4A A8 2D 81 5B 6B 3B FF 00 06 63 E3 B1 69
 47 A1 D2 6E 40 9D EB 56 CF C0 B9 60 C3 D7 FE 0F
 B2 0F D6 15 59 A1 34 9D DD 2E 90 94 BE AE D1 89
 ED FB 4B 00 07 2A B0 92 18 66 3F 2F A3 29 F5 A6
 79 80 F3 46 4A 8E 33 5B EC 84 42 A7 38 B7 69 27
 5E 33 ED AF 7C 10 E7 AE C1 14 E2 7C 29 C7 21 D9
 0E 95 8D 44 DC 35 5E 6D 2A 48 4C F6 27 68 D5 96
 2F 0D 24 3B A2 49 37 94 A4 F1 C7 60 25 DF 3B B7
 76 4A 1F 2F 0E 31 36 35 00 73 17 31 5C 8D 7E 77
 43 6F DB 09 3C 75 FF C8 94 D5 5E 6D 1A 88 34 7C
 8F 21 C1 6C C6 BE A7 3C 48 F2 60 E5 C7 B7 FB 42
 D1 E7 FD DE 80 66 0C 13 89 95 A4 81 83 37 A4 47
 34 20 19 46 4B DB 1C FB D4 73 D4 40 6F 3A B5 5F
 AD 36 55 6A 8C 51 EB 6C 29 AC 63 C3 73 6C B9 7F
 4A 8B AF 41 73 9E 27 20 8B 4E B7 D2 AB 61 20 AB
 38 04 62 C3 A2 AF 41 D1 A2 DC 8C E7 6F 35 8E E2
 DF 23 38 FE 89 64 47 2F 64 D9 68 BE 14 E2 D7 C0
 AF F5 07 16 A0 1D 3A 5F 7C 90 3D 53 E2 AE 36 72
 4E 97 58 EC 7D A0 90 D8 C6 C1 49 48 D2 8D 8F 1C
 10 98 2B 51 D8 B6 2D 0C 9E EA F1 FE 61 5A CB 3C
 54 8E 06 B7 93 7F 86 61 79 8A 05 3C 5A F2 DE DC
 B1 F8 14 F4 A1 06 C9 1F 69 34 56 12 B3 0D FD 60
 D4 98 6D E3 9A 25 67 A7 4D EE BE 16 21 C6 8D FD
 AE 01 09 C4 8D 6A B3 AE 53 FE B7 7F 33 C8 2C 35
 98 8C F2 54 1E 12 72 7B A8 28 17 23 78 C0 83 9D
 36 F9 20 6D BF F4 FC F1 2A C8 6B F0 19 CA 35 2E
 6E 67 42 56 B9 44 88 6C C5 64 A3 03 31 3E 58 C0
 5D 87 61 7A D9 CC ED 23 13 85 2D 25 D3 39 FF 4B
 D7 AB DE B5 A0 84 51 82 F1 0A 13 9A 30 3A 83 89
 75 8A D1 82 34 64 EA BF 47 BC E1 9E 48 D7 33 00
 52 F7 2B 51 72 26 7E 32 C2 66 07 DA B1 DF 25 1D
 FA 82 63 43 11 AB 3E 5B F8 42 86 38 6A 35 B4 1C
 AD D6 5B 03 EE 3D EA 6F 23 B2 96 40 B2 78 51 6D
 EA 92 32 CD EB 02 5C 53 60 37 78 3D B7 8B D3 0F
 DD 11 40 6A 1D 80 B2 CC A2 8D 71 83 55 F7 00 F2
 32 41 9A 3D 59 B7 CF 70 C6 A8 40 11 42 A4 1C 90
 78 CE 1B 8B 8B F8 EE E9 43 D5 4C FD 9D E5 70 93
 84 2E B5 3F E6 BF 89 2F 08 7F 02 D6 B6 8E EC 3D
 66 3D AC 26 6D D6 58 20 90 74 39 92 2F BC CA 02
 D1 68 29 67 29 08 73 AC EF 3B 95 AD E3 6D 3B E3
 C2 87 D0 E1 0D 2C 49 DC 94 E6 AC 46 3C 7D A0 E9
 3B 13 40 52 EF BE 15 3F 96 88 B5 ED 15 B8 6B 40
 AE 6E AD 17 29 ED 6F BF ED 95 FA 4C 51 05 54 95
 CE AF 1F 6F 62 60 F1 63 A5 39 EF AF 91 62 5E F2
 5F B7 F4 10 63 D5 16 D4 6B 52 5C 3C F0 23 C5 38
 B7 01 B2 AF 5F 06 E5 F7 0D CF 18 92 F5 46 25 00
 6B D0 68 75 AA 57 CF B6 EF 64 EE 72 8E ED EF F9
 3C 22 10 59 1C 6A 7B 37 37 08 4C 44 7A EA 1A E1
 80 7E 43 31 73 A9 D2 1A 1A E6 02 84 A5 15 F8 7D
 B9 B9 5C F8 AE 1A 7D 91 90 6F 04 1B 1A 72 A7 AD
 14 84 E3 66 46 3F 71 57 CB 32 C2 D0 5A B1 71 1F
 DF C3 91 82 1F CE C2 9A 41 37 71 0F 33 FC 5A 46
 B0 B6 0C FD 08 A4 C7 77 11 0E D2 42 1C B4 C5 20
 8F 8D 87 94 0A 89 D7 46 BD DF 2A 76 3F F0 E6 4E
 7D 39 9A 82 C2 0C 1D 4C 1A 04 FE 46 D7 E5 FD DB
 2C E9 D7 98 10 3D 82 C0 DE 34 35 8B 7E 22 CD A3
 B9 CF D2 C4 C0 DC C1 7B D6 27 35 D6 B4 62 2E 42
 D2 2B E8 A6 A0 6A CD FC FE F4 9F 5E 2A 81 A2 8A
 29 68 A3 32 09 AD 38 BF 2D 4D F4 18 A8 5B 8A 4E
 76 82 E7 5C 39 FB 54 43 8C 54 FD D3 EA 28 B4 37
 DA DA 50 B1 99 6D 2D 37 B7 36 07 EB 2E A4 7F 17
 50 54 52 D9 F2 0F 75 AE 34 30 8E E0 01 D9 6D 75
 26 4A 3D 42 79 16 B1 FD 7E B2 C5 AC 14 DA FB 13
 A9 F2 1C A9 2A E9 64 AC DB 5A 19 8C C3 4B A5 19
 6D 99 04 82 19 1E 5D 00 09 AA 29 9B 26 3F 17 5C
 A1 41 F0 65 F8 A8 18 D8 A0 70 1F A5 6F 86 C5 B9
 4C 70 6E FD 22 F4 F9 2E 3E 1F BE F5 B1 32 FC 23
 E3 3E EB 06 C1 F4 42 AE 9E 02 86 8A DD A6 6E 91
 2E D8 88 4C 1D F7 FE C0 DC 17 50 E4 7A 5D 26 67
 71 45 E2 85 BC 86 C4 1D 31 BE 11 91 61 5C 92 51
 C8 9B 5B 99 06 43 47 6C FE D9 BB A7 DD 5E 9C A9
 43 41 46 95 A3 C3 99 52 FC 3E 29 89 86 03 C0 25
 9C 3D D4 A2 D0 CA 12 5F E7 71 F9 E5 04 1F B9 5E
 8B A3 88 47 4B 3A 50 24 7C CA 37 D1 DC AA B0 91
 FC A2 6E B6 8D BB 76 FD 26 DE 51 E3 AE 87 7A 81
 63 A3 6C 13 33 2B 71 B8 B4 74 DA E0 6E 3D 97 77
 36 96 E8 11 BE 95 D4 32 B4 0C E4 A6 AE 43 9B AC
 FC D7 56 9C 7B 14 35 2A CD E9 28 9B 98 03 1C 3E
 75 6D C0 B1 9B 47 F0 C1 CE B2 24 1D 70 77 98 D2
 54 00 80 E0 25 7B B6 08 82 68 4D A5 5C 1D 16 30
 7F 5C 25 BA F7 D1 19 E5 80 38 5C 77 EE D1 AA 79
 31 F3 77 5C 84 A4 BA 83 DE 92 F2 7B A4 2A 59 ED
 35 18 F9 9D 16 A5 2D B1 1A FD 3F 90 88 F2 FD D1
 FB 15 AC 6F 95 9B 5E FA 22 5F 2C B9 B4 0E 1F 49
 BF 4F 6B 7F 19 A0 DC A2 6D D8 C3 DE FB 45 64 64
 A6 FB 0C 1A D6 4F D9 F2 03 D2 71 FF 39 2B 79 7E
 0C 8A DD B3 7E 40 DB 3F 44 02 87 F7 DA 2D E5 AC
 92 93 37 4F 3E CA 0E CE FF 88 1A E4 2C F0 0B 6C
 75 BA F9 90 97 2F 20 0E 6E 93 5D 42 05 71 BA AC
 46 D6 03 D8 15 56 8C AC 64 E7 35 A2 9B 01 CC 94
 3E E0 CD 10 DC E7 D5 C0 2A 75 F5 86 7D E8 A9 28
 F8 B1 22 66 8E 62 D7 87 06 AD 18 62 74 9A 53 72
 CF 89 CA 7F F8 89 D3 80 77 E5 AB 03 12 DA 05 E3
 F3 42 E2 8A A4 20 36 FF A6 C4 9A 76 D3 52 73 3A
 E3 74 66 48 16 EA 5D 84 8B 8F D7 74 8A BC E4 97
 1E F6 E0 F1 9F CA 84 40 37 F6 17 47 4F 89 F1 3A
 CF 76 78 89 D3 DF DC CA 26 DD E4 35 0F 10 B7 50
 E9 85 E0 3C 22 00 E6 D7 22 9C AA 5A 95 8E 9A CE
 C9 3D 08 19 E1 F8 CE C7 77 CB B5 1A 86 71 C7 17
 D4 F1 79 0C E5 2D 23 95 07 B6 DE D5 81 C5 2B 25
 7A 84 47 1D 12 7F 3F 58 48 7E EA 6D D0 CA DD FF
 E7 26 7B D1 DD A7 8D 45 2E 47 D1 41 32 E3 B1 41
 6A 43 DE 65 3A 35 44 40 2B 57 08 98 25 6E A1 13
 24 29 80 04 56 13 B5 7D 7C 5A 5E 83 CC 94 4C 59
 FA FC 81 D4 BB 90 2A 72 77 EB 13 53 5D 24 9B DD
 C8 10 EF F0 8B 77 6B 89 BD 48 44 A5 B2 F8 6B 96
 72 8E C3 9D BD CF D6 B9 73 5B EC 28 95 42 1D 4D
 A6 2B A9 E6 F2 AB C7 CC BD 39 68 94 FE E2 7E DB
 28 69 63 0B 27 56 65 FB B7 DA 15 74 11 BA DB 7F
 C8 D5 A9 54 9E 6C 65 3F 5F B9 E9 A3 66 29 05 4A
 D0 69 C1 86 E9 01 2C C4 1B 27 A7 51 33 D7 ED 1C
 58 CF CC 5F 8F 42 53 D6 08 59 FC C9 4E 71 69 DC
 79 40 71 F3 74 74 8A 90 29 57 7E CA 7D B6 F6 F7
 57 A4 AE 5A 3E F9 27 A8 78 70 28 BD A9 1C 36 1E
 F3 8B 0F 33 33 89 EE CB BF B4 2D AA EC 4C 00 57
 8A 84 38 55 85 A6 FE 58 68 F7 80 66 66 A3 56 73
 02 AA DB FB 62 4D 6A 49 81 37 4B 86 CD 69 09 D7
 0F 16 EA D7 2E E6 6A 22 C0 21 E3 BE 66 55 75 3F
 84 53 37 46 E2 5F 39 DB F9 2D 0C 0E F9 C0 CC 38
 5C A4 47 ED 2B 10 AF AD 34 6A 48 E7 87 52 4F 19
 61 F9 98 EA E7 2B 94 9A 52 CA 00 0F EF FF 9B 8D
 CD A8 91 73 31 C9 2C DE 5C A6 33 79 79 08 F4 6A
 72 56 8C 93 45 D1 CA 29 7E 50 E2 B3 19 3A 31 C8
 AB DD 1B E9 01 62 81 0F 02 46 F1 9E D5 83 B8 54
 CD EF 63 19 B0 C6 19 7D 0E 4F B2 D7 CB 51 97 8C
 5D D8 FD 16 E6 CF B1 FC 6C CE E1 EA 12 AB 50 0C
 28 A3 D0 77 CF E6 21 98 A3 96 1F D1 34 30 5E EE
 56 3C D3 2F DD 05 2B EE 84 59 CE 4C 96 A4 49 2E
 B9 54 28 C2 40 2C DF CB 00 AA 5A D7 EF E2 58 0D
 1F D4 59 6C B0 02 0D 89 37 94 C9 85 AE BA 6C 08
 28 5D 25 10 B2 FB 43 E6 BD FF 3F 8A 67 BA 8D 7E
 15 CE 40 68 D0 DE 93 1D 4E 23 25 D3 65 68 35 C5
 48 9C 56 8E D9 72 FB 2C B1 CF F0 5C 34 93 F1 B3
 27 EE CE 5D C2 FF 93 6E 29 92 1C 9D E4 B3 F0 0B
 99 72 DA 26 9F CD 7D 55 18 38 24 21 DD EE BF 37
 84 4B 60 91 AF 04 0E 65 80 11 78 1D 83 E5 73 84
 15 9B B3 D1 85 7E 7C 9D A1 D6 C7 BC DF 9A 81 3F
 DC F5 4E 6D ED 35 DE 58 F9 02 92 EF 01 C5 50 20
 32 BD 22 00 AB 0F 55 D8 BC A1 B4 0D E8 72 7E 6F
 98 98 6D 41 80 17 9D 69 25 20 FC 0A 99 4C 58 E9
 A0 57 78 7E 9A 77 15 BB 09 C6 24 8C 6E 82 0A 6A
 C4 24 99 04 A0 E8 F7 5A 15 AD E1 91 8E FC E4 69
 46 6B DD 4E 36 BA FB 0B 42 76 58 3F DD FF 34 4D
 69 D4 A5 4F 26 96 73 CC 43 63 C7 A6 34 6B B2 80
 06 F9 37 CE B5 4A E7 91 2A 1A B2 17 6E 5D 29 15
 11 40 41 27 90 9D 9F 2C E9 F0 5C 17 BF 4E 4F 2C
 70 2D FA FA 84 F1 C1 02 ED EE 10 63 CC 8C BB 73
 9E 14 EF 07 95 2E 46 CB B7 52 D9 6C 1D 12 7A 2A
 2A 9F A4 4F 20 9C 59 18 63 68 9A 18 E6 A5 C5 F6
 87 DB CC 9A F7 5E B3 DD 1D 08 D1 2A E4 0B 91 B9
 D3 0A DA A3 54 4B E2 28 B6 7A 6B C1 AE CC 3A 65
 B0 5A AE 25 61 78 D3 34 16 00 22 3F 64 B8 09 82
 1B 05 AC B9 1E 5E 54 C5 E9 54 BB 36 C7 88 91 1C
 7D C2 3C 7D 5F A7 2E 57 4B C8 48 A3 F3 08 77 B5
 99 10 86 CC 57 BC 7B B2 11 B8 FB 60 4F CF 94 4C
 AF 64 AB 8F 71 44 91 CE BD 61 DA 2D E1 51 A9 9E
 97 98 80 6D 4D F7 C3 AA 79 FA B5 A1 38 FE CC 63
 99 97 5D DA F1 53 28 9B 9A DD 84 F8 CD FE 32 51
 C2 AD C0 D1 08 EE 7D 27 72 09 AF FD B6 21 D5 27
 F0 86 D3 13 E3 21 CF 98 C6 29 40 80 BE 17 B0 67
 EB B9 9A 89 8F 6B 2B 30 9E A8 89 76 75 CF 7B 37
 31 2E 25 94 02 E6 81 82 59 A1 9E 00 66 34 F3 FB
 84 74 EF ED E9 B2 99 B1 39 C1 CA AC 82 2A 37 9E
 19 0F BF 9E 8C BF CF 5E 8F 2A 55 22 59 DA 0B 34
 DA BE 28 E6 59 9B 0E 9E BF 70 C5 3E 0C A2 8F 88
 DA 54 61 E4 2A B6 A9 44 AF 13 26 18 8D 17 78 73
 D3 FF 97 F8 59 8E B6 AD 2A 88 DC 23 95 99 4D C8
 A3 6A E6 1C 4B 39 0B 6D 5F AE 07 2B 02 A7 C2 F5
 5F 90 17 5B 0F 80 96 47 26 4B 89 2D B9 A5 A2 73
 DD 05 D0 F3 82 8C E8 95 D2 44 EB 24 90 00 4A 4C
 2C F0 E0 4C F3 A5 8B 03 4D 47 19 CE 7D D2 BF 55
 2E 88 0D 6E 62 D1 ED 7D C2 EF 9D FF 4A 54 5D 32
 78 6D B7 A2 33 85 0E 56 CF 6E E5 87 DB 06 6E 7C
 3F BD 54 1C 63 4C 85 FF 9F 69 52 6B 86 AE 51 88
 A9 C0 BD F3 F8 08 00 4C E4 3D 4F CF 22 62 BA 76
 E2 22 79 85 56 6B 9A 22 93 1B 4A 5C AE CD 0B E6
 41 4B 31 2C CC D9 C0 89 FB ED D8 86 2E E1 64 BD
 A5 8D A3 45 31 3E 2E DD 12 B4 90 1B E4 7F 9C 46
 47 38 C3 B6 B8 7E 20 62 90 EF D9 84 3F 83 2C 09
 4A 40 3B 6B 79 10 BC FF 93 1F 08 30 55 DB BC 1F
 0D 2A D5 03 B6 DD AD 70 09 D2 01 7E D7 2C 96 39
 AA 1C 19 1B CD A2 B9 AD 5A B2 15 C5 FF F9 47 2C
 08 0C 20 3C 9F F0 19 DE 7C F6 49 C6 8F 1C DA C5
 3B 98 40 3A C0 FB 73 DD 15 13 9D 28 21 A7 7B 7C
 3D EE 5E 7B A5 32 8D D8 88 61 AC FE CC 67 7E F9
 3D 1D 82 22 A6 77 D9 AA 42 ED CB E9 D8 24 A6 3D
 49 0A 06 8A 96 EC FB 9E 55 C8 15 94 E4 D1 13 83
 82 97 F0 F0 69 93 EB FA 05 C5 B4 93 33 D3 6F 28
 F5 06 14 00 78 15 37 7F 3F B5 2A 94 A2 47 79 90
 22 0F A3 D3 07 59 DA 3A 47 7A 9F 38 A1 FE 42 5B
 BA 31 B8 4C 5C A2 3E AC 3C 8F CE AB 17 54 FE B7
 F2 6D 8F 06 7A D2 25 D2 24 33 E7 A9 FC BA 0F 8F
 82 DF 17 22 7B D3 2B 2B BE C0 FA C9 C3 BB 24 EC
 BD 0B 47 56 B7 01 F6 8D 72 CB 1C 06 6E 47 C6 47
 F1 9E 21 43 99 61 D0 ED 5E DD E1 B2 82 3B 72 46
 0E B0 E9 86 5E 96 A2 3D B2 5C B7 E8 4D 17 FA 00
 61 6F 7C 94 73 02 6C D1 FC 98 F5 51 5C 31 B0 52
 DE 04 7B D9 D4 03 83 41 30 DF EF 8E 67 0F FA EA
 98 03 C7 C7 0D 17 B6 A4 FB F5 28 5F 2C 5C 32 F9
 23 D5 8B 9C 13 DC 95 56 39 61 A9 D5 B6 1E 81 37
 A5 07 93 B4 D2 87 72 45 18 F8 EB DB 35 F9 81 97
 7C 49 80 37 D0 9C B2 0E A6 5E 16 69 79 CA 8C B2
 FC 7B A0 05 4A 87 9D DA D0 7D 68 96 C3 AB 6D CA
 28 DC 04 57 4C 97 03 84 70 66 F9 82 52 19 C9 C6
 5E DD 3B 8F FC FE 83 15 96 3E 5C 97 15 1D 36 04
 91 87 68 C9 9E 71 9E 4F A4 13 D3 4D C5 AE B2 B2
 06 4B 7C 73 95 6D 02 53 07 F5 7E 92 08 CE 20 9C
 FF CD CE 31 C3 50 13 F6 19 84 46 7B 66 ED 8B A2
 8B C0 6D EA B9 BB 47 07 0C 51 5B EB 7E 8B FA 7B
 93 B5 D0 44 28 F7 65 34 33 3B F9 10 D0 70 E7 BF
 F4 D7 F0 91 24 8B 61 73 57 83 53 D1 CC C2 6B 13
 28 F8 00 54 5C CD 63 91 9D EB 40 79 3F 6A 44 74
 21 EB 86 E9 88 C4 03 5F 8C 72 7E DB 54 35 78 9A
 9A F8 C8 18 30 58 35 75 14 F0 C8 E5 85 14 E9 EB
 5A 8C 58 5D 34 59 A9 94 A3 FE B4 09 D7 F6 6F 58
 BE 05 D7 A4 86 76 AE 68 36 97 6B 4E C4 C4 37 F1
 F0 3E 30 C0 BD 72 6B F1 74 43 03 0B 67 90 66 B1
 9C C5 2B C6 A8 C9 34 8C 4F 6A FB 48 64 FC AA E1
 DE B5 D4 44 74 E8 E2 82 20 16 29 CF 6C C0 5E AD
 CD A4 11 16 2D 9D 6A 7C EE 60 75 D0 A6 79 82 F0
 9A 5C AF 90 28 30 54 12 42 BE 95 AE C8 C1 08 E0
 DA 2D 12 DC C8 9B 7C 73 EF EF 99 7A 79 95 A8 0C
 22 CD BE FD EE 54 4C 2E E4 14 E6 63 65 12 7C 5D
 FD 36 62 0E 1C 6F 91 42 28 BD 38 68 3C 96 37 7A
 37 98 EE 7C FD 90 88 34 8E 0E 88 EB D7 0B FB A5
 CC 7D B3 5B CC 91 3F D3 CB 5E 61 0D 4C 5E EF 29
 63 CE 37 94 A4 75 91 56 14 9E 60 65 8D 32 86 56
 60 90 65 82 DB C9 2C AE B6 1A 7F 29 41 E9 F5 98
 49 30 2B 35 EE AA 1B 42 18 6A E6 1D 68 06 95 43
 CB CA 7C 58 13 CF D3 75 7E CD FF C8 4F 66 A3 A5
 B9 0E 31 6C 81 75 9A 44 6B 8D 2E 4B 51 3B AF A9
 6F 60 4C 8E 07 A3 87 69 01 BC 56 DD 98 7F CE BF
 CC 0C CC 14 5C 69 2E AF AE 0A 85 38 8D D9 DB AF
 77 7B BE 10 56 51 58 08 B6 3C 73 DE A9 AD 6D 2A
 20 2B 32 B4 50 34 56 33 18 3D 71 8B EA 19 6B 9F
 0D 27 DD 62 DD 34 0B 6F 94 3C 0D 02 DA CB D1 99
 89 C2 DC 02 BB 16 3A 05 83 DE EB 39 91 44 32 8D
 F5 E1 9E 22 2C D2 AB 6F 22 18 03 15 D4 76 EC E0
 03 09 E2 F2 51 01 C4 EA 4E AF E4 86 0D 8C 3E DD
 A7 30 EA 8D 0B E0 74 88 ED EA 04 D7 04 34 0C 03
 FC 54 8D C9 F9 82 B3 8C 46 C3 65 1C EB 63 35 D7
 B7 A1 BC 14 97 E6 02 9B 3C A1 F9 3F A3 87 FD D8
 56 EB E8 35 E6 7D 17 1C C2 A8 20 87 25 61 D6 04
 1C 83 2B 84 82 68 D0 A7 E3 B7 D4 F9 60 DF 3D 18
 6E 5E 06 E7 08 FF 0A C6 D8 01 82 15 5A 44 55 A0
 9F 9F BB D6 78 A4 FE 1E A6 EF 29 5C B2 50 0E 12
 04 D8 75 44 54 E1 ED 3B 2C E3 01 A6 24 95 77 E6
 BA 02 69 26 8B 69 F1 CE DA B3 BC 0A 83 D4 6A EB
 D3 B2 39 03 B3 E4 DF 00 05 8A D0 1D 92 84 43 18
 3B 47 7D B9 3A 4E 1B 73 33 3E 53 FB 5F E7 F8 B7
 02 03 75 48 B2 5D 2F 70 42 F9 65 36 8A 6C 40 61
 01 31 F5 5C B3 3D E3 0D FF 9B 78 5B B5 40 1E ED
 0F B4 C2 1D D3 D7 16 C7 37 CE 86 EF 65 A7 E1 23
 53 40 1A FD 9C E3 22 85 ED 9A 76 16 60 0F 85 4C
 9E 1F F5 BB 46 1A 07 2B 80 7C 1C CA FB 78 2C 90
 CB 1A F2 44 37 59 C2 A5 7D 98 B6 14 46 8D 99 48
 CD 7D 65 D5 34 FB 2F 69 05 60 1F B2 BB B9 3C 4F
 47 44 4A 72 4B B4 3B 00 71 A7 EC 4C 1A 57 EE 7A
 CC DB B7 12 69 F6 80 5F 51 A8 88 E5 6B 18 1D 92
 17 16 CA 96 84 92 95 DD B6 37 06 5D B1 2E D0 4A
 91 C9 94 0A 5E D9 70 43 59 04 D3 F8 B5 3A E4 29
 C0 01 08 AE 2D 74 51 05 BE 46 86 B8 D3 92 EF 27
 17 C6 13 B5 E3 80 F8 A8 3E 19 BD 33 38 1E 43 DC
 8A B8 8D 13 D3 08 02 8B 72 ED 39 A1 4B 53 2D 1D
 32 94 71 12 8A 80 A6 55 C3 84 75 FA F8 B8 CA EE
 AB C3 AE 02 A6 D9 21 22 D1 F9 BC 25 B9 DD 90 83
 A0 94 72 8A 7F 37 97 A3 12 6F 4A 30 8B CD C8 61
 D3 BB AA 6A D5 77 78 9A 65 AD 00 16 CF 73 E2 0D
 DB 2E 11 09 24 89 D3 BD 21 9A B7 03 FE EF 70 A6
 88 35 ED B1 CF 50 68 C7 CB 26 0E E6 BF C5 B2 C9
 4A 43 FD A9 49 5E 8A C0 4C 35 88 35 75 F0 67 1C
 1F 25 57 F6 BE 7E 3B 5C 60 C2 6A B6 9D D4 24 87
 23 69 75 6D D5 0F 77 92 27 DA C9 88 D8 33 62 6C
 15 E6 88 CB D1 BC 7F 04 99 DF AA DD D1 9F 74 D0
 F0 F3 76 13 2D 4F 69 15 30 B9 05 6B CB FA 3C 15
 DC 45 98 F1 3B A5 2E 99 16 5C 1F AF AE 62 31 48
 9A E3 D7 8B 67 F4 18 41 B1 EC 1B 0A 30 40 51 E7
 77 70 E2 F9 0B 84 40 35 E8 DD 5A F8 E4 6F 02 7F
 A4 5E E9 C9 B3 64 B3 15 36 62 A3 BC A1 99 C0 C0
 0C 24 98 DB 39 D7 D8 4C 6D 1F F0 8E 10 14 40 55
 62 35 44 14 A5 75 63 0A 70 3C 4B CC EF 2A DF 7C
 1A 45 A9 FA 4B 72 2B 86 0B 15 3A B9 CA 4C 21 FC
 63 DE 21 69 5E 79 AA 79 70 FB C2 7D 69 E8 C5 84
 AB EF 15 FD B6 F2 8C 77 B5 A6 22 C2 2C 70 D0 A0
 4F CE AE CD 9B 82 A5 54 A6 2A 1F 91 31 7B BD 7D
 37 BE 8C F3 F3 02 80 2B C1 31 9E D7 78 5A 3F C0
 0E D2 D2 81 8D 3A 4D F0 8D 8E 1C 71 CC F3 14 56
 5F 1C C4 0B 94 CC 92 25 3E 5D D5 2C 7F 1F 52 94
 62 24 66 9A 72 AF A1 49 1B 32 4F D7 FB 6D C7 D5
 ED 8D 77 2E 43 25 A7 69 76 5F 4B B1 29 2B A5 3E
 0F 78 FE 24 94 91 29 98 A3 29 19 AB FA B7 52 9C
 FC A8 42 4F 67 14 13 67 73 82 92 57 11 00 E8 99
 E4 ED 36 40 A8 40 34 B2 1D 49 37 4A CB EB 19 D7
 FB 14 87 AB 09 E3 57 DD 6D 0F A0 04 33 CB 49 67
 27 8B DA D6 8C 59 B9 85 93 2F 2E F9 88 8F 28 04
 C8 2C CE 1F A3 B0 85 65 3D 0A C9 A1 FB 72 48 0B
 42 D9 19 99 56 D3 61 21 0F 16 B0 CB A2 C0 D6 AA
 2C D8 96 71 B0 D8 09 EF 1B 5A 9C 4C 9E B3 9B 72
 59 94 2F AF DB 5F F7 5F EE 9A 22 2F 3C E1 FA F8
 29 2C 8A 60 D2 5D C0 92 46 A9 13 3D 8B 72 3D 71
 79 1E D1 C8 92 78 84 48 23 F3 57 33 D0 F4 38 03
 C5 33 E7 BD BC 3D 51 98 49 29 27 0C 8F AB 9F 12
 F5 45 B7 3B 82 0C D4 25 BC A4 0D 68 59 E8 B5 B4
 6C A3 45 4E A5 64 70 BA 51 B7 E8 4C F5 FA E3 CE
 85 37 9E A6 14 D6 8F 2C 84 83 F6 8C E6 B8 61 F8
 2F 61 08 12 34 E7 CB 16 D5 3D FA 9F DE 2A 81 E5
 1B 2B 20 79 C4 4B 50 31 8E AC 9D E1 5A 1D 0F E7
 01 74 C3 1B 0E 47 E4 DB 4A 42 62 5B 06 4F B6 AA
 60 7E FC 02 B2 F0 6D 9D AE 08 61 7E F7 50 1A 81
 5D 8F 54 B2 0A DD A3 82 E1 53 D2 64 27 38 89 82
 CC 4F 74 08 E7 31 31 70 21 FB FF 81 0E 07 7D C6
 61 3D FA B7 C3 58 BC BB 9F 74 B1 A7 80 22 57 BD
 37 AD 69 07 18 55 72 37 B1 A9 3B CF 4B EA 7A 76
 47 8B 1E E4 EC DE E6 62 DC CD C7 19 E2 F0 AC BE
 67 5A E2 50 29 00 70 E3 F6 34 32 74 36 B1 41 DB
 55 EB CF 21 8B E7 22 8A 2A B2 37 A5 3D 48 C3 9D
 36 18 00 02 24 8B CF C1 67 10 C3 29 3B E6 FC AA
 FF 91 6B 6A B0 7F F7 7D 6C A6 FB DC 9A 29 09 18
 94 E6 CE 60 0F EF 8E D3 06 BE 02 EC 89 F9 8C 24
 A2 60 04 A6 4F B4 01 6B 16 FB 20 78 50 6B 19 CF
 35 C5 D2 01 17 FC 8B B3 11 FD F6 B5 35 24 D4 05
 29 8C 5F 4F E9 A9 2E 17 4B D8 4D B2 CE AA A7 28
 87 21 0C 56 2B 56 AC 7A 37 61 B6 61 D5 9C EC B5
 A6 54 F8 8C BD E3 B6 F7 75 0D BA 36 58 A5 B6 14
 6B EF DF 67 C7 21 59 8D B8 F5 47 0E D4 56 B7 A7
 49 07 6F EA 2F 20 50 90 0D 36 9E 08 3F 67 BF 55
 7D BD 3C 7D 86 7B E8 8B 01 26 E9 3F 78 3A 58 2B
 A7 2B B8 C3 36 02 0D 8D 42 A2 75 F6 8A DE C1 A9
 88 C2 70 0D 1D 06 E3 C8 90 2C 1B 03 53 C7 C5 74
 0B 43 4C DE E1 38 27 B6 E0 47 20 10 8E 4C F4 E3
 51 91 69 5D B2 4F 49 6A 28 0B FD 4D BA 04 5E FA
 DE 58 7F 98 46 59 EF A4 57 9F 04 BA 9D 3C 13 AE
 E1 40 38 A8 1E 4D BD A0 44 3B FA EF 91 79 86 6A
 36 24 FC DA 06 12 F2 6B 80 1C 73 BA 98 03 22 65
 75 40 89 E9 83 3E D9 8C 83 30 72 D2 37 06 08 05
 A0 3F E1 5E E9 53 10 43 EB 2B A1 74 91 7C 6F 56
 BD 94 4A 0A D2 56 E0 1D 19 CE AD D8 92 34 49 F1
 E1 3E 92 6E BE 28 DF 8E 69 A8 00 C9 94 10 7B AE
 8C BA CA CC 33 6F 73 37 05 44 88 A1 D3 49 CA BF
 4E B3 77 D4 F9 FD 2C 46 5F 25 D2 38 4D 2A 38 71
 E5 09 39 F8 28 10 6A 0E 4D E3 5D 1F 1A 52 F8 9F
 C7 A9 38 65 DC F3 1A AC 3A 93 6F BE D5 56 63 22
 11 D5 69 E0 94 8E AA A2 D2 E5 FF 0F 2E DF BF 7D
 8B 3A B0 10 77 93 30 3D A2 E0 BC BB ED 0B 40 40
 2C EA 3F 3B 09 C9 CB 39 DB EF DF 4E C2 E6 5F 61
 12 A4 FF F7 F6 CB EF 78 1B 6C 4A 09 06 BC E3 D4
 58 6D 52 47 A8 9B 3B 16 ED E4 B7 16 EF 66 27 19
 92 CD 1B B4 2C 9C B2 47 F7 A3 B7 F3 63 AA A5 AD
 1B 70 FF 4C 5C 5F 24 16 36 1B D8 B4 B9 0E EE B2
 F0 60 00 BB 3D C8 21 FE F2 B4 CE 42 72 60 07 FD
 9E 6B 38 44 40 41 64 4C 38 A9 DE 91 E8 A4 EE F7
 69 F0 2E 55 91 7B 50 9A BA 4E 49 D0 97 85 6E 7C
 7D 11 2E 42 45 F2 2E 63 F7 DC FE E5 EC 58 71 28
 37 E0 F8 03 02 08 5D 77 0F 60 F2 E9 85 8E 9B 1F
 97 1A DD 50 1D 0C 1A 9C 8F BD 34 8A 59 EB 4F 3C
 D0 57 FA 46 CC 6E 2C 16 98 A1 DB 05 F2 AF F2 B7
 2A 0F D1 E0 36 49 AD DE C4 C7 20 98 6F C8 31 7D
 AD 7F 51 29 33 6C 4E E7 6B AE 18 7E 9E F5 34 D4
 30 A8 2D 81 6C 0F 93 33 E9 26 7C E8 9A BA 11 88
 CB 26 14 42 C2 02 BF 1F 59 98 3A 19 DB 40 9E 86
 A2 A5 00 9F 52 82 F0 18 0B 91 B9 0B FF 7D 78 80
 7A 90 D8 7E 13 49 FE 73 CC 21 6D 8E BA 69 AB EF
 89 AB 61 31 6B B9 BC 66 87 E5 7B A3 36 E1 8A CF
 D6 5E D3 A1 9E 05 AA 57 98 A1 01 4D D4 8B 92 4A
 2B 04 DE E4 03 F2 3A C9 C3 BA 5B B5 B3 A2 DB E8
 84 92 7F 74 06 C4 70 20 82 EF E6 A5 99 66 AC 84
 30 90 ED E9 4E 85 7F 55 12 A8 24 90 A0 ED 1C 34
 84 82 6F 46 1E 37 07 43 78 AA 55 A7 7F C6 B4 BC
 06 C7 C7 A7 C8 52 EA F0 68 A8 AC 4A 53 B4 3C 52
 74 E8 E8 6F 28 92 96 AB D3 8B E4 35 26 6F 93 35
 C7 16 FF B8 BD FA 0C 2D 5D 6A F7 D1 2D 4F 5E E6
 FD FC 05 43 C2 62 A5 27 3E 8F 74 16 44 0B 82 D2
 D2 5E 32 FB 7F 62 36 6E 19 60 0C 39 57 EC DD 2B
 AC F5 3F 96 31 6E 62 82 B3 6B B1 EB F7 C6 1D A1
 9F 8E 5B EB 27 DE BF F6 1D 58 A5 9B 76 01 0D 6B
 70 91 52 6A 96 36 1D E1 9C A6 C9 97 E5 04 44 5B
 DB 0F A6 F5 D6 FA 57 9C C5 FD 6B BE 73 CA AF 5D
 2E F2 38 46 92 2E 54 85 DE 18 E9 E5 BA 0C 49 7E
 D0 B0 DF 50 F7 CE AD 50 E7 96 D0 A5 6E CD AE 15
 FC 81 2F 99 AE 64 63 C5 0B E1 C3 A5 96 10 09 EA
 96 D7 4C CE 9E 0D B2 07 18 79 11 CC 9B A5 E1 62
 C2 89 9B 4E 30 84 14 A9 47 39 1C FF B4 F4 BE 29
 25 16 A7 06 49 22 B6 FA D9 CE 20 47 A5 7F 1B E5
 C1 B1 3A A6 15 40 B9 B0 5B 65 80 8A C4 2E BE 80
 B2 66 F7 B4 72 97 56 26 8E 39 37 BA 2C 4F 55 03
 E4 77 D6 7B AB 7E D5 63 0A B6 A4 55 E3 DF 81 CC
 E1 A0 17 F7 A1 49 0A 31 F3 DB 5F B3 A7 E3 A4 86
 28 4D A2 AF 0D 84 FF 44 67 30 13 C1 43 81 C2 C6
 12 D6 70 7D AC 7E 82 26 FC 20 36 36 57 F7 8D 61
 6B 2F C2 6B 92 4F 2A 2F F4 48 61 14 31 A8 5F AC
 98 33 C0 79 6D 24 51 DF B6 4F 3A 82 AC F5 CC 0A
 1B 89 CA 49 1F FC D6 22 93 D9 DF 07 33 38 F4 43
 76 15 5F 5B 3F 77 38 9E F0 A9 9D 85 E2 D0 40 12
 8C D5 74 DC 3E C8 4A FB 5A 94 66 7C D6 F8 0C 1A
 76 AB F4 DD 67 D1 28 85 6F 7B 99 82 3E F4 06 08
 59 59 FE 08 AA 89 43 C8 CE 47 E2 8E 0E 2D 9D 49
 73 82 A5 DA DD 8E 9B 75 BF DA 2E 8E C0 CE 2F F4
 F7 F6 D2 3A B5 73 90 31 2A 8F B5 42 56 19 69 76
 54 90 C3 03 91 DA C1 09 52 36 C7 B1 48 74 A1 6C
 59 2A 2A DE BD E8 43 E0 52 B2 D7 57 22 60 9F 32
 AB E8 DA C2 8A C4 D3 B5 D2 8D 1E 6D 04 8D 34 9F
 0F A6 CF B2 B1 51 1F A0 CF B6 22 54 58 51 CE D4
 31 61 EB 3E 09 B7 10 0E 79 DF DD 8A C6 1E FD A0
 E8 6A 9C 7F 5F 30 B8 25 57 92 98 22 19 5B 93 04
 79 24 5D CD D5 97 D7 B3 71 F3 52 CD F1 EA C5 AA
 50 E0 F8 69 FC 87 75 5F 57 0A 18 A8 20 38 F3 82
 30 9D 77 26 34 F2 C5 0C C7 0C 41 7E AB 05 C0 98
 49 83 71 E7 4D 22 08 E5 D2 F2 D8 5C 1A 18 FA 5D
 0C AF 1B 1C 72 85 BE A8 31 2D E6 27 5F 82 64 B5
 8C BA 94 57 A7 BA 3A 9F C4 8F 92 3B 18 81 32 1F
 E2 B3 23 03 5B 1E A0 CC 84 7A 57 C7 FE 7A 6A 0B
 D1 1E 99 5C 66 13 AE 82 94 CB E9 73 C1 79 F8 DC
 E1 92 E6 11 C5 12 5B 85 91 CC 5A 44 3C A2 B3 B0
 97 E8 E4 7B E4 9C 2B 97 6A DC D2 AE E7 85 F9 2C
 0D B0 D6 EC 99 3A CE D2 81 0C F0 59 5F 8A 4D 95
 11 D3 F8 9B 05 CC 3A 72 F9 F6 41 6B 8F AC 2F 95
 CD F7 8E DD DC 60 61 85 76 85 CF 87 EB D1 AE 17
 DF 1E B4 3B BE 00 19 0A 4B 70 53 69 67 0B 9F 60
 CE D9 1A 65 6A 6B 7A D8 BF 61 16 F6 A8 CD 32 F2
 B9 7A 55 3F AD 23 B0 23 E3 7F 50 10 41 A6 63 28
 86 F9 68 51 CA 5F 46 03 7F D8 11 92 73 B2 15 EF
 70 46 83 66 88 0B A7 97 20 6A 54 F4 C6 DB C7 9D
 B3 D8 B9 E0 46 48 86 90 23 CB 57 A6 ED 66 87 50
 A6 50 A9 12 53 7A 6B 80 48 62 7A 0B 74 82 63 16
 A6 DE 9C BB C9 2C 2E 9D 4E 4E D7 EA 94 2A A6 EE
 6C 09 75 EE 20 EB 27 AB 5C 4C 51 96 83 F0 51 56
 BC 84 36 59 D7 FD 28 3E F6 81 A8 4C 28 C0 9B F9
 E0 C7 FF 4D CE D3 6B CE C3 1E 4C 8D F6 E1 CA 85
 9D C5 EA DA C3 91 B1 5E D9 56 59 EB 0C 8F B6 84
 E7 FE 60 D0 D6 97 50 E3 9B 21 91 BA 95 12 01 A9
 5C 21 1A 26 0B 85 6E EA C9 9B 2B 44 49 15 82 AA
 3A 33 B9 A8 DE 8F 0A 6A 4A 51 9E 2C A6 57 FD DC
 4B E5 5D 76 5B A6 8D C0 DB 7D 99 BA FC 9B 07 E8
 22 A5 D5 7C 6B E7 BC 1C C5 7A BC 9F BD A3 62 66
 06 A6 34 3F 44 38 AB 65 D3 5F 17 BD AB 4D 43 03
 65 76 D5 77 27 E8 C7 7C 74 0D DC EC 6F 0D F5 AC
 E6 E5 91 F7 7C 7C 76 B4 D7 53 B4 D0 0A F5 16 4D
 C5 4F EB 38 09 BD 2B D9 38 A1 83 04 92 7B 11 5B
 2F BF 26 21 C9 71 A5 C5 1D 01 3C C6 07 CD 2E 08
 D2 2F 31 64 11 87 DF 7A 26 DA 7F CB DE 2A 6C CE
 58 7F 42 B3 4E DD 71 E2 24 DC 80 F8 7A 8D D8 25
 43 8D BA 2B C4 5D 99 F9 58 38 01 0F 69 5E 8F D8
 D0 1B 1C 8A E5 C4 18 A0 2E 41 A7 7B CA 74 E0 97
 A9 B9 17 BB 30 C2 E5 EE D2 1A 60 99 60 E1 A2 96
 14 D5 49 64 B2 0C E2 0B D7 86 9C 86 D6 9B 12 67
 FF C0 FE 12 9A 67 22 75 D4 6F 79 C3 DF 66 41 6B
 39 D0 F9 37 1E F6 8A EB 08 92 E4 E7 9B FC E5 8A
 F7 2E 11 75 1D 3B 30 A1 5B 65 92 15 2D 0A 1E 4A
 C6 8A 1E 57 B8 3F FE A0 65 89 33 59 36 2F 5D BE
 18 82 6D DF 01 59 03 4C 6D 98 60 3C A8 D4 5F B2
 FA 4A CA C2 FD D5 91 0B B7 8B 67 03 D9 52 B6 40
 25 98 30 2E 9B 7A 2C 48 1F 2D 46 5C A9 31 91 44
 14 6A D3 69 03 23 81 02 A8 CA CF 06 6B C3 D1 BC
 ED D7 12 6B 97 66 37 DD 48 33 7F 87 49 C4 24 51
 7E AB 77 09 A0 4C C6 F0 40 C4 8F 48 6C EC 9C 93
 B1 C5 EB 02 B4 20 35 DD 23 D1 44 64 AD A2 26 A8
 B3 E2 5D 1B 78 7D 29 64 E4 AE 56 E2 7C A2 F0 1E
 AB B3 FB BA 6C 19 A8 7E BA 8E 0F 6D F6 AF F4 D6
 25 98 6F F7 00 30 E8 5C B2 89 21 52 42 D7 66 8C
 A2 43 46 41 FC 75 A6 46 E4 BB 6E 8A C6 DC 67 2E
 90 86 28 E2 DD 0A D5 D1 5E E1 42 0D FF 70 5B 90
 CD C9 E0 59 67 4A E2 E7 3B 2B A1 6E 6E 38 67 EF
 8F 97 91 4F 1A 30 5B B2 74 F6 62 6E 84 35 AD 36
 03 C3 4C A2 BD 65 EB 75 33 8C A0 23 17 AE F3 8C
 68 81 D2 D0 84 FB C9 E6 43 48 61 9D DD 2D 47 E7
 79 BA B8 D0 31 F8 C9 C2 FB A7 BB F2 AD D5 15 97
 13 F4 D8 0A C0 36 FB 1F 92 41 58 22 90 DF 0D D7
 BA 7F 12 38 49 11 A7 62 0B 84 F5 68 29 BC A2 2D
 BD 60 2A 2A 7F 76 63 B9 01 F0 69 35 89 3F 2E 0A
 CB 76 03 B5 B0 F1 65 6B EA 30 B6 55 DA 02 1B 4B
 B0 B6 09 AB 1A A0 8B 00 9B B7 B4 CB 6F F1 8E 70
 35 24 5C FC C9 BC 0A 12 FA AB 9E 9C 63 17 CD 29
 96 1F 41 2B 62 0F 9A 29 8E 4E 84 C1 CB 4F 40 3B
 6A 48 73 5E E0 63 3F 0A FA 62 67 BA FB ED 42 C3
 37 F9 C9 4C 3E 27 95 B4 B7 F3 B5 F4 04 FC 3D B1
 33 63 77 BC AD 2F FF 66 A2 19 21 E5 BF 4F 87 D8
 35 A3 1B C2 B2 84 B1 6A E5 9C B5 21 B5 F7 B8 E4
 99 8F 17 94 30 0E 30 CB DE D5 99 26 38 13 D5 62
 44 76 3D 08 A5 2C 5C E7 5C 0D 95 A2 28 C2 FD 9C
 05 44 BF 76 E8 5B BD AF DD C0 1F DA 84 D9 87 76
 8B 3A 05 85 DB 54 A7 DE 16 A2 A0 90 07 05 BA 5D
 8F 6F 59 03 27 7C 4C C9 12 42 D3 B4 0C 14 47 FF
 BD 33 AE DB 4A 65 4C 54 42 A4 BA 10 9F 1F 2F 5A
 ED 5B 1E 18 2C B9 9C 05 F7 0B 38 21 F6 85 9E DD
 59 55 E3 7A 65 C4 ED C8 C5 4D 15 F9 99 46 0B FC
 98 BA E5 74 A9 CB A9 98 C6 72 04 46 29 0B 77 E3
 0A 3F 53 B6 13 96 F2 84 7B A3 EA EE E9 B8 47 45
 88 1F 8E 22 DE 67 6B 75 55 CC 3B 04 C9 42 70 A1
 2C C8 8C 30 E9 A5 4B C0 31 37 2D B2 B3 E9 45 00
 40 48 10 B7 54 B2 D4 FD 4C 0B C1 19 D1 9A 45 21
 36 2E A4 8C DB 28 30 1D B2 49 6A 98 3E 31 0D A3
 C5 32 E8 48 3D B2 C5 D2 95 B4 5F 06 39 EE BD FB
 0B A8 C1 76 AD A0 5B C0 14 C0 8E 45 41 CE DB 2A
 2B D4 B9 25 C6 EC 0C A7 11 4C 74 50 66 A4 A3 C6
 C0 81 C0 F5 4A ED D5 74 E9 5E 23 AC CE F4 02 77
 21 5D FE B4 34 8C BA 25 0E EC AF 1C 7C 1A FE 0E
 E9 29 2B 2D E0 3E B5 89 1A 7C E4 78 23 A3 77 86
 B7 B4 B0 A7 6F 26 00 56 60 2D 99 9B 63 4E 8F 8F
 6F E0 3A 34 BB 68 71 FD ED DF 75 E3 6C 8E 41 6C
 51 72 CD 84 F2 3C D9 1F 6D 38 A5 E3 98 13 7E 12
 F7 09 94 BF BA E8 03 04 9E F8 1E 9C 0B BF 49 8A
 F0 A4 8B B8 C6 90 DD E0 38 DE 77 1F 4E AF 9A 8C
 8F C9 47 4F B4 67 FD CB BB 16 83 39 0A 56 54 F5
 25 63 FE 5C A2 AD 84 55 67 E1 AD E1 2C DE 23 AF
 41 0D 0E 4A EC 8C 66 38 33 B8 98 00 B0 66 8E 6F
 AF D3 5B E3 06 B2 5A A8 6E EB 90 11 4A 4C C6 01
 0D 63 22 70 3F F1 68 95 BF 3D 67 B5 C2 8F 7F B3
 A1 8C 0E F6 C9 BA ED 7E 44 1A CA 42 A5 01 71 4A
 8D FE 7C EB D6 C9 0B 1F 47 B6 E7 E2 7E 9B 64 03
 8E 2D 74 79 83 E4 68 48 84 0F C8 6B E1 71 F9 D5
 DF 08 2B 74 40 3E 6D 59 EF 62 8A C4 A5 11 A1 8C
 46 EE 99 6C EC CD B9 AF BA 91 5E E3 4D 9C 82 3D
 19 DF 9E 72 4B 55 FF 50 09 41 11 1C 52 6A 33 6A
 B6 15 A7 41 16 7D 14 40 F7 18 04 17 7C 55 E5 1C
 09 A7 51 9E 6B 94 3D 04 4E D1 0A 0F AF 2D A3 34
 E1 7A 7F BB A5 DA 2F 99 C4 48 F5 EF 9C 4C DB 25
 6A 4E 08 D8 05 B4 BB A6 53 60 0A 72 B5 0A 84 C1
 8D 3A 94 36 EC 5C 03 2A DB 0B E6 F5 5E 36 97 27
 46 BA 61 5F CA D2 D0 05 66 3E 9D 85 47 4C 8F E3
 A6 9B 0F 30 D4 0B AB 3B 87 60 F2 7D 92 F7 E7 E5
 50 D8 DC 51 AF 6A F4 CC A7 CF 5F 62 F7 38 C5 D5
 CE 87 69 EB 16 D3 CE 60 38 B3 60 24 8B C3 D7 55
 DC 35 FC 72 3A FB C7 3C 65 22 33 C9 1A 2E A3 47
 AA 23 46 52 81 E8 02 5B D9 BC C0 C2 6D 4D 06 CC
 43 DB F7 09 8E 45 53 0C 64 7C 8F 2C 9D 7C 80 B8
 12 8C E6 39 75 87 4C EF E1 67 D8 C1 06 02 C5 1F
 16 05 36 91 E1 70 FF 7C BA 71 B1 70 B0 2A 22 13
 34 E0 4E C9 3F CA F9 08 AC 49 B5 53 FC CF 86 5A
 6A 32 C5 FE 4A 7F F5 E2 81 6E 60 89 88 05 C0 C3
 1C 58 C5 06 21 CF 0D 39 4F CC D7 D2 89 F8 42 55
 8F 23 97 30 5B 23 1E 74 C9 28 2D EB A5 2C 11 42
 05 DE F3 5D C9 A4 84 71 76 30 D5 42 D8 45 65 C6
 82 BE EE 86 20 3A 94 8D D7 EC E0 BD 93 3D F4 18
 B7 B5 A1 30 9E 29 4C 66 3B 3F B9 38 E0 40 84 CE
 6E AD 19 A2 C1 B4 3B 21 93 93 84 A5 C7 FB 1C A1
 DC 46 75 DD 86 19 10 32 EE 73 69 58 3F 07 0A 63
 49 89 75 8B B2 56 FF 7E 5A 94 8F 99 55 0B 1E 59
 EE 5F 41 25 35 5E 1C 99 FD 61 5E 3F A0 C9 3D 17
 49 6F DF 5F 8C 7B 55 26 0D 7E 52 46 E4 07 C5 69
 66 A3 B3 C8 EB 91 87 84 AC D2 32 23 9C EB CD 1E
 2A 0D 1D B1 E3 84 67 36 93 74 61 B6 5E 34 09 A2
 76 E2 9D 18 CD AA EA 1A 36 63 44 D0 F9 AB 72 95
 12 B1 EB 36 09 22 7D 28 F3 A1 68 EC AE 65 8E FB
 87 80 89 94 58 A7 06 18 51 03 38 35 71 52 04 64
 D5 6C 77 F9 70 10 53 C3 B8 3D D9 C9 C2 76 FC F7
 AD 4E 7B B0 2A 4A 40 C6 83 0D 75 4D FC 5A 60 1D
 85 27 EB 57 28 F1 68 0C 5D 26 F0 7C 8F 98 95 25
 96 ED 1E E8 D6 7B 1D 5F 70 32 7D AF 6C 34 2A 01
 2F 20 75 3D 89 F0 A5 C6 32 65 63 96 DF 82 84 E6
 ED 34 AF 9E D6 82 2D D7 9C E0 C7 A2 33 66 3A B8
 F2 DD 76 A4 9F 50 07 61 3A E7 BB E7 A1 12 DB EC
 A9 BE 12 97 CA 24 4E 80 AD 23 DC 78 CF 8E CC 3E
 3C 0B E6 30 21 5F 42 BA E0 37 78 C9 9E 0D BD CE
 3F 9E 73 3F 8C E6 BE FC 02 9F E2 10 DB F1 91 EE
 3A 9C C6 51 74 C6 71 CF 28 2D 0F 06 12 07 5D CA
 31 A8 2C F7 95 1D FC 9C BA 63 F3 82 FC DF BC C5
 3E 96 F3 EE 3F 85 36 FE E3 FC 4C F2 79 F4 A2 57
 3F 00 A0 B2 E9 3A 39 67 B2 22 B8 FD D3 8A F8 00
 D6 39 3A C7 76 25 D1 3C 0B 6A 21 65 2B 83 44 8C
 54 2A FE 8A 68 1A F9 1D 41 22 17 3E B2 46 FC C0
 2A 86 35 1E DC A7 7F DC 10 73 57 5C 11 53 68 43
 79 05 20 ED AE F0 A4 25 44 CC 32 DF F1 99 2B 1F
 F0 9B C1 EB 71 3B A6 D1 C4 BE 0C 17 A8 C0 EA 95
 C1 D7 A5 70 47 0A 1E C8 2D 64 D4 0E 54 09 1B F0
 73 1A 9F C8 DF 62 74 A8 15 B7 25 95 92 51 67 1C
 25 5A 16 7C 24 5D 02 68 28 86 00 5C CE E1 32 34
 ED F2 21 D9 D7 06 77 88 C0 CD 3B 4F 40 AF 93 CA
 21 66 BF 2D CA 87 91 4B B6 DA AA 09 4D A1 A9 36
 43 15 B7 78 B0 D0 E2 1F C1 7C FC DA A0 AD CE F6
 17 58 77 85 79 56 F1 5F D5 8E 2A 66 F2 68 A9 C8
 86 6F A7 0D FB D8 60 7B BD 26 11 5E 4F 39 7F 4A
 B2 F8 54 EB E9 4E CA F3 9E 43 86 23 93 5D B2 3C
 80 3E 60 05 E0 4E 72 6D 03 77 0A B2 B8 18 6E 7E
 29 B9 4E A4 F7 66 1C 4E 50 7F 4D CC 5E FD A8 FC
 69 AA 68 17 55 C6 8B 31 C4 5D B6 EC 4D 37 7D C8
 3E D6 3A A5 BE CC DD 11 18 43 AC E4 AD C4 8B 91
 43 61 8B 3A BA E3 FD 71 B3 8A A9 C7 E5 0F 3C 64
 88 C3 51 6A AF 63 A1 38 71 A4 F2 B2 52 DE 04 6F
 AC 45 4B 91 55 23 AB 73 57 09 13 94 75 69 98 44
 E0 DD F8 36 83 48 3C 5B 23 8E 79 D6 2E 88 D0 4A
 BE 68 44 2B F5 E8 AC 52 F0 B2 D8 39 88 6E 6F BC
 B7 B7 97 8D 98 1A 75 7A DC 86 F5 12 99 5D 2E 27
 7B DF 08 49 07 EE 00 E3 38 E8 80 A9 14 41 94 8F
 11 C2 23 51 6F 77 34 3E B7 F0 7B 23 47 ED 0E 3E
 9C 6C 9F A3 CF 06 7A EF 2B 79 98 BB DE 8E 8A 99
 ED 73 86 49 6F 0B 37 20 0B 24 A8 64 51 22 C5 E4
 44 0D C4 F3 82 BD 8A A2 6C 5B B9 B7 6C 44 1A 34
 CB F6 0E 0F B6 80 65 EC AE 73 ED 9F 50 C8 9E 57
 3C 0E D2 7E 56 8E E4 13 9C 15 32 38 03 9E 5C 95
 5F 5D 2B 74 19 5F ED FF AB AE 41 B8 52 A6 69 32
 11 A6 B7 0A A6 70 67 CD 7F EF 26 F5 62 C6 C2 94
 82 19 C0 35 2E A5 CA 26 AE 67 03 E1 CA C8 51 EF
 5C A9 2D 92 63 00 CF 1F A8 23 7C 13 F3 31 46 8E
 21 17 03 13 80 ED 91 25 CB 87 FA AD 6F D6 EA 96
 BF 8F 71 03 86 A8 6A 20 CC 56 B4 67 BE 17 20 46
 00 67 3F A9 23 AF 2F BD 79 6B 13 63 77 38 38 7B
 0D 9A D0 46 C1 4F 33 54 41 33 EF 06 D5 06 3E AC
 04 CA 02 B1 0B 95 0C 28 26 3F 6A E1 A1 76 AA 30
 D5 BA B8 A5 E9 11 B9 3A 83 68 45 15 4E 14 25 54
 BA B8 D0 41 C7 D5 D8 06 29 0C A9 22 D8 2B 8B C2
 3B 8E FD 30 5E B1 5D 10 30 0D DF FD B2 5C 80 A4
 5A 08 C3 1E 45 40 02 6A AA 10 F2 E5 31 9E 3C 7D
 0B F0 F6 3F C4 90 40 92 66 BE 52 52 3C 6F 02 20
 1C C7 B1 54 2A 84 A9 7D D1 08 77 63 D5 56 6E 23
 ED F6 72 14 84 CD 9B B9 EB 70 58 61 F5 48 C0 72
 68 9C AF FC 74 A9 6A C9 39 DD 9A 0A 02 81 3B 4E
 36 AE 47 79 3B 95 22 65 E6 2F 19 27 FA 21 3C FD
 C7 8F 91 48 1F E7 45 2D B5 79 7C 8F 35 44 61 86
 7B 2D E2 34 EB BC D8 A8 EB 10 34 D7 AC 9D AA 5C
 5E 13 CF A6 01 EC 6F 13 AC 93 49 79 53 F0 E7 A3
 AF EC 6C 98 DA 29 16 E0 37 59 70 DC 58 CB D1 FA
 28 A5 CB CD E1 24 35 9B AD 2A 75 57 2E 54 70 5F
 7C 2B E7 DA 45 80 15 7C 90 45 40 AF 77 B1 5C 3A
 F2 D8 6E 19 E6 4D 5A F6 78 A4 F7 44 A9 66 2D 71
 6D 13 F4 88 0B 3D 68 87 F1 9B 80 E0 F2 60 99 F3
 F4 7F 49 71 46 F2 53 3F C7 20 C3 7B 40 CD F1 C8
 52 1A 09 BD 3C 7F 46 EE 0A 54 EE E4 A5 54 AC 59
 3B C7 7C C3 E1 CB 31 C6 AF D4 E8 15 AF 76 E6 2D
 60 CD 86 17 CB BC 47 4A 38 1A 9C 97 CA CB 00 A5
 F0 D5 FF A5 16 84 95 AE 34 7A 49 EF F1 87 A1 A5
 41 F4 B2 77 BD 67 9D 7D 2D 28 82 87 5C 6C 22 1D
 93 A3 6D 24 18 BC 84 B1 B2 DC 31 CB 35 6B A5 C5
 AA 8B B5 A3 AB 61 09 15 CF B6 31 EE B0 B8 D8 73
 88 0F 86 AE 4D 54 49 3E EA 5F 8E 49 40 64 4F 74
 2B 70 BF EE 37 B1 50 EE BA 85 5E 0F 97 30 B2 86
 5A 5B 16 65 CB 75 0B DA 89 73 E5 1D 87 CB C0 1B
 0F 20 B9 7B 2C A5 34 F9 E4 9D 5B 25 D3 28 4B 34
 3A 19 21 19 1F E4 22 3D 48 3B 96 68 F9 3B EF E7
 0A 7A 14 17 E4 C4 1A FE 00 3D F5 76 D8 20 BC 4E
 4F 54 48 BB 7C D6 A9 D1 36 B1 52 67 F4 C0 9E A2
 2D 71 28 AC 34 85 87 EC B7 1E DF 41 79 D3 77 F2
 17 9F 23 EE B1 06 1E DD B0 14 CB 39 83 80 F3 57
 B5 FC 22 FB 30 2A 7C FC 3E 84 43 EC 3D 82 97 58
 26 1A 0E C5 53 50 01 2C 16 A7 09 75 0F D0 AF 2B
 BA C0 58 9D 35 70 79 A8 6A 70 01 54 DF 3F 07 D5
 54 DF A3 64 91 C3 29 56 D4 04 42 1D 29 95 E0 EA
 68 B3 8B AC 9A 59 08 3E 31 FC 98 79 9D DA A4 D2
 D1 82 29 C1 11 E6 AF 4F E2 41 6F FA FC FB 25 2E
 D0 2B A3 CD 47 2B 52 6E 8A E5 07 04 22 5E E3 E8
 EF D2 7A DF 81 91 35 62 1F D2 01 A7 78 A2 3C 43
 D8 55 B8 8D 5D DF FA 5B 5B E2 D2 0F 10 0C D3 27
 20 57 55 38 76 40 55 D9 82 1B 89 FA 5E 7E CC BE
 22 1B 8E BE C4 17 4F 07 CD 05 84 79 BF 3C 25 60
 03 B8 40 D1 B6 8E 3C 31 A9 1B 7D 49 45 A7 18 EA
 84 C5 0F 2E FF A4 7B 23 98 47 56 E6 A4 F4 6E 68
 FD 3B 95 3B 04 04 6C 30 DB 40 F7 BA 27 F6 EF 1E
 4F C4 F3 6B 0E 66 2A 19 5C B3 28 84 DA F4 BE 35
 BF 7C 10 38 54 BD 0E 02 53 34 A1 BD A7 87 2A 46
 26 56 09 AC EC F2 BF 45 21 51 A4 C7 0B 2B 0E 0B
 C3 BC 9B FE 30 A2 19 D6 D3 58 43 C8 15 32 AE 59
 38 9F C5 30 72 86 3A 97 2A AC 45 61 D0 B5 98 9D
 C2 E0 0F 8B AD 00 A9 FD 38 74 34 76 E1 83 65 9C
 AF 2C 60 86 4B 62 C0 B1 1F 81 9A 44 B2 41 BE 0F
 0B C2 2A 30 BA E5 68 8C D3 11 B4 A6 56 AB 22 7A
 FF 6C 2E 97 8C DB 0E 7A E2 35 AD 14 9D B8 8B F2
 91 F4 70 3F 0E 9A A1 0F E0 DD 3A 9E 21 AC B2 19
 A7 95 E3 AF DF C7 E6 19 C4 11 44 7E 32 17 A7 BF
 6F 84 C5 6A 0D F0 DC 33 3E C6 76 B1 9E 2C 6D 07
 A9 72 26 C8 5E 15 CA 62 E4 CA 1B F4 A8 E2 EB 0C
 B9 D9 10 18 64 8A 56 06 21 67 4C 69 B2 3C 41 B4
 E6 08 10 F7 EA 69 F0 19 EB FD 5B E3 33 D5 22 E5
 AE BD 9C 4D 9B 38 A8 F4 F7 F6 B6 6B 7D FE 93 5D
 CC 77 A0 1A 5C 87 4A 0F A5 1A FC 35 11 11 9C 79
 D7 95 FC B7 31 A5 60 95 87 95 A7 B0 21 6A 19 A2
 E6 04 EE F1 10 21 7E 74 7B 95 1E 45 44 D0 5C EC
 65 48 4C 5A 42 61 EC C2 44 4F 0E 98 B3 28 98 6D
 26 E3 8E A5 C2 FA 4F C6 20 C2 52 1B 80 9C 85 A8
 47 85 7C 83 AD D2 3C 06 77 00 31 3C 24 AC 59 E9
 14 9D 9B D3 B6 79 FE 47 A9 CB 64 19 4F 51 0A 16
 33 41 FB 35 34 48 CF 05 F8 55 A6 CF E4 57 D4 86
 90 51 B0 E8 E1 0D E7 08 F1 70 F9 D1 32 50 2B EA
 0C C3 C8 86 9F 02 BE FC 7D 88 0C AC FA 06 74 56
 BD 55 75 BE E0 D7 AD B3 58 EC DF F2 37 43 28 84
 F8 A3 43 70 AA 33 75 4D 01 2E 3A A1 CB F5 3B 00
 E5 24 E4 15 62 AB 5B 8E 27 9C 8C 4C 45 AD CF 84
 01 F5 91 A0 16 B4 70 D3 76 06 B5 C4 FF 9D 8B C7
 1F 44 EE BC 41 92 52 1A 33 25 C4 5D CB FD B9 0E
 3E 03 E9 A8 33 6C C9 83 90 83 72 34 BF CD CF 25
 1D DB 63 BE 97 6E B9 59 CA F6 13 5C A2 72 F9 15
 7D 0E 1A 4B 62 22 8F D8 64 B1 D0 9B D3 F0 A0 E3
 FA 69 E4 13 17 FE 50 89 74 77 6E BD E8 81 AC 94
 AE BF 71 F6 82 E2 52 D8 39 0A B8 31 35 93 79 4F
 B2 20 F1 CE 18 C2 B6 C5 15 3C 16 8C 61 75 72 62
 1B F5 9C 62 18 FB C4 4B 3E 0A 55 BF C7 81 D5 82
 A0 D1 91 90 1E 58 E4 9B 18 B9 18 FA 6F F1 9A F6
 B6 8E 03 79 AF F3 A6 18 78 40 D4 F7 45 1D 2E EB
 16 07 56 4C 89 32 8C 09 10 A1 0F EB 77 26 35 8B
 8A C7 FA AB 4A 5F 2D 44 DF 20 5E 17 85 E3 2B E0
 D0 A3 C0 BA CD 6C F2 3D 3A 32 D3 20 5E 1E 1A DF
 57 6A 05 92 B5 0F 7D 9A D2 00 8A 41 93 95 D2 0D
 A5 AB 94 5B DC 46 2D 9A 5F 75 10 D2 0E 64 30 83
 53 EE D5 59 9D 35 C7 C3 D2 D4 6F 57 4E 95 24 CB
 98 D0 50 8F 7E 1B 17 9C D9 48 B1 92 22 D2 3C A9
 DE C0 3A 3D D8 41 46 D7 0E 6C 29 7C DC 45 51 C8
 DF A9 E3 CE 3C E9 96 2F 5C FB 9E E4 DF DD 74 5B
 8A 2F 7A 56 3C 88 D9 A4 34 9E B4 73 DC A5 14 68
 31 F0 6E 23 8D 5A 6E 6E 4D 11 15 22 9E DD E9 9E
 18 E7 9C 4E 24 F7 2B 71 99 D0 5C B8 B7 34 5B 85
 69 2F 2D 12 B7 86 0A 67 F9 F5 8C F8 DC 3B 66 B7
 68 3B E0 16 11 6A 35 0B 87 CC 6B DD 3D 46 6B 17
 7B 27 6A 29 BB C8 E4 91 11 2B 42 D8 89 09 FC AD
 0D 7F 3D A9 2E FA 6B AE 0C 2B F4 C6 7E C3 53 FA
 21 50 3B 52 DA 4F 4A 9C AC EC 68 9A 55 2A C5 C4
 BB 26 44 E3 10 EF A8 2C F3 24 C0 39 97 63 79 C7
 79 7C 88 15 6A DE 03 80 B4 6A 58 28 A1 52 69 FD
 5B A0 C0 92 E5 40 47 96 AC 28 B3 7C 0C 99 C5 FD
 3F 1A 16 79 77 CD DE EB E9 4F FF D3 39 7A 38 80
 E1 9C 0C 45 05 90 A9 F6 E6 60 E7 A6 6A EE B4 F0
 4A 09 9F 3D 7C 7B 80 8F EC F7 B6 00 7A D2 3D 0F
 F6 C8 E0 68 D3 81 46 48 03 34 4B 4A ED A9 2A 8F
 3C 0F 9D B9 8F 3B 29 4A 4C AF F1 9F 84 99 44 E0
 CD 14 42 D1 03 72 FB 07 26 39 59 52 41 20 DD 30
 14 04 06 D4 0C 53 BA AE E5 91 8B FF 5F 75 94 B4
 E0 D0 C9 A7 4D 03 E2 13 0F AC A1 97 A0 88 20 55
 08 FA 7A 50 32 64 E0 19 6D DE 52 02 D4 A4 4A E6
 CA E6 04 8A 3A 8C C5 72 2B E7 D0 6A 9C 37 B1 DF
 B4 FE 17 E3 80 9C 32 6B 80 1B 3E 9E 72 F9 A7 63
 C9 E0 40 A3 19 40 76 60 80 37 EA EA 5D 5C 77 AB
 80 91 31 AB B5 96 9C 87 DE 20 FA A2 92 E2 DC 6C
 37 8F B1 BB 1D C1 8F 52 8A C3 D1 0F 89 D3 3A 73
 9C 1A D4 EB 7A 83 18 74 1D 68 A2 21 D6 CC 6E 38
 27 F9 DB 8E 59 6A 89 EF 81 B9 4C 22 8C 08 FE 96
 B1 1A FF 2A 1B BF 1F 8D 02 8B 65 13 16 22 29 F1
 F1 62 41 BF BB 40 0D 56 F7 27 BB 68 CC 15 33 0C
 67 C6 87 9B 4D 87 D5 CE 6E 6B 04 37 C9 62 6C 0B
 1C F6 3B 3D 91 DE 70 77 0D 0F DE 1C 71 8B 4B 09
 FB D7 B0 BC 21 DC 32 AF 31 7D 9B 52 AD 72 8C 9D
 03 FB EE 7D 1F D1 A2 0D 1E EA 90 2F D6 5A 6D 19
 C7 37 FB 34 DD D4 AA 4D F2 EE 79 C1 68 60 BC 4F
 29 FB 0B 89 8F F1 A2 BB 95 20 FE 34 CA 1C 97 B3
 9B 47 A1 34 84 12 48 E5 2D 97 77 DC 5C 4F 0A 90
 FF CB 40 7A C3 5D 10 27 2B 51 A4 94 46 E8 B8 A3
 4B E5 1B 76 F8 5B BF 40 1C 28 F8 8E A6 47 13 87
 D2 20 07 25 57 8E EA 21 CB 8F 7B CD 2D 92 F8 A4
 97 9D 63 FE 85 38 EF 4A 23 2A 20 95 52 09 FB 0C
 4D 14 E0 C2 65 14 CE 32 8C A9 F5 AC 2B 8C 04 AB
 CA 05 83 C8 00 CD 93 D6 52 CB A0 75 21 FB 97 B2
 C1 EF 4D 06 6B 1A 62 B5 08 7B 0B 33 75 00 99 73
 2F D3 1D 76 26 D7 A6 44 B8 D9 38 D2 62 B2 DB 19
 12 4D 5C CA 36 5B 64 D6 F3 B8 F5 82 FA C1 BE 76
 F6 30 3E D1 02 D1 0E 4C 87 BA 71 50 86 84 B8 1D
 74 8F 4F 2E 34 76 C1 C1 C4 BA 31 EC 3B F4 52 97
 D9 3C 8B 27 9F 92 F3 4B 18 5B A6 D4 AB E4 D4 E5
 9A 83 1B C9 DF C9 ED 18 E6 AD AA 48 E4 02 3A 80
 F1 3A 5D D1 E8 10 52 23 D8 1C EB 02 D1 AA 84 D6
 58 8D B0 47 27 E7 F1 57 21 70 A7 24 D5 18 DC A6
 06 E2 09 B7 C1 38 BB B2 78 A0 54 0A 54 64 A1 F0
 7B 20 70 7F 56 BC 73 40 B3 7D D4 A8 21 58 97 7B
 45 E5 80 0D 2B E1 2C 4E 12 59 5C 10 C8 0E 3F 34
 79 48 43 38 1D F4 31 0F 91 FB F0 40 5B 0E A9 69
 E2 9B 95 48 9F 18 E4 EF 6A 0B 1D 18 83 3B AE B0
 E1 7E F7 74 D0 6F AD F4 00 E4 E7 37 65 77 E5 11
 A0 7F 89 1B B9 A1 91 B4 67 E1 3C 76 81 D6 0A 1C
 51 61 CF EC 0A 6F 67 60 96 00 DE A2 83 2B 29 7F
 57 F7 56 F6 EB BA E9 03 D1 13 96 98 98 6C A7 87
 95 BB D5 A2 8F F3 B5 1E D3 4C 13 F4 76 49 B5 7C
 C8 3E 58 82 DC 4A C8 0B 5E EF D5 38 C1 AD CB 69
 F9 4E F5 26 CF D4 D7 66 F6 07 F3 3B 27 33 CF F8
 42 60 E2 BD 14 D9 F8 DA 46 66 A1 1A B5 34 43 A5
 64 E6 EB F0 BA 67 49 28 1E 98 24 44 12 62 01 77
 D5 CA 93 70 FB 05 58 FF 65 A0 8A 64 4B F7 12 94
 79 83 AA 9E F7 3F 46 13 4F 2C 8E 19 E1 9F 47 6C
 C7 7D 7B 26 89 0A 9D 9D 3E 04 B1 2C 54 F3 CB C7
 9F FE 69 C9 7E D2 18 32 7C 78 55 3D A3 65 D2 4C
 72 99 F5 39 DF 38 39 44 82 41 6C BD C5 EE 70 36
 10 7D 09 C3 B7 C4 2F FF 15 B4 47 C1 43 C8 B9 F8
 3E 35 04 B9 6B 99 B9 96 7E 3D F6 9E 3B 98 86 7F
 88 EC 78 69 E0 6D DB B6 32 E2 99 75 BC B5 51 83
 29 B7 55 D2 DB 3A E7 74 C7 03 27 2F 43 52 65 EB
 D6 0A 2A EB BD 22 FD C4 5C CB CB 2F AB 96 05 90
 60 EB 05 89 B8 9F C3 9E 9F FF 4E 06 CF 28 ED 9D
 A9 46 8D A9 14 19 86 9A 28 8A F5 2E 5F F1 B5 D7
 91 64 92 43 CF 7B AF 9A A4 EF FB 74 F6 14 6B 17
 03 58 CD 50 0F 5C 94 31 55 94 2B 3A 94 36 AD BE
 85 80 F8 C9 52 C3 28 26 42 13 15 11 E5 C0 2E 92
 8E A5 2C 11 22 53 42 51 9A 88 B7 7F 36 C2 FF 6C
 27 9F 18 A1 80 2D 1E E8 2E AF D1 26 86 4F 83 A4
 C4 09 8D 57 83 78 C3 CA F7 47 58 36 99 32 32 54
 0A 3B 2C 2C F6 E2 B2 7A A6 08 03 D4 DD 07 91 8B
 B0 29 3B FD 72 0D 55 7C 7A 26 F2 14 DB 51 D8 A0
 21 86 39 69 CF C5 AB AF DF 28 96 DF 74 AA 7D 89
 EA 4A 75 41 BA 4A 80 95 8C 98 76 64 83 D7 25 CE
 8C B5 55 2D AF 65 13 83 C3 72 F0 60 43 D6 48 C6
 92 A2 43 5D 7C 09 75 44 86 B7 C0 95 20 C1 E2 19
 14 0B CB 51 0E 71 DB 1B B0 4E 75 03 C2 C0 4C 99
 8A 71 86 CB 6F B9 D8 72 80 68 A3 98 7B E3 38 14
 6E BB A6 EE 84 A4 13 3D CD 8A 47 0F 6A 5D AC C8
 AB 76 84 26 7C 1E B3 74 3B 66 FC 15 7E 00 67 6D
 71 28 E1 75 5F FB EE 8C A2 DA 42 78 AB A1 A2 19
 1D FE 15 77 6C 57 7C BF 99 9F E8 00 63 ED 99 BB
 CB 83 40 08 4B AC 83 D7 59 5F 2F EB 97 81 34 25
 EF D6 9C A8 95 B9 1A 3F 96 F8 66 F5 94 D5 F7 40
 FA D3 E8 87 A2 91 DC F2 C3 10 B1 1B 2E 35 0E 63
 C0 C3 38 C6 3C F7 06 E5 E7 C6 05 F8 29 70 6D AC
 BE 6B 95 C8 25 C6 1E 33 3C 20 52 C2 27 38 C6 B6
 A8 D5 CC C7 57 7A B7 91 49 89 16 21 D0 08 BF 48
 D2 46 B8 69 98 29 90 50 8B BF 87 51 7C 02 6C 07
 3C A9 0A 02 D8 EA 69 74 29 A2 1E 3D CD 0D EC F1
 D6 F1 9A E2 03 27 34 12 07 E7 B3 62 01 1F 71 AF
 CC 98 E2 C7 38 4C 0A 5D 72 5E D5 75 13 0C E4 23
 37 D1 DF 5E A4 D9 F7 32 40 0B 03 45 5D 35 9F A0
 51 98 F0 6E 92 50 72 A6 5A FE F4 63 BA F4 2D 5C
 97 3D C5 6A 94 CF 30 DA 5E 52 E8 36 68 34 45 FC
 A0 DA 82 D1 B9 84 47 D0 4F 6F 3C 27 70 3C 31 03
 C7 3F 95 ED BC DB 91 D5 33 9E 6F 79 D3 48 8D 58
 53 30 91 3C 8B E8 CC 3B 67 B4 4C 6B 26 B7 C6 3F
 6C 40 77 04 77 66 4A D8 23 16 32 07 F9 66 D7 45
 4C 02 81 A3 29 4B ED E9 1E C2 BC 8B 8E 1A C8 75
 C2 74 C7 34 46 24 64 51 1E 4D 70 72 C5 C5 F5 16
 9A AD C8 63 BF 2F E0 CD E1 97 0A 9F 91 CE 3F F9
 CA 05 C7 35 72 DD 5B 97 5B 56 EC B8 83 48 B7 90
 13 0D FC E5 58 58 B9 72 82 E6 29 6A C3 96 55 54
 ED F4 1A DE 3A A8 21 DB 13 53 30 B6 5B 5E FA AE
 C8 AC 7C C7 00 FB 3E CE 9E D6 17 F7 03 09 D3 5D
 9F 47 5A 7F D2 4C F0 94 3D B9 41 45 D4 7C 78 0D
 81 48 B5 E5 EA 6E A7 24 83 A9 84 3B 1D C2 1A BC
 8F 20 76 45 39 D2 88 56 77 A5 A4 08 09 1C A1 70
 DC C1 F3 8A 53 42 09 70 37 5A 4A 1D 00 60 51 01
 C8 15 BB 61 6F A1 74 90 38 33 D7 11 15 D1 BA C3
 7C 2A 9C 35 10 F6 20 4A 81 B3 B0 8F 2A 3D AF 41
 B6 E6 2B F5 D1 44 0A 3F 95 3B 77 C9 7F 55 22 7E
 F3 68 BD A8 6A 9A FB B3 39 C3 6B B4 1B 02 98 99
 7D EE B5 EE 82 8C EA 89 AA 59 68 04 1F B8 16 EE
 4C A0 16 F3 11 2D 68 1A 69 37 95 1A AD B5 AC 18
 F1 3D E9 FF 41 E5 39 E5 7E 1D FC 2D D5 05 4F F8
 59 4D 05 D3 DB CF EB 36 D1 27 58 52 90 B5 B4 38
 F4 8D 37 44 C8 CE 2A 4E 5A 3C 9E CD E1 E4 BF 2E
 44 C8 F4 61 29 F4 FA 37 25 94 EA 4C 90 5B 42 47
 C8 1B 60 E8 6C BC 55 AA C9 E8 47 CE D7 5B 64 C5
 31 A4 40 52 B7 FF 69 5C A6 C1 F2 0C E1 51 DE 84
 2B 46 61 C9 17 12 78 60 1F 70 3B 54 8C AD A3 B7
 5D 1A A3 DD F5 74 30 30 B0 71 7D D0 04 4C E0 6B
 B8 32 75 75 E2 BD C3 BF 76 24 D3 23 C1 46 B5 83
 DC 28 2D 10 A1 3D A6 96 6B 0E EE 9A F7 F4 37 8F
 51 8D 3F ED B3 EF DF 04 57 1A B3 0C C2 96 19 A3
 E9 31 97 CB B1 CC 3A 6B DD 8B 2C 36 94 A0 D1 63
 D4 78 21 86 3C D4 08 AD 5D AC 16 60 FD 5E 22 CA
 5C 1B 54 88 C3 12 35 A7 00 4C 5E 37 6D 3E 87 4C
 55 3A 05 3B 33 E6 E6 1E 82 BA 9B 0D E7 EB 54 00
 41 88 93 DC 50 F9 AD 4B 3C 7E 30 6F 2C 14 D3 AD
 28 08 CE EC 9B 46 F2 F5 D8 5B 90 01 F8 79 CE D2
 5D E4 F8 18 1E 35 F4 16 6E 46 42 E2 13 CB B5 38
 95 2D 8F 54 01 D9 3F 7A 18 22 91 86 B5 3C 39 AF
 4D A3 18 58 77 CA 53 00 17 5F D7 71 0D 99 C6 8C
 78 6E 5A 5B F1 16 59 79 D5 3F AF 51 E9 21 7B 97
 51 A5 D9 02 96 F8 CF DB EA 3F 02 74 9D 86 AB B2
 29 FB 67 8D 30 3F 0C 9F 2A 8D 29 82 EF 45 67 F1
 B7 CE A8 B8 96 30 22 79 0C 18 13 F2 2D 03 C5 68
 0D 4B A4 0F 1E 49 E8 45 7D F5 5F 37 E8 9A 4D 5C
 47 FE 0D A6 A5 BF 79 4C 3D 10 1A 14 FF E4 66 2C
 21 06 F1 70 BB BA 9B 72 2D DD CD 5F B2 D3 17 E7
 0B C2 DC E7 2C 89 8D 1B 59 59 97 0C 68 23 D1 8F
 A8 F3 C3 BA BC 36 31 24 2C AF CD AE 06 BF AF 9A
 07 9E 05 82 50 DC 18 07 1E E6 8B 6D DA BC AC 37
 A0 38 0C 4C 9C 90 A6 3F B1 D9 6F CC 21 CE 68 BA
 22 98 F5 86 E0 58 0F 30 CD B6 94 52 37 F8 1D 5F
 6E DA 88 15 33 FA 2F B2 DA 1C AF AA 7E F9 44 54
 6E 04 FB CD 72 C8 59 34 26 50 43 26 AC 48 B3 6E
 35 D7 AF 80 CD 3C FD A5 D1 D9 82 E4 9A 55 E6 B8
 CC 92 A2 4A ED 65 F1 B7 32 B3 70 AA 4E 06 AB 4D
 CB 8B D6 B8 2D 93 2C C7 E1 13 0B D6 FF B9 0C 04
 27 4E E6 BF FE 46 C0 33 A0 55 8B A2 47 E5 C9 4D
 F2 29 E7 75 82 A6 7D 99 17 5D F2 D9 B2 E5 21 C1
 CE B3 12 6B A9 AE 55 86 19 84 BC 25 A9 D8 90 8A
 EC 4C 0A 49 16 A7 C5 29 65 80 F5 12 70 AA 2D EA
 BF 02 27 F9 CF 10 D1 90 B9 6B 83 57 7C C0 09 40
 DE 05 D9 42 FF 10 B2 FE 4C 3E 38 BE FD C1 15 B1
 C3 8C 84 CC 14 8A 17 B1 B1 31 3C 10 EB 5C 41 74
 F0 1F 01 7E 0E 13 73 AE FA B4 DB D0 EC A4 BA D5
 6A 20 86 D5 E3 5E DB CF 66 3D 60 7A 76 FE 03 21
 75 D5 88 72 20 32 67 A2 B0 D7 18 BF 53 43 C5 4F
 FE 40 E5 01 60 63 75 45 92 FD 59 3B 64 57 EE 0F
 A0 B8 EB C2 1B 17 E9 E4 E8 B9 18 BC 2D 02 05 BD
 0A 61 D5 E4 1A 36 21 0F D0 AC BF 7A 11 33 CB A4
 7A EA F3 6F F5 8A 1C 9C 57 60 0C 17 3A E1 61 D4
 BB 9B 90 72 1C 01 37 EA 49 F7 59 D2 BB 16 75 53
 C2 E4 03 EB 26 1B EC 4F A8 E6 A1 61 62 1C 47 F5
 02 67 EE E6 1A E7 4D 89 B6 EB 1C A4 0B DA 9B 77
 D3 CD 86 40 CA BF A5 84 9B 81 85 A1 84 CD 13 CF
 0C 5C FE 7B 4A E8 B2 53 04 23 B2 D9 3E 1C 7A 5C
 D3 EC E4 42 42 66 F2 A9 D6 58 06 26 C3 A0 EA 5A
 3F 65 43 64 79 78 49 E0 9D E1 13 A8 44 22 F6 94
 6C A5 7A F9 29 16 3D DA 64 46 12 A9 97 EE F2 5C
 49 E7 62 50 AF 43 BF AE 6E D0 73 E5 C2 9A 57 A1
 AA 47 84 6A 26 9E D4 BA 50 1C F8 A7 61 F9 E2 E1
 E4 CE 4E ED 28 A4 8E BF DF FD 44 73 22 88 5C 29
 3C 75 E4 9A 20 2F 5D A3 A2 93 9F A4 B6 54 91 73
 F8 35 CB DD 0A EC 5F 29 1D D7 DF 4C 12 B8 A9 5C
 BA 4E 7A A7 61 B1 71 D5 25 8E A3 CA 41 8A 82 2E
 DC AA 1E 01 04 47 72 B0 54 25 16 88 57 41 72 26
 BA AF D5 25 20 C9 5A 5C BF 85 D3 97 10 CD 46 D5
 B8 0B 4A BE C1 5A EE 2A 5C 60 C3 23 30 FF 53 3D
 C6 EB 26 28 51 E3 06 29 0B 25 F4 74 EC DC 70 B4
 0C 5D 49 94 22 E8 3D BF E6 10 DF 86 3A 63 8C 57
 DA 59 0A 99 BD A3 32 BB 09 5F 2A 49 CC 16 C0 77
 37 11 36 F2 EB 50 FB 28 41 0D 0F A8 7D F9 87 6F
 30 B1 DC 3D 8D 14 24 59 9A 64 07 08 08 6B AF A0
 98 0D 69 B4 C3 B8 88 4E 5F 25 40 F8 E8 A7 31 87
 37 E9 98 9D 56 9D D0 BB F1 D4 BF 6F 10 B1 C6 4F
 FB F9 F5 F2 1F 59 90 BB AC 5C 26 2E CC A5 E8 BF
 27 21 04 8D 48 37 23 0B 9C 60 E9 EE 0F 4F F3 54
 67 8C 6E E2 DC B1 61 4C 8B C7 01 71 68 DA 25 B4
 D5 AB 08 52 22 F6 DF 1B E5 41 15 C4 A3 F1 D1 6D
 AD C5 06 C7 48 03 44 6A 54 0F 73 94 93 89 BB 36
 3E 41 48 BA 8C 06 CD 05 3D D0 56 E2 D1 BF E6 8C
 3A 02 F4 05 5C 1C CD 4C 8F 70 F5 40 88 FB F7 D2
 5B 26 39 C5 0D 03 C4 F9 33 AE 8B 8D A0 DB CC 8C
 10 07 CC A1 A9 07 5F 47 7E A1 1C F8 97 D6 C3 CF
 97 78 E6 B0 B3 ED 39 9A 79 47 48 D0 E3 15 44 6B
 6B A3 3E 55 FC 4E D4 D2 AF F8 D4 24 13 81 2F 32
 2A 6A 67 9F CC 96 D9 B1 43 9E 9A 00 B7 F5 4E 04
 90 AC 54 26 A6 17 61 53 7E 3C 4C 2C 20 1F 73 E1
 AC 04 F5 4A EE B8 DE 26 9D 30 4E F6 F7 35 C2 FA
 92 61 AB 14 E2 FE 37 80 43 12 EF 89 05 31 39 B2
 9F F1 AD E8 C0 95 A2 10 57 DB FA 53 B1 D9 A0 4D
 8F CD 1F 59 00 9C 21 69 3A D2 C7 1F 4E 73 AA 49
 EF E8 FC E5 DC 4D 91 32 AE 0C 2C B4 8E 73 E7 70
 38 20 B9 19 3E F7 95 F3 C5 EA 08 36 64 26 3D 0D
 1E 9C 2C 53 8F 8F 0A 04 CA BC 08 F9 EF 73 38 92
 C7 01 AD C4 2F 0E 2D E5 16 A6 FA F1 62 B7 64 0B
 79 B2 3E 85 97 D6 DB 60 A3 CC 2A 1B 10 27 58 4C
 FA DC 41 01 03 F8 1E 0E C0 2C 8A 2A 61 AF 76 39
 17 DA 3A 0A 07 6A C3 E5 B6 BB 2B 98 9C EA D4 59
 8D EA CC 93 D9 5C 80 DC 83 1D 65 BB D9 CA 95 8B
 22 3B 08 11 C3 9D F1 46 30 D9 81 CF FD 3F 7A 4D
 58 22 00 44 D5 B4 59 CA F1 F2 99 FD 14 BF 1F DE
 56 C4 7F B8 AD BD 8B 94 23 11 43 1D ED CC 44 6D
 DC 27 12 C1 C4 55 41 B3 F7 7A 22 B8 46 50 FA 90
 18 52 39 60 AE 05 2A 98 1E 4E 1D BC 98 D0 62 94
 D3 54 74 BD B2 0C 58 9E 09 09 9A D9 9F 08 2D AD
 37 69 1B 17 52 22 D5 BD A2 8A 6C E2 1F B0 D1 3A
 59 28 40 8F C8 0D 9B 13 43 2C F2 18 6C DC 45 D7
 93 58 B1 06 7D 2F E9 F9 6B 46 12 71 64 5D 8B 97
 C6 46 59 2C D7 96 F2 38 45 96 B2 1B 33 0C 5E DE
 14 3D BC E7 09 32 53 26 CD 90 11 89 31 DC D0 2C
 FD BD D8 F8 0D C5 61 60 26 27 0A EA 55 89 CB F5
 D3 13 BE 97 2B 12 C3 C5 71 E2 A5 B0 A5 F7 63 36
 E0 FC EA C8 5E 0C FC EE 66 08 07 88 DB 00 40 26
 86 85 6D A8 09 78 4D 93 72 37 5D DB 38 BA 66 29
 11 FA A4 89 F3 72 E0 9D 85 01 77 29 57 0A BD 7B
 DD E8 F0 7B 48 10 F1 33 90 F1 E6 BA D0 CB 1A 3F
 F7 7C CA A3 2B D5 80 5F 94 7B F3 5D 67 6D F4 55
 59 83 E2 9A 33 0D C5 85 2B 42 69 B7 E5 23 76 99
 5E 1C 6A B3 ED 68 3C 5E 38 DF AA 6D 88 EE C0 99
 70 7F 36 22 9D D2 3D E2 70 AF F9 68 76 3F B2 1A
 49 21 7C 18 87 15 B0 4A BE F9 16 DF 79 9E F8 6A
 E5 9E EF BA 1C 85 E2 49 4F DC 66 D9 51 7F 7F EF
 9D DA 1F 8B A7 B9 AE 6B 99 F7 55 13 D1 23 BD B7
 95 33 B2 B6 CC DA 04 CE 1D EA D2 AB FA C8 10 FB
 AF 15 82 DB 4B 44 BD A4 56 77 06 7F 8D 57 23 39
 4F 8C 95 4B 11 AD 59 C3 BD 80 AB AB 06 FE AA 1F
 78 3A C2 C6 20 D0 92 7A C7 81 02 B1 B5 EC 5B B3
 29 58 A7 34 5A D0 07 4E 1F 92 98 19 19 EA AB D6
 F0 11 F6 00 98 FA D5 9D DD 04 9E 55 96 2C 32 2B
 92 8A 20 2D 7E D1 CD DC 62 7B 28 D9 45 E4 81 55
 CA 87 AE 30 D1 08 CD 92 AC 23 89 7B A7 C0 80 08
 1A BF EA 09 AD 7B CA FC D6 1B 0F EE E0 2B C1 F8
 F8 1D 6C 2C 58 51 5F 65 83 8F 9A 95 78 D8 02 95
 3F 36 79 9C 80 7A 8F 56 4B 4F 64 EC 0C 21 4F 5E
 C3 E3 00 A9 FE 25 EC 0C CA 10 90 96 AD 1C E9 3C
 81 3E BA A6 6F DE 65 42 07 F8 E4 84 85 42 68 01
 DD 11 C0 C4 47 26 23 EC A7 6B 45 93 6E AF 2B 82
 FB 04 12 A2 59 11 9E 85 F5 81 17 0C 10 F7 F2 23
 66 A5 AE 27 74 08 CC 62 9B 16 01 C5 40 58 E1 A5
 61 08 DC 71 43 71 84 39 FC 17 70 CA DB 26 55 1F
 2E D3 13 E6 EA 45 85 8C CD 7D 1B E2 6D 45 83 BF
 88 5D 1B 9B 22 05 40 8E 2D 07 EC 93 45 C3 66 5F
 66 7C 62 B1 A0 24 9A AF 75 8C A6 1E 21 0A FE 81
 4E 0F DF E8 4A 23 68 13 41 27 74 CA BD AD AE 2F
 F6 A8 C2 6C A8 81 FA EE 88 29 1A EC 15 C0 C0 2A
 86 F0 24 C5 79 35 E3 C1 06 C7 44 28 05 04 3D DA
 C9 4B 68 01 FC C0 D1 D6 B3 57 13 B7 0F CD 77 66
 98 C9 5E 11 B2 D4 22 15 51 AC 75 52 8C F1 FC 53
 FA 41 7F 28 D1 7F 1F 59 67 A5 04 8A 8F FF F3 93
 F5 17 0D 69 EE 04 2F C8 25 7C 0C 34 88 0F DC 04
 DC CD A0 AF 2B D0 A7 23 E1 5E DC A0 98 DD E2 54
 48 FC 17 C3 4F CA F8 7E BB 86 6A C9 BD 62 65 DD
 05 50 86 9D A3 68 BD 5D 6D D9 FB D5 3F B5 C7 63
 3E 68 DD 18 76 2F 33 2B F2 BB AA 9D 9F AE 39 9B
 39 6D B1 96 02 95 68 C6 03 AC 7D 52 21 17 B1 8A
 8D F9 B7 86 C0 33 4B 4A 8B EA 48 68 73 7D 22 63
 81 30 AF 36 A1 3B CD 04 0C 48 8C 77 29 E1 60 F1
 52 C5 C7 EA 39 D6 1B B8 97 5F F6 A2 E3 DA 40 AA
 BE F7 D3 9E 8D EE 30 A9 0A 41 AB FB CF 68 54 35
 F8 56 CC 74 6E 26 57 B7 A8 12 CB 72 46 14 BB B1
 26 F4 0E 2D 9B 7A BF 12 31 C8 01 4B 89 5B A2 35
 42 32 D4 3E 21 E0 9B 7E 61 ED FE D6 3E 4D BF 9E
 1E AF 81 58 B1 2F AC C3 76 F0 4B A2 0F D6 95 6F
 F5 8F 81 08 BA 69 AD 4F 63 71 F4 C1 FD B5 D5 4E
 89 65 4D A1 38 0E 4E 4C 81 99 B2 C4 DA EB F5 BD
 FD 6A 3E 3E 7D 4C B0 95 B3 B5 9B 71 06 14 3B 2E
 64 79 BF 04 5B E4 BF C5 D1 06 7B 4F D2 6C DA 34
 E8 9A 98 58 DB 31 23 42 A1 B0 70 90 58 DB 1A 93
 F4 66 CB 8F F1 27 BB 50 FE CB 2F 19 2D 1C 7E D5
 B3 36 2D 13 42 0E 14 F9 7A 70 40 5B 70 D9 A1 EC
 85 FF 8B B5 9B 01 72 A7 70 B4 68 67 9D 4B 47 EE
 64 C1 B7 C5 4D 87 F7 DE FC 1D 21 26 CD 25 79 DE
 22 71 56 7F B8 EA 2B 9E 85 13 96 11 69 D3 89 33
 8E D0 DA A4 DC 6C 2F E5 7F 56 4A 8D 2A 3E 64 1D
 FC 6B 14 9A 95 40 44 28 5B A7 1B C8 82 84 BE E4
 13 CA 26 D6 8A 56 B0 26 39 B8 50 E4 3E C3 7C 47
 F2 98 D1 CB 26 95 09 A0 D1 69 80 75 4D 55 53 E8
 9C 3E 9B 99 56 13 6F FE 66 43 64 DE C9 30 4E 03
 31 E3 8A D4 77 1F 2C 3E 24 3F 97 2F 5F 45 B3 B5
 5E FF CF 48 57 A0 BD 4F 08 2C B6 42 1D 18 C1 25
 41 AB 30 B4 2D 61 99 13 CE 2A 1C 93 F2 12 AC FE
 1F 1A BE 6A FD 27 04 59 49 51 42 DB 57 D1 CE F5
 F1 E8 80 95 4C F5 0F 52 8D B6 B0 D7 0A 6D 4E 8F
 F8 56 48 00 63 9F 36 BF 25 C1 63 AC A6 24 22 B2
 3D 4A E8 BC FA 67 4A 31 91 03 E2 68 98 6F 11 9B
 06 2D 5A 46 DF D5 C2 E8 12 BF EF 32 74 8D 70 10
 10 DF 34 78 7D 09 6C 5C 42 CB 17 BF CB 27 27 B5
 B3 10 17 26 E7 2F FD 3A 03 00 B1 47 48 C6 CC A4
 06 1B 43 4C F0 74 58 AD 4D D0 5A FF A9 58 A5 C9
 C5 7C 2E 04 FF 42 CE 5B 3F 73 05 C3 22 3C 72 C1
 5C 45 5B 20 E7 57 AC 00 55 0A 3F 05 97 94 6B 04
 3C 0C 1A FD 39 40 56 B5 6E DB 74 34 DC AC 5F 17
 F1 6A 15 C9 55 BB 6D 74 EE 2F A5 8D 4F 50 97 F1
 38 64 42 66 D3 BD E2 70 C1 3C 49 F6 A8 D3 70 E6
 91 2C 34 B4 99 40 50 E1 37 4B 71 13 7F 48 5F E8
 6E A8 8F 28 82 99 91 E9 30 40 0E CB 6D D8 9B 1D
 31 2C A3 1E EE 88 6A 76 73 DB 07 A6 53 5D 71 B4
 D5 48 D0 5D D8 0E E2 9F 0D BA FA DB 39 FB 88 A6
 4C 47 03 B7 DB C6 D1 03 BB 61 B8 AA 25 7D F7 BF
 05 73 8E BF 22 7E D3 6D B1 B7 18 89 B4 DD 38 4F
 40 BC 81 F7 ED E7 1B 68 58 0B FC B7 AA AD 8C 7D
 DC 57 39 B5 68 FB 36 D3 3E C9 40 8C 63 E8 5E 5E
 D5 6B 02 DE AB 72 2B D6 9F B1 30 3B 4B F3 4A D9
 16 19 4D D8 0E F1 78 75 55 99 0D 23 9D F1 7C 56
 01 1C 2E D7 B0 EF 7B 29 D4 66 38 6C ED 18 BF C0
 C3 B6 87 7B 20 99 E5 8D CE D0 6B 07 24 25 B0 24
 A0 A2 5F F0 C8 11 4D C1 D4 01 93 B9 6D C9 27 A3
 8B 42 AD 93 67 70 CB D7 DF F3 12 2C 52 16 AA 8C
 FC 39 1A 64 83 BD 2B 5C E9 37 FF 93 57 F8 60 FD
 FE D4 F5 BA 17 F4 F0 01 91 DB C8 0C C9 29 1B 33
 E5 D0 C7 20 34 14 32 B5 10 AE 0A 30 21 08 33 EA
 43 A7 03 20 6A 9E 3F 58 C1 24 FB 0C ED 3B 54 B6
 08 2F F4 5B 2F F2 A3 D7 77 EF 6A A2 8B 4C FF 4F
 25 AA 7C 49 C7 27 09 C8 BA 0A B8 4B 7B 9D BE DF
 8E 3E 40 11 74 BD A5 BE 83 F8 5A 52 D6 3A 65 E8
 E8 EF B1 FE FA 71 22 53 3C 7F 45 4A 9C 8C 18 3A
 C4 C6 80 26 27 79 23 B7 9E 57 E2 41 B0 75 B5 70
 75 D5 ED 7E 66 42 F4 79 BD 3B 86 B2 FD AB 45 C8
 0B 12 E3 BF A2 96 99 51 A6 30 EA 3A 50 31 3B 47
 AB 4C FE B2 3A 6B C8 93 E8 02 35 93 6E CD 65 DE
 28 C9 4E 98 4E C2 BE D2 59 B7 C7 4F 61 01 C5 69
 38 D5 26 2A 21 98 52 C6 2E 89 0B 35 CE BD BA F9
 EA 59 48 CA 3B 43 56 F7 A9 A9 63 72 AF 8E 48 F1
 46 34 27 8C 80 B0 78 28 C7 4D 0E 9B E7 B6 7B 3F
 C1 69 E5 E1 AB 5B 88 61 B0 36 16 EE 7A D4 2E 95
 0C CD 39 21 6E A6 85 69 EF A3 18 79 C9 A5 38 40
 4D 18 EB 76 FF AD 2A 71 96 BB DF 9E 19 89 8C AC
 EE BE E2 C1 86 7C 7F 8F 76 33 B3 B5 48 93 6F 0B
 F6 D9 FA EA 31 59 20 1E 58 96 F5 DC C5 56 21 64
 D4 35 CE 90 C7 D9 76 DC C8 F4 69 A8 2C 4B 76 A6
 66 13 B9 A3 A2 A5 EA F2 B7 4C 36 62 E9 E1 1B 0B
 CB 29 28 66 40 6E B1 82 BF 0B B7 A1 78 98 62 55
 57 C5 19 33 54 84 67 CB 81 34 51 F9 45 BE 26 0F
 22 51 4F A3 43 0E EF 3C 09 06 4E D5 FF 96 7F B6
 38 F2 6C F2 9D A8 C6 6D 71 E6 AA 37 BA 0C 98 FA
 6E 34 18 A2 2B 57 37 1D 80 E0 4A 81 D0 77 7B 49
 A6 73 5F 75 D9 56 05 A2 75 53 D6 F6 C3 B8 1A 8C
 40 78 2E 94 61 76 98 8F 1E E3 CD 4C DD 39 01 C7
 3B 8D DB DF F8 41 12 9D 6D 58 32 AC 38 1B 62 4D
 45 10 46 05 39 6B DE 63 E7 10 FA 14 86 F4 34 9C
 CA 62 9D B3 6E 32 94 D7 01 BC B6 78 3F CA 9E D7
 C6 7C 52 85 69 46 F1 E4 43 66 A8 C2 1B 72 88 A1
 DD 1F 8E 5E CE 14 32 5F CC 7A AE 33 EE 59 D4 95
 74 AC 43 71 8E 50 2F 6C BF 78 37 E1 DE 79 53 46
 14 FC 3E 8C 52 3C C7 E8 26 58 5B BE 99 5F 8F 19
 27 19 EB E6 2D 00 91 75 BA DF 68 B0 60 70 C5 3A
 78 89 33 9D DC 15 E0 19 78 79 62 A4 6E 0E 52 58
 9D 55 CD 58 15 86 FA 1B 13 C0 01 18 30 A6 6F 26
 E8 39 66 08 C7 F6 5E 16 06 06 3D 31 A6 43 86 37
 13 32 28 2C FE F5 9A 13 C1 49 06 00 D1 4A 02 01
 37 45 DC CF 2F 82 77 71 62 70 E8 90 4B CB 99 9F
 92 58 56 D4 6D BB C9 FD 0B 54 9E C1 3A FC 2C 23
 5B 04 D3 F6 4F F0 39 D5 83 22 2C 24 F3 52 56 68
 47 9D AE 2B 10 19 2C C1 D9 F1 43 87 7D 2C 1B 51
 D0 94 24 6D 86 10 4D 9F C7 BC C1 77 BA C5 7A 23
 41 6D 11 BA BE DF BF EC 87 79 5E 6A B8 76 2A CC
 D2 59 29 D7 D6 27 9F 71 FC 1B D6 4F 77 EE 02 DE
 CA B7 25 17 36 F9 61 33 83 3E 9E 35 92 83 ED F7
 FC 9E AD 0F D2 32 01 78 53 D9 47 53 68 53 44 F3
 C0 7C 8F B3 F3 D7 8B C5 56 A9 A9 20 D8 7F 67 85
 68 BA 22 B7 60 CE E4 90 18 AB DF A2 40 A1 E4 AA
 F9 A7 03 8A 80 2F BA EF 27 48 C7 A5 0F 74 69 62
 F0 26 10 E8 C3 70 AC 91 0C 7F 5F 40 31 4B 64 75
 97 BC 96 62 4C 61 C6 FD 97 0C 28 59 18 BB 0E 09
 ED 25 59 7C 14 34 F7 97 FE 85 0F 0E 8A C9 F0 82
 F2 06 D5 47 CA 98 2F 93 ED 02 BB 5E C9 F6 17 85
 EF 78 1E A7 09 B6 C8 72 00 69 39 1A F0 43 9B FF
 DB 8E C3 E0 1A 52 FE FB FB 7F E2 D7 40 E4 41 E8
 DD 3F A4 86 9A BC FF 79 06 F0 D5 4B A6 DB B2 52
 7C 8B B4 2D 99 19 66 87 B2 1E C7 46 31 B5 65 21
 51 D3 66 BA 68 46 90 8B 4B EE FE C4 17 9E A6 E7
 F6 A4 2D 8E B3 EB F9 3F 72 FF 69 2B CB 50 4E BC
 D1 77 64 23 D8 90 93 D5 FA 8C A5 83 2C CD C9 2A
 C7 B9 A7 65 CC 7D C1 39 FC 8F 2B C4 92 44 31 3F
 67 EF 91 AA 4A 61 C7 14 C0 D6 08 BF 96 6D E2 3A
 BD DB A3 75 5A 53 02 19 CD 7F 6B 0E 07 06 50 D6
 65 79 67 9F CD 2D 2E 86 48 0F 2E 88 39 E7 32 4C
 19 F6 26 48 DC 59 4F BB EF 06 22 10 17 41 66 2A
 6A F2 EF D7 3D 4A DD 60 2B F5 69 A2 C2 EF B7 18
 A4 70 9E 23 85 5E 1C 89 CA 9D 47 82 74 41 1D 53
 51 53 01 2D 9B EB EE B4 F6 D6 06 2D D2 77 95 C1
 50 4E 60 BD 81 44 8E EF DA 7B 5A 35 32 5E 50 B1
 5C 5F A1 CC FC A3 BF 10 DF AE 54 64 2A 0F A8 02
 2C 41 23 C5 5D 04 91 90 9B 3A 96 16 8C 1A 89 55
 AD 75 70 37 E5 F4 85 C7 EB 59 0C B3 B9 75 CB 69
 02 91 2C CB 26 F4 51 1A C2 0E EF 02 BE DD 7B 67
 D8 A9 0C 9D 40 01 EC B0 40 52 21 14 C9 F0 AA 9C
 25 D2 DA 03 5A E9 51 C8 24 97 E0 01 C7 12 91 C0
 24 68 D7 79 DF 90 5E F4 5B 17 0E A9 79 60 ED A6
 E5 4E 55 9C 81 36 04 A7 DC 52 B1 98 60 73 F5 50
 35 77 A9 9C F1 D2 77 58 E8 4A 68 E9 37 1D 28 93
 A5 FA F8 0C 4A F7 FF 0D CB 63 37 58 6F 4B 1A 77
 FE C2 12 2C AD 36 06 77 EE A7 67 4D C7 AC 0B C6
 97 18 62 04 99 67 3E 2A F3 3F 1D 31 F8 C7 23 84
 CB 11 D4 1A 68 4E E3 B6 6B 01 17 9B 72 9E 35 2B
 CF 1C 4E 94 BF 9E D3 DF 55 B6 23 F3 35 39 66 85
 06 42 5A FE 2D B8 7D D9 79 A7 B6 E5 15 85 B1 FD
 42 B9 07 45 95 4A A5 81 33 CF EA B8 CD AC D1 E5
 EA C4 4B 9D 41 5D 7E 84 6D B9 B2 43 54 E3 82 7F
 EB 2D 4B AE F7 50 68 9B B3 4E 83 FC 89 7D 2C 98
 B9 23 02 87 9D D2 97 A5 C6 14 6D 26 B5 09 77 2E
 AC F2 D6 31 F5 51 55 8B 5A 76 68 55 45 6F E2 8A
 A6 61 8A EC 2E 6E 8F 62 77 BD C4 F7 25 A7 7E D4
 39 CC 7A 02 DE 7B 42 B7 9A 64 01 0B 53 80 CC 07
 9C 6F C4 06 2A 3C A5 9A 6B E2 01 BA AC F0 F9 45
 BA B9 DB B1 D4 A0 E7 B1 E8 30 82 F0 3E 16 A9 A0
 DE E2 73 18 E4 89 DD 04 38 EF 5D E4 BC AD 40 B7
 52 18 0E 4F DB 63 BF CE 0A 14 6A AA F3 8F 3A 54
 BB 3A E1 AA 7A 1B DD D7 BF 08 16 9B 0C 85 43 63
 25 43 A1 7E 68 FB 86 B9 AF 8B BD 83 3C EB 48 E0
 8C 80 B6 77 2B D3 48 0C BD 4F 9E 26 E6 B3 D7 36
 D7 3C 8E CA CF E2 2B 11 83 FD 48 DB B8 C2 2F 75
 6A E2 0B E5 90 8B 1C 93 66 F9 2E 45 32 1F 8C 35
 19 7E 85 13 F1 BA A9 46 DB 9B D4 5E 6F D1 0E 7C
 88 40 D2 4A 06 1C 5A 3B EB CB 8A E7 7E 72 77 CC
 C3 22 22 73 01 07 61 2B FD 64 2F 58 B3 FF EC 89
 C9 FF 48 C1 62 17 40 DB 5D 99 C3 6B 87 1D AA 10
 16 DB 94 9E C5 14 F4 C3 17 36 8F 71 37 4F A7 75
 0E 07 6D BF CB 4E 0D 55 CB CF D6 81 DC 81 6A CD
 AF 31 B3 C7 7D 42 31 09 16 57 11 CA 82 01 11 EA
 5F 8E F2 66 2B 45 64 7B 18 CA 54 A7 DF 70 B6 D2
 3F 64 68 86 B3 F2 DF D0 4A CE 53 29 93 A1 E1 D4
 83 D4 4D 44 11 F3 B8 7C B0 62 21 4A A3 40 6E 72
 95 58 C0 C9 3D 15 BF 03 6C F9 1E A0 21 81 EF 74
 91 DB 0F 37 75 AD A1 AB 95 4A 54 9E 0D 6F 6C 2E
 68 D9 C7 22 26 93 93 6D 74 D2 0C EB B9 09 BF F8
 50 DF A1 F5 77 33 19 3B 15 98 80 94 E0 F5 C5 80
 95 24 9A A4 CE 2E 26 49 71 CA CE 8E 63 DE 10 43
 54 FC 1F 15 91 F0 86 B2 C5 BA C1 C0 5E B6 3E 58
 C3 8A 46 1C 76 84 22 21 47 94 F5 FC 43 5E 69 3C
 99 37 36 32 9A 69 0F 8E F3 B2 91 EC C0 94 C8 BF
 74 F8 40 A9 09 4F 7B E3 C1 CB 87 C2 6F 93 49 84
 C0 69 FE 40 60 11 9F 16 0E 08 7C 16 48 5E 15 8E
 E8 DC AB 31 19 A4 F9 C4 CE 55 7C 24 D0 64 91 18
 6B 16 D8 72 4C 85 FA C7 62 B2 E9 42 FF 20 61 57
 A5 82 26 50 DA C4 BD 14 B5 01 A2 04 60 E4 0E FE
 2D 61 8B 24 47 79 48 88 78 A4 81 AB C8 3E 44 BA
 33 15 07 B9 6A 03 00 C0 3A 31 EF 0A 71 D9 F7 26
 7B 9E 0B 97 6D C7 03 DA DA C4 E3 DD EC 05 13 11
 9C EF 87 68 BC A0 AF 04 E2 0F 73 1F EA C5 D4 37
 A7 F7 8F 69 B0 FE 41 FF F0 02 81 26 79 9A 27 CA
 4F FE DC 89 80 69 E8 9B 75 7B 34 DF 35 2F 43 7E
 AD 09 B6 53 EB 78 76 67 0C 5F 4C AD BA 4A CE 33
 E3 C5 38 62 E4 BC 55 6D 89 AE 2D 17 7D 6A EC 0D
 BB 9F 95 DF EF 63 F1 40 E0 89 0C 25 5E DB FD 61
 46 6B 76 DC CC A7 82 7A BF 28 1D 0C 0F 0E 59 8A
 AD 0C F6 8A A6 DE 57 68 B6 FF F2 66 FD DF F5 F3
 60 DB 42 3E 04 D5 FB B1 C8 60 FF 5B F2 E8 01 61
 E1 07 C9 C0 78 41 58 7C F3 07 3A 06 C4 27 92 9E
 44 61 FF 64 E4 84 91 8E 41 20 81 F8 21 FF 85 32
 BB B7 B0 96 C5 CF E2 74 EC C4 31 D7 D6 7C C2 92
 2F 90 37 86 07 A7 9C 36 30 B2 51 50 BD CD B2 66
 1E 3A 8E C0 CB AC 0D 8A 66 6D 68 E2 01 E7 03 AF
 9C 27 D2 31 B5 DC 4F 6E C6 FF 1F 05 B3 3F 80 14
 0B BD 7B 6B FF CD 95 F8 AF C3 D8 39 FC 19 7D D5
 C7 C7 76 86 F5 27 13 4A AE A8 6B 30 DC 54 5B 14
 76 17 10 94 6C 7E 12 29 D8 50 1D 88 90 31 C5 B1
 DF 42 8D 0A F2 4C 4F 0B 20 B0 E4 DB 22 CF 5F F6
 5D 0A AB FF D4 A2 3C 03 92 DD DA 71 5D EA 65 07
 ED 90 40 15 6B E4 DF 99 8B 8D 4C ED 0C B5 25 A2
 C1 56 7B 0A CB 1D A3 33 16 FA 5F D5 22 A6 54 51
 79 C5 C8 C3 42 76 62 26 24 E3 AB 8E 54 F1 E9 7D
 64 A4 68 F5 FD 23 9C 67 BA FD 8E 0C 74 1A DF 5F
 24 1C 63 74 B9 82 CD CB 8B CF D4 44 97 44 60 98
 F0 1B F9 AC F0 C4 FE 58 DE 70 93 F3 60 BB 52 B6
 25 F3 97 C3 62 AB C2 84 EE B9 81 D7 95 CD CA 19
 54 25 DF 89 D1 0D 07 E1 68 F0 5B 05 57 91 8B 00
 67 B4 FB 37 12 32 5A EE 53 B0 AB C4 E1 7A 2B 4E
 2C 99 99 08 49 19 29 C3 1F 7D C3 6E 35 63 44 A6
 24 43 F7 5A 16 FA FF 0B F5 1F 66 15 02 D8 65 71
 89 B0 33 19 3C 80 6E CD 94 65 F0 35 6F D7 7C 60
 B9 0C F2 03 BD 3D A2 1D 05 3A 40 AC 3B 06 C6 B0
 DC 52 63 01 CC A3 E0 0B CF 28 83 97 D5 B1 38 B5
 C7 F5 1C 64 7E 8D 83 5D FF C9 77 DC F8 B8 BE B7
 09 47 75 86 8A B2 68 29 F1 10 AF E7 44 55 37 6B
 B6 F6 02 73 A7 0F 7D C5 0B C7 0F C4 57 CB A3 B7
 58 14 50 53 9A 46 6E CC 89 04 AA CC 27 9B D4 EC
 4F 15 85 F6 9E E5 58 6C 8F 4B D2 23 E8 FC B9 36
 51 B3 E1 77 4E 5B 3B 77 F8 28 4C 98 E1 A1 3D A2
 14 20 D3 43 90 09 00 5F 84 C6 F2 F7 39 56 0F E6
 5C CC 8D 12 8A 14 3C AB 3D 30 C2 54 1C 22 96 B1
 28 BF 11 09 F9 CD B2 8E FD 58 84 F9 C8 D9 B2 48
 BC D0 BC 0D F2 24 F7 9D 89 2E 45 9A 68 7E 80 D0
 BC DC 2E 84 87 F3 5C 72 95 B3 7B 15 9C 8C 94 6E
 C5 1C E8 D4 80 68 DF E8 11 19 18 37 99 D6 2B B5
 DC 63 D1 95 50 54 48 A2 11 7F 4C EC 05 4B B6 86
 7E 78 98 54 99 65 79 9F 6E E8 99 82 14 A9 06 AC
 7E A4 BE BB 7C CC 10 BC 61 5C CF 07 A0 5B 04 80
 0D CA BC CD 60 B3 40 2C 03 28 28 0E 2A F7 84 40
 FB F8 E4 5B 17 A2 D4 F0 92 B9 5D AC F2 A9 6F 8E
 D0 D7 2E C6 0F 26 DC 34 DD 71 FA C2 89 91 D5 AC
 27 93 29 78 AC 74 14 59 9A 43 F6 3A EB DD 66 B4
 E7 BB D1 65 BC A0 E6 83 DB AD 90 3C FC 4B B1 9C
 42 FD FC 33 DA DB C2 91 EF 30 12 A3 E4 C5 32 4E
 93 38 3B 33 C2 38 EA 8E 1C DB E8 ED ED EB DA B9
 34 EF 2A 99 C2 21 FF CB 3C CE D0 25 C2 3A 3B C7
 78 F1 61 02 3D 70 FF 8D D9 BF F4 29 24 0A AE F4
 0B B7 6A 83 C1 17 D8 6E 53 3B FB 92 33 43 67 70
 DF D5 0F 59 26 CC 87 7A EC 4B 7D 54 0C 36 65 7A
 C8 8B 88 79 7E 6C 81 5D 46 A4 DE E8 AB E3 B4 1C
 1C 06 54 3A B6 1D 6F 5F 2E FC 36 D7 F9 97 C3 ED
 21 5B F5 E4 41 A2 53 ED 52 77 F1 1E EA 3F 35 00
 41 5C C5 0D 18 85 1D 1A CC AF F4 20 F2 6D 4A 23
 DF 59 A9 68 9B EC 81 69 D5 DE 9E 03 12 04 26 94
 97 22 BB A3 64 66 3A 09 C1 0B CB 5F 77 F7 CE 46
 34 FC D4 7C 44 90 BA 7E 9D 54 09 EB 38 47 4F D7
 40 1D ED 63 9F D6 08 23 7D 5A 4D A6 DB 08 CC 07
 ED 44 48 1C E9 86 8D C9 57 2A 54 BD 33 DE 74 6C
 47 B0 CA E7 27 63 C0 E9 C3 34 42 84 20 5A B9 9B
 76 66 B5 A3 EA 08 BE 72 C3 63 3A 41 75 EE 47 DB
 E4 5F 99 F0 11 C4 CC AF 83 37 28 C5 F6 BF 35 CF
 64 05 7B 2A 6D 82 4B AD 55 94 6F 99 C5 2B 49 FE
 63 A3 61 60 96 71 81 BB AA 86 6F D6 BF 46 74 68
 5D B2 CC 03 41 60 59 AD 48 67 63 11 61 23 6A 67
 7E 5A CB C4 94 D2 5A 77 49 66 B8 E2 32 90 76 50
 92 AC 49 50 EB 72 CA 3F C5 87 C6 30 32 4A 13 5B
 2C 79 E0 30 96 70 06 9F F1 8D 7E 0F D9 F3 21 AE
 BF FC 23 AA 77 12 27 56 A6 B4 E8 9C 52 69 86 5E
 2A 16 15 67 BF A8 70 71 63 57 C7 D6 DA 2E FD A0
 76 11 1B A8 10 76 30 D1 74 44 23 F0 76 B8 48 16
 CA 7D 6E 7E 7B AD B6 6A 53 FF 30 10 92 F3 BA 2E
 8D 0C 23 EC A0 C2 51 2D 2B 9A 0C D2 32 B8 93 51
 29 67 AA 1A 05 4B 42 F0 6D A3 07 BF 03 AD 55 0E
 19 6F 9E 45 22 B6 96 FD DC E5 73 61 DE 7E 13 53
 26 3D B8 EE B2 90 9F 7B 15 C4 77 7D 4B 60 8A EB
 CE D6 5B 89 B4 C5 72 40 59 8F 5E 1A 96 74 E0 B5
 40 3D 15 24 25 79 E1 C7 18 4B 66 AD 56 BD 3D DC
 18 C4 76 36 B6 D3 27 91 0B 24 32 AF F8 BA E6 0A
 A7 92 4E 43 65 1C CD 74 A1 2B CD C2 AF CE 70 CB
 8C E2 A6 58 0C 70 7A 00 03 CC 20 FD C3 70 F8 B6
 62 25 EC 7A CA C4 6E D2 2D 9F 9C DA DB 40 56 26
 94 3B 31 40 97 02 5C 06 DA C3 B6 C2 2D DB AF 5F
 CC F9 A8 14 6F E9 B6 EF 88 6D 01 8F 86 34 92 4B
 95 80 EF 01 04 39 C8 72 AC 59 16 59 48 72 84 3C
 57 D6 D0 B4 08 C2 26 C6 44 73 30 D9 E5 91 7B 51
 AE 84 E1 54 8C 9A E3 CE 84 8A 8E 44 B7 D5 06 07
 01 CA F8 9F 60 DC 98 DA 68 27 E5 2C 48 80 98 90
 27 E1 4B 56 23 8A 06 DB 07 38 09 28 98 E3 0E 91
 3B C2 D2 CC FB 2D B4 0B AF CD E3 3F 19 2A B5 DB
 13 B0 C9 74 8E EF 22 80 CD E0 9E F7 AD FD 48 8A
 97 62 EF 37 66 F7 10 AE 9D C6 CD 11 47 CF 52 52
 6C 11 88 68 65 46 4D 5A 13 72 10 A2 93 6E DF B1
 55 39 1D 65 24 77 E3 98 9A D6 9F 11 DC 75 06 85
 D7 9A D9 36 9C AC 42 5F B9 34 C2 B3 9D F2 0C CD
 B3 C0 62 C4 31 CE 12 4A 46 3E 8E FF D0 65 F1 61
 4B F9 6D 34 6B 63 C8 0A 08 21 EF 79 8A E2 70 2B
 B6 A4 7E 6F A2 CF F3 13 8E F5 04 1B AB 82 98 5E
 71 98 E8 26 7C B2 40 08 09 CD EA F4 4E 91 3E 90
 85 F0 68 B9 4E AA A1 25 01 1C 09 04 53 07 B5 9D
 DC 25 50 49 B3 32 F3 E6 E1 88 24 AA 03 7A 48 73
 59 73 F2 39 C7 70 F0 28 95 50 27 90 01 1E 67 F3
 B3 83 AF 8E 00 28 74 09 3A B8 E9 D7 6A A0 F2 32
 33 7A 08 25 04 46 E9 4F 30 AE B1 B4 AD 29 27 CF
 48 9D BC 9F EB 50 87 8A 9C E5 21 35 5D 6D 50 D3
 FC 7B 42 57 3D E7 94 5F 4E 7E 6A C2 57 26 A9 41
 C4 A9 D2 DF 4E 63 53 9E EE DC 1A DA E4 0E 25 C0
 F5 D8 33 0B EA E5 14 1D 46 32 05 2A 4C 48 3E 96
 16 BD 00 C6 C0 24 89 CA EA 9A 0F F5 23 44 66 48
 49 29 4A 49 E4 13 72 A3 72 60 7D F9 97 49 60 F7
 BE 90 2B E9 2D 52 D2 9F A9 2E 71 65 DB 3F 22 64
 19 47 88 2C 52 D4 5C 41 DD 4D 2F 0F CB BE 4D C7
 A8 80 84 D6 EF 37 EB 13 34 D1 2C CC FC 04 52 03
 E7 26 94 50 35 D9 F9 23 39 7C 14 19 CC AE 0F 27
 53 A0 3A 04 BE 8E 29 25 F8 23 2C C2 E3 92 5A 0F
 0D 38 E5 C5 73 7D 02 47 B8 CA F9 6A CE 5B 18 D7
 43 55 60 68 0B 96 DF 68 19 C9 07 C4 E7 07 06 F7
 B7 05 DF 5F 23 F7 3E 7B E5 F3 78 F5 A3 8E 43 29
 C6 02 9B DF 66 4A 0A 4C 68 1E 94 41 A8 47 19 11
 36 2C 09 70 C3 5B 09 3E 05 3E 9B 10 20 A2 36 55
 84 45 DB 52 6F CB A4 88 A6 70 0F D0 3A 3A 03 63
 84 FC F4 FE 7A AB 90 3F CA 0D 22 0C 17 96 ED C7
 7D B2 BB 15 F6 55 66 BE 6D A6 F6 28 F3 57 1C 26
 B6 FA 5F 8A E3 E0 7E FB 42 10 EB CE 1F 2C EB D2
 B6 26 14 DE 59 E4 87 95 59 FB 99 D6 10 75 E8 5B
 C2 A2 6F 0F 08 46 B2 52 8B 88 C0 7D E9 9E EB FB
 8E D6 B7 64 23 4B DA 3A A7 A2 53 23 24 43 B1 7F
 94 CA 78 E4 37 2A 08 BC FD B2 B5 82 23 42 CB 5C
 07 9B C6 15 B4 27 03 51 76 F6 AB 55 13 19 2F 37
 EA C6 4D DC DD C6 EB 62 E7 8A 5E C2 EA 54 5B 15
 B4 4E C2 31 E7 63 15 53 B4 6E A9 C4 13 FC 1D 25
 F2 E7 63 9F 07 69 8E 1D 5E 51 4B 85 FB DB C6 BC
 C5 21 7E D1 D5 F0 46 3A 57 BB 8B 77 E2 6C AB 95
 B7 3F B3 6D 78 EC F8 AA 95 23 8D D6 57 5C 2E 22
 D3 1A BF 76 ED 6C 83 D4 BA 70 7E 7E 6F 51 12 18
 6C CA 19 DD 26 FA 69 58 D1 C2 61 07 8F F7 28 D9
 F1 D3 28 01 3D FB 0D D7 F1 53 91 13 DF 82 9D 58
 29 7F 46 67 DB 70 95 DB 39 84 C7 4F 09 51 4A DF
 FD 54 93 92 27 4B 0C E5 E6 2B E2 EA 52 49 89 49
 1F 30 38 2C 11 8F 51 5C D9 A1 49 6D 80 92 6B BC
 43 64 F5 89 58 DB 7C B0 7A AF 31 9D 2D 2B 0D 5B
 69 7A 9B D9 D2 5F 2F E2 3A 45 B1 3B 2A DE 2E 4F
 EB EB BC E4 54 A8 1C D5 4D 3D 33 37 D2 53 79 25
 E4 DF 0F 1B E0 3F F2 E0 D6 B8 0F A5 92 A0 E7 92
 22 7F 73 41 C1 8F 60 03 56 05 DB 50 44 AE 42 76
 89 B9 68 C2 90 D2 F6 AE 36 B0 51 01 32 46 D2 1E
 8C 03 22 59 0E C0 FB C0 73 DC FB E3 70 76 2C C0
 78 79 0F B9 59 A8 82 67 B8 89 90 B5 09 93 90 0B
 95 F6 C2 00 38 C4 87 EC 5D 56 1B 83 3F E5 2C A5
 DB 7D B4 DB C5 B9 F4 EF CC EF 4C DB DD C3 B4 A6
 48 0B 9F 73 4A 97 8B E3 6A C7 0A 72 D6 6F F3 53
 F1 95 95 DF 2C 81 EC FC BF 70 76 1D 12 23 7A 04
 9A F7 B6 EB DA 55 FF 70 0D 07 CE 84 F0 9F 25 C9
 9D 6E 57 2F 24 24 6A DB 56 70 3D 99 D6 66 08 28
 1F E1 89 B3 2D 3E D4 21 DA 48 94 B1 16 56 72 16
 B4 D2 7A 7C 06 63 EF C7 87 42 C7 4B 0A FD 7A 48
 08 36 5B 66 14 4F 04 E3 1A 0B 12 3E 62 80 2D E0
 9F 40 E9 87 E8 64 64 88 CA 4C 84 F1 CA 55 D9 53
 CC 12 06 21 A3 99 AD EE 73 5C DE EA 9A 00 02 38
 DA 25 AF D1 D0 CA E2 7D B6 E5 16 9C F8 71 95 A3
 7F 58 AF AA F2 9A 40 B8 70 E2 59 AE 43 1F 65 2A
 10 22 A7 5C 9F 90 20 A2 D2 9C B8 3A FA 47 EC F6
 49 2C B6 E8 0E A9 1F 16 37 C5 23 0F 6C A7 E6 06
 33 DA A2 ED 79 C2 1B 39 E6 82 52 7B 08 FA DA 79
 94 97 71 F4 D8 9F 03 67 02 56 2E F8 0C 05 C2 48
 AD 51 79 4F 72 DE C7 05 64 0D EE 56 26 FD 3B 32
 78 41 E5 3A 05 74 C5 61 0B 02 4D CE CE C3 B8 94
 62 D2 83 1D 55 4F D0 6F BB 9F 1F 76 80 0F CE 13
 07 44 01 F0 51 8D 3D 46 55 CD 7E D2 18 E3 47 FD
 B0 2B 56 EF 78 10 8F D7 5A B7 F4 CC 9E FD 33 FA
 7E 4B 32 B8 4B 3D AF C5 0E 64 07 56 66 8A 39 90
 32 C7 05 24 14 19 9B 99 6A DA A0 77 07 4A 54 67
 97 28 F2 68 D7 EF B0 EF 39 28 FB 11 1A 16 FF FB
 49 18 41 30 7F 49 13 7D 4D 4E 47 03 73 8D 45 EF
 1F 2B 56 FE E2 9E EA 6E 3A 37 55 EF FB 04 01 BA
 C3 73 0A 55 74 89 68 B6 9F B0 0B 49 F3 51 6E 9D
 BA 1F E0 DF 62 8C 3A 7D 68 6D BB 0A 04 24 0E 3B
 97 AB 39 BB 03 87 34 C4 59 91 40 B8 09 BF 38 F2
 57 F2 9D B4 4F 80 EF 6A AB EA 7E 70 E2 88 6A 76
 BB 95 1D 81 88 5B CC D6 34 7C 0B 95 24 D7 3E C0
 D7 3C C9 6B CC 34 83 EF 68 C4 CE B9 A1 87 3A BC
 D8 9E 2C 0D DC FF 9A 04 30 5C 42 9D 97 60 D6 D2
 17 E7 24 90 4B B3 E7 75 7D 38 25 BE 50 1B EA 01
 86 29 65 9C 3D 57 F5 E3 E3 90 D7 B2 23 B6 1C EC
 87 2C 46 01 FE B0 88 19 20 90 19 45 1E F6 D2 BF
 9E 14 09 EC 6E 85 A4 42 57 26 CF 55 9C 4D F4 AB
 1C 91 5A FC FC 30 AB 4E 22 9A 14 B1 8E 02 C4 E1
 30 B4 97 5D 81 2E 84 50 C5 95 89 30 07 33 C0 3C
 B8 D5 25 9A D1 8C 3A 0B FA 57 49 21 E4 EA 8A DA
 08 C4 15 F3 43 98 0E 68 6A F7 4D 67 5E 2C 78 A8
 77 D8 16 18 21 2A DA 6D 85 70 79 0B 10 41 17 F9
 26 97 88 DB F7 DF 3E 34 7B 11 99 18 E4 AF 8D 39
 8D 90 1B 8E 3F AB 56 C8 7D 11 DA 54 56 91 5C AF
 B6 80 03 6A 3B C7 30 B5 C1 CC 49 EC C1 24 2B C8
 CF B5 09 02 28 E4 EA 27 82 D3 59 B3 AF C5 9E A8
 5C 17 B5 BC F0 D1 47 A9 91 09 B4 F2 79 92 B7 26
 25 65 D8 DB 6A 40 AE FB A1 C9 93 4A 76 2A 6C 51
 68 F0 49 2C 71 F5 4E 0E B9 9A 4D 9F D2 EF 67 54
 E3 EB 66 56 FC B7 FF 77 15 19 D9 2C E8 38 86 20
 F9 0E D9 E0 87 A5 72 16 27 1B 06 01 FE 67 13 2C
 9C 2B 95 5E 8F A6 D0 C5 0F 8F 7A 0D F2 E5 8D 54
 DC 65 CF 92 65 C2 E7 C0 6D 8F 28 D1 D5 14 B4 A0
 A6 26 0B 6F 19 35 33 97 DB 59 A4 E3 76 F9 29 6D
 57 25 D2 3B 7D 05 7E DB 37 56 18 D5 CF 90 EA 61
 70 62 32 0C A2 B6 64 5E 65 50 9A B4 46 D8 A2 76
 26 62 8D A4 4C 01 AB 3B 68 F4 79 9C B3 4C 6D 82
 17 79 52 D2 BD 25 FF F1 C9 23 B0 BE 11 11 47 96
 71 6A B5 F2 17 2F 4C 19 25 F0 A3 27 97 B9 2D 3E
 1D 47 B4 AC 2D F1 1B 98 66 FE 77 69 0D 94 67 3A
 8F CB C3 BC 2E AF B7 69 07 20 A8 1E B0 01 5C 27
 7A B1 B5 C3 3D B1 83 C4 42 CD 0D 3E 4E 9D 0D 53
 C0 A5 19 BA 95 B8 C0 88 32 04 AA FF 82 38 3E F6
 4F 19 04 66 D0 76 0D 68 E8 84 A5 F4 8B 98 1A FF
 50 11 6A A3 9E 20 80 B0 2A 1E 80 ED 18 52 E8 12
 C1 32 6A 7E 32 23 DA 6D 65 10 9B D9 26 BC 8F 6D
 5B CA C1 A0 E0 BF 53 AF B3 53 F6 1D 49 97 33 04
 26 11 7A 7D 0B 9C 27 E2 A7 1C 66 8B 69 35 74 B8
 A6 79 2C 86 BF C6 83 6B F6 50 D7 EB 92 D5 65 75
 F6 C3 16 E0 CD 5F 8B AE 4B 8F A1 5D 2E 13 ED 88
 DD B7 3C 43 8C BA E2 27 7A 63 09 E0 77 B1 B3 29
 B9 60 B5 8F A0 22 3D 50 35 96 DC FA 7D 9A 76 EC
 A3 C2 BB 94 43 3F 8C 33 B8 FC 0B AF F2 80 7B A6
 07 20 92 F9 B8 34 B0 BF BA 8C BA D7 8F 31 05 74
 4F B6 1E 3D EE 9C 9A 75 8B AF 93 C8 F8 F0 31 E6
 84 20 D2 4E C0 BC 52 C2 4F 7D 47 EF 34 71 DC 68
 93 CB F2 02 64 E8 B0 BC 13 2C 3A 70 28 11 62 E3
 F5 4B 79 56 82 35 A9 8D 66 DE 0E D0 3D E3 48 1C
 5D 57 A2 06 11 B8 51 3C CE 4F 30 AC 58 F8 BA D4
 C1 A4 BA 5D 4F AB 2B B5 63 9C 12 56 A5 85 30 4B
 80 06 BA 9C AD 78 69 EC 0F 59 41 28 09 86 D0 CA
 83 32 36 10 24 1E 10 DF 24 9F C4 37 C9 E4 F7 33
 D9 92 E4 05 A7 BA FE 6F F0 39 0C 10 7B 38 5E DD
 02 71 87 20 5D 63 2D 27 9A 63 04 AB 34 20 AF 0C
 12 1C A0 4A EE 0E 56 3E 68 F4 33 BE AC 1F F1 7E
 69 38 AA 04 7C 56 21 69 96 5E 76 02 A5 E6 67 72
 A2 8D 31 2E 70 A3 CD E0 FC D4 C3 6F B1 91 1D 76
 86 81 3C B7 6D 1F CF 13 A5 EA 01 0C 8F 5E 0F F3
 9D 91 22 CC F9 CA 37 0C 5D D7 0D 94 7D BC A8 C6
 6A E9 F1 E2 2E 43 DA 66 B5 CC 11 BE F1 F6 0A A4
 9A 96 81 CD ED 88 7F 71 BB 5E 0D 23 59 52 5E 14
 D2 44 A9 26 27 BA ED F6 D6 4D 77 6E CA 5E D5 49
 51 D8 50 09 24 F9 5D 4B 3B EF 72 26 22 FB E2 C2
 DC EE 4C 50 45 00 92 59 27 2C 47 E7 3F 73 5E 9D
 A5 58 ED F3 5B 15 F9 F6 49 92 D7 1E 2C B6 E2 87
 55 5A 31 19 52 03 6E 56 9D 38 40 0F 63 DA 1A 0C
 FA AD 2B E7 6A 03 15 EF AE 54 F6 64 A6 B4 96 87
 86 08 CD 6E 02 6E D0 6B 8E F8 90 86 16 E8 44 99
 84 5A 8F DA 79 C0 BF 49 C2 C5 46 9F EB 9A 80 EE
 4F 0B BD F1 97 88 C6 FA D1 DB 00 4B 94 71 C2 AB
 96 B2 9A 97 2B 58 20 61 A7 14 47 BE A1 70 FF B7
 CF CF 38 6F A6 8F 15 BA 33 F5 52 B5 34 A5 BD D2
 49 DE 13 1A 23 BF 94 81 64 FA 1B 51 97 93 AD F1
 C8 A2 67 3E A1 88 5D 75 A1 A5 8E E4 4A 6B FB BF
 B6 F8 F1 D4 25 B1 EF CF 7B 7B 96 E4 D4 97 8F 03
 A1 9C 8A BD 66 7B 0B F7 F5 F6 98 09 27 AB D2 1B
 B4 16 81 D0 02 65 6C DF 0F 04 37 70 D6 7E D7 02
 84 B7 A0 89 AE 6F 29 EA 08 BF A9 34 36 85 4F 77
 6F 04 C1 E8 AF 32 D2 54 73 01 24 DB EF E7 DA 08
 B4 FE 11 BC 51 02 D4 4F 43 E6 B7 8C 4D BA 63 44
 C0 38 3A 68 6E 07 36 3D 84 17 16 D8 87 55 09 12
 AD 42 02 E3 FC 84 48 AD 75 DD EE D9 74 59 A5 BC
 67 82 CA 84 81 CA CC AC 80 93 52 5D A1 CC C7 75
 45 3F DA 69 CC E0 E8 84 47 E3 78 F8 39 BA B5 14
 AA 23 11 58 FD 1B 18 AB 9E B9 16 1B 7B 46 99 C7
 53 D3 38 11 BC DF 4C 55 08 33 00 E4 6E 9F FA 72
 02 C5 1A 7D 91 44 95 B6 C1 4C C1 2D AA 5E 15 18
 0C A9 E4 27 17 57 D2 0C A8 80 BA 2B DD 8A 76 BD
 48 77 3B 73 DB 74 A7 42 A6 8A F3 81 63 84 F7 E3
 83 EA 14 BD 1F FC 48 30 66 11 6B 02 62 6B DD BF
 2C DB D2 D0 A9 E3 C2 60 09 51 1A 91 A8 5D D7 8D
 3F 1C C5 44 FD 04 F3 67 73 AC FF 75 14 FC 58 34
 A0 3C 7E 86 71 E6 49 43 51 B4 69 37 C7 19 C3 D9
 C3 8B 4E 8B 19 29 F9 22 53 F6 15 B8 F2 92 4A DC
 AF DB 00 01 E6 7F 07 6B 69 AB 67 A1 4F 28 14 63
 BF 0D DE 72 CA 89 90 4A CE 68 34 79 CF D8 8D E2
 86 75 E4 A4 38 2E FD 9A 7C 75 9F F0 01 BE 16 D1
 45 2B 7E FA 58 73 88 AC E9 F9 B9 F3 DC 67 F8 B5
 D1 94 D8 E0 33 7F 6F 2D 69 4E 94 39 5A A5 4E 09
 47 1A 3B 86 4D 9A FC 8E B5 D3 F4 D0 67 1F 97 7A
 13 D6 51 F9 C8 54 7B DA 7C 2D 14 5C 84 05 CC 57
 AD B6 20 64 69 8B 67 8E 2D D2 A1 6F FA F4 FB 50
 16 AF CA 95 47 97 19 28 D1 8D 6B DB B5 D5 B7 6F
 F4 EB 7D D2 D6 93 C0 9A A0 CF 08 58 F1 09 14 E7
 C0 CA 65 27 D6 20 AA 12 46 D3 4A 79 BF 67 F5 5F
 31 1E D7 22 2F 60 9A 21 1E 8F B3 6F 14 4D 07 7A
 DD D4 E9 19 30 5D CA D3 20 FD D3 35 69 8B 7B 03
 9A 57 7A E7 A0 0E 93 2B A7 34 BA 79 E0 1B B6 ED
 67 C2 A3 54 E0 EF 6B 17 50 1B 58 EF 66 A7 DF 1A
 6D 31 BB BC E4 4B FC FD 9F 68 3B 3F 8D 9A 7C C7
 8C 1D 2B 4E F9 C2 80 E9 CB 00 EF F6 86 C7 10 12
 E0 EB 30 D6 E5 17 50 E5 2F F0 89 0F 4B CF A0 6D
 AD 07 D3 E9 FF 56 29 8A 57 BA 15 18 57 65 5F C5
 27 D1 86 A7 75 3A 6A 3C F6 DD 0A 61 13 26 1D AF
 F0 07 16 B4 7D 73 F4 6C 22 29 61 03 62 F2 78 09
 FD FB CE 59 85 84 AC 13 9B 16 7F D7 BE 5D 7B 95
 EA D6 CA 31 F1 00 15 7E 08 66 E7 43 58 70 B2 A0
 4D 68 47 FE 15 6E C6 68 2E E3 34 46 DC 28 C6 D2
 BC 22 9C C0 F1 0C 14 CB 7A DA 50 C8 58 D7 40 9C
 60 B9 FC 4B 99 94 23 49 88 51 B4 8D B5 27 69 11
 1E 66 B7 EB AD 95 AC F2 44 53 DA 37 EE 5A A1 07
 17 99 DC 11 27 4C 75 F9 01 0A 0D D1 E5 84 29 7F
 84 BC 4C 6A F9 60 7A BC E9 86 56 06 65 3C 4D 23
 7C E0 3A D9 0A 2E BB AD E8 D2 77 76 1F 4A 09 23
 B3 BC 5B F0 62 A4 57 A8 EF 06 C9 C5 49 95 64 C3
 C6 50 3A C0 58 A3 01 9C 26 49 06 C6 36 C2 1D 2A
 4B 39 81 06 13 AB 52 55 27 31 61 6B A2 E6 24 AD
 FE 56 3B AF 5D 3E E3 91 34 F2 8E 7B CA 53 B5 43
 6F 55 16 2A B8 A1 82 12 00 22 BA 98 60 42 1F 02
 3B 2A 29 DA 98 03 79 2C 60 B7 88 07 25 72 A9 89
 D1 DF 09 56 10 1A 4F 91 89 FA CD 47 68 B9 99 09
 D6 73 BA F8 74 21 A6 1C 88 E8 35 7D 76 CA C0 9F
 B6 BE CD CB 91 A8 13 43 64 4D 1A 42 40 44 D4 B2
 EB BB C7 65 38 FC BD A4 6B 7F C9 33 AC FC 40 85
 13 B1 76 7B AE 2E 16 76 F0 32 0B 30 D3 DA BC 36
 56 71 EA B1 3B 1C 56 ED 54 8A CD 19 30 42 BA 10
 4B 8D 60 0C F3 E0 E2 82 89 1A D1 74 22 65 A9 D4
 B0 5E 04 0E B6 A6 B9 BD 8E 49 8B B4 1D F2 58 A4
 FA 65 6B 5A E5 AB 22 27 E4 CE B3 F8 26 FC 33 06
 70 51 AC F2 2A BF E8 39 A0 58 13 94 BD DC F1 81
 12 90 00 1F 48 21 B0 D0 C7 18 79 D5 CD 21 3B 2F
 28 4D 1D 7F 66 1B 01 44 66 C5 F5 36 90 E4 F6 BC
 34 10 4E C0 4C FE C9 0C 22 F3 64 60 30 22 7F BD
 E5 04 93 83 AB 5A 30 E3 12 EB A9 F2 ED 7E 52 DB
 83 1A 14 6B 54 BD 63 7A A8 A0 FD 30 53 F2 22 91
 FF 84 6C 20 A3 76 2F F5 57 45 29 2C 08 C3 28 FA
 91 43 49 C6 80 54 E4 F2 29 B8 A3 D4 C3 21 20 BA
 E8 51 A4 FB EF 48 B2 4C 31 1A 4F 5E DE 96 10 A9
 15 93 83 EE 0C 1A 2D 71 79 83 10 BC 8F E4 3D F1
 5F 35 AE 61 41 4A 1F 80 04 AB 63 D1 55 4E 5D 13
 2E E9 8F 09 A5 12 B3 EC 16 3F 8C D8 6C 6D 7F 6C
 26 F2 32 08 E5 16 18 D6 D6 A3 B6 4B F1 05 C4 2F
 05 5A D9 E8 0E F2 27 58 5F 09 0D 2E B4 A0 08 ED
 2C E0 ED BC 52 52 20 87 B8 47 DD 10 4D 5C D7 BE
 03 1A 68 A6 5D D8 A4 AB 26 97 0E 2F 04 3F 08 39
 92 26 0A 43 E7 51 88 B0 38 64 56 BE D6 7F CC 43
 84 81 DB DC 3D 27 73 A0 F2 D6 4D FC 4F C9 6D 8A
 EC 9C 13 0C E8 CC 80 99 78 2F 95 B4 BE FA 71 C9
 D1 6B C4 B1 18 48 4F D9 85 1A 64 CC BF AB 2D 75
 F8 3F 87 E8 C6 5F FE 3E 67 1D EA 45 30 5C D2 D8
 0B 5F 9A 22 2F BB AE 90 28 C7 9F 27 BC 1D 58 70
 F8 A3 4D 5B 61 26 EA 87 5E DB 2C 1D 61 CB 85 2F
 08 8B 4D CD 89 9B 74 87 CD 4E 4D 86 1F 36 03 4D
 F5 77 5E BC D6 F5 B9 B7 09 99 63 A9 C5 1D C0 C7
 C8 7D A6 EB E9 99 60 9E FD B7 6B 22 24 3D 2F BA
 1A 9C 03 28 96 F8 4D D1 4C 49 E5 88 3B 7A BF 46
 6C BE 05 22 B8 3D FA 21 AF 2E 17 B3 F4 B5 35 FF
 AF E5 82 FF 48 D5 7D 3A 11 26 1E 14 52 45 CB D4
 A6 1A 76 1B 1D 27 C0 83 75 33 2F 4E F8 E0 1A B8
 3A D1 D2 F7 32 48 8A 20 4A 89 CC 90 42 1C 78 7D
 D2 FC B4 D1 EC 79 5F F6 34 AA FB 4E 7F F7 46 C4
 24 46 A3 98 9E 23 88 23 9D 5E 2B 5B EF 9F 3F DF
 2F 7B 35 36 96 EB CD D4 F1 06 0F B5 6C C7 DA 84
 C7 7E 93 FD 01 70 6C CB 5A 3D 2C 7D 94 92 57 0D
 27 75 59 14 CC CF 37 79 E2 6A CA 27 F8 D6 71 55
 A4 A4 AE CB 63 B7 28 33 AE 7A 54 6D FB 69 49 74
 C1 14 20 75 03 2D 38 4B 25 B4 B5 CC 38 27 1D 84
 85 4A AE A5 DD 19 59 DD 21 95 32 19 92 B6 97 8C
 DD 2C 46 97 25 51 79 0E 99 24 5E 25 5C 11 D8 9D
 6E 72 FE 61 19 4D 6F A0 A7 A3 D3 D8 6A DF 26 99
 72 E3 09 5F 6B E6 5D 55 A1 CF BA F5 89 67 6F 8F
 33 56 26 0A 7E 15 0C D4 81 48 52 E1 7B E3 15 76
 E9 D9 85 5F 99 AD 31 28 B9 78 8A 8E 07 4E 91 8E
 BE 6F CA F2 FA 76 94 C8 AA E6 E9 38 A1 42 D9 19
 D2 E0 C6 40 46 76 80 55 22 2B 9B 3F E4 49 8D F2
 D0 EC 8F DA AC 46 D0 30 89 15 A4 B2 0F 8E F3 62
 CF 0D 16 39 BA C7 10 43 38 DE 98 9B 9A 0E 58 B3
 E6 AE 93 19 67 23 8A 5A 1B 61 2D AA 4B 63 19 E7
 C7 EB E1 2C 39 40 55 9E 42 42 D7 BA F9 60 51 50
 A8 CC A5 FA 92 F2 35 18 2C B4 E0 8E 2C 6A C1 BC
 7C 5C 35 3F E5 14 C7 A9 D6 DA 6D B4 6C 1C 33 28
 B1 AF F4 9E EC B1 BC A7 79 75 9D 52 57 52 69 C3
 1D 5C 64 64 D1 BE 8E A5 D4 20 3C 62 2C B1 CA D5
 E0 DC 75 DA DB 37 97 D6 5E C1 41 59 4F 92 B4 9F
 CD 40 65 1E 35 BB 3C F0 28 FB AA 9E 02 86 BA B9
 21 5B 6A 36 20 6E 53 47 CA DF D3 39 0E FC 2A 86
 4F E4 3C E5 90 91 EA 90 68 12 AB B9 19 3D 9D FB
 D0 AF A7 10 3E A1 74 3E 1B E0 3F 5A 86 1E 87 DE
 DB 7A 0C 38 1E F2 8C D5 F7 FA 42 7E 9E 9C 45 A6
 5A 25 75 6F 2A C5 C5 F2 0E 38 D6 11 C2 EE 8A 96
 A7 08 FE 56 C7 7A 1E CA B1 C3 9D 35 8E D4 6C BF
 3E FD 0E 36 3B 2C F0 B8 C0 B3 D8 9C 40 29 70 6C
 3B 50 32 EE E4 89 18 06 15 E9 EC 8A A1 41 F9 EB
 6C 67 DC 91 F8 46 22 81 F4 43 64 AD 3B A7 20 AD
 88 EF 43 29 68 6D FE 8F BA 90 A9 77 D0 6C 49 67
 D5 85 9E 08 98 DA 73 AC 77 03 8B BA 12 32 EC 23
 3D B5 50 20 BB 33 E2 F9 C3 5A BD D0 D2 5C 06 A2
 94 0B AF 56 9E 41 E1 91 80 F3 25 ED 67 3D 12 A9
 30 68 66 D8 7E D2 B3 DB 6D 0B 97 E6 46 7A 1D 2B
 1B 3A 74 8C 67 A2 B0 B0 DD 30 69 FF 07 75 AB BF
 EE 6B E7 FA 2F 6F 54 E5 7C 96 96 A7 E3 30 65 6A
 40 60 AF FB 31 C5 D0 F4 52 C7 1E C8 E3 67 52 5F
 20 8F ED 60 5D FC 7C 5A 6F 09 BF F3 D6 05 7E FA
 82 B2 35 C7 5D C7 1B 93 29 80 23 5B 73 6C 10 A3
 0D E5 F5 F2 42 C4 C9 D1 EC 4E C6 1A 22 74 AE C3
 4D 37 67 15 4D 65 26 FD FF DE 39 C0 64 D5 E7 7B
 B7 24 13 D0 9D 16 46 32 79 51 68 35 5A BC 32 19
 20 B3 B9 CA 3F 7C 56 11 02 6D B3 7F E0 6A A2 49
 76 D5 3E E6 37 31 5B 92 84 2A AE F8 7B 5E DD CC
 C0 45 89 39 1D CB 20 24 64 71 D5 B4 04 BE C7 32
 F0 71 FB EC C3 83 48 2D ED 10 95 73 9C 56 3A 10
 5A C5 BB B5 5A 84 24 27 65 C9 45 29 C0 DA FF 5A
 0E 08 9A D2 59 C6 9C F4 FE 91 71 D4 C5 72 2C 77
 0A 65 3D E8 CA 9E FF AA 08 39 AB 8B 23 BD 86 CF
 B5 4F F8 24 E0 08 DC 99 D4 E2 FC B5 DB 26 D9 6B
 B7 E1 3E A6 4A D8 E6 77 64 A8 01 47 C0 7F 9A F7
 78 D2 DC EC 4A E8 01 23 65 D3 6C 01 8F 06 EE 6C
 B9 C0 F2 98 4A 11 77 11 AF 12 D9 7F 1A 83 C9 40
 9A BA 63 90 25 E6 B7 26 C7 8C 12 0A 5E 23 3D A5
 0C 6D 20 51 BB 85 72 43 FB 24 14 EB C9 C6 52 E9
 39 D7 55 21 49 4A 49 B3 25 70 4D BA 07 6C 05 A4
 0D 02 3E D0 08 37 36 02 39 C2 0E 74 F8 83 37 E8
 E8 47 6E 52 B7 19 1A 8A A0 2B B5 27 F2 06 D2 69
 64 A6 0C AF 95 D8 C6 DA 13 AC 88 05 B2 02 2B 65
 EB 0B 83 06 ED 8C 50 E2 35 F6 74 77 53 62 A1 89
 E5 CC E1 97 EF 67 4B A6 06 4B 0B 01 4E C7 9E 18
 AD C8 E6 DA 7A 5E 2A C9 2C F8 A8 FD 89 63 F3 BC
 9D 7E B3 71 11 3F 3D F5 D0 36 3B 20 73 9A 78 73
 AE 80 5B E6 AA F9 E8 3D DA 57 F3 74 EC 6D D4 55
 A6 86 F8 BA 13 10 31 65 E4 1E 32 6B 68 57 EC C1
 1E B4 A4 FA 60 6F 14 18 C1 F2 A9 04 33 DC 95 9A
 5A 95 4B D9 E4 BB 1F 4D 7B 31 9D 4B D0 C8 1A 46
 53 7B 91 2B F4 48 C7 EF 64 0D 2D C0 B5 AD 76 68
 93 D0 55 17 D1 C4 33 85 B0 F2 3A 53 F9 E3 09 70
 7E 6A 82 3B 98 00 13 CD F0 74 2D 3B 76 90 8F 8D
 7B 33 34 3A AB 28 B9 56 6C F0 40 6A 5D 60 F3 FD
 AD 40 09 C7 AA 9D E0 06 29 90 71 FC D4 53 D4 06
 1E 50 A8 6C 4C AC 7D 64 05 83 04 E1 EB EB 97 04
 6E 0A 32 B0 47 E3 65 78 99 C4 0E 0A 4B 45 CD 7D
 3F F7 6D 32 A6 C4 54 2E 8D 42 7E 12 39 28 8A 56
 04 0D 4A 60 54 10 AB D0 7E 7E AB F0 53 32 19 96
 CB 11 2F 07 4C 78 9B 8C 86 0F F8 DD 75 40 5C 75
 F9 71 D0 5F 2F 5E BD 70 DF D7 77 5C 03 CA D8 DE
 08 C0 16 7D 52 38 04 16 EF 97 AB 64 16 5A ED C0
 4D 92 A1 8D C9 18 69 30 3D A8 5E 17 D9 9C 68 F9
 6A 0B A0 D1 4B F2 4D 30 23 DC 12 44 7F D5 10 29
 92 6F 15 2C 75 E3 BA 6F 33 5B 6E 85 0A C0 21 4A
 46 CE 44 CC 89 1D F4 FC 65 D5 5E 25 C5 67 31 B1
 5B 1A EB 79 D4 BD 44 BF FA 0B ED E6 96 0D 12 48
 89 6B 98 23 F3 8A 12 86 DE BB E0 94 AB E3 2D 8D
 84 E1 45 E5 48 C4 B8 8C 56 97 35 7F C7 82 E3 EB
 B9 01 66 DB 32 94 05 CC 0A B2 F0 2A B5 63 B9 12
 BF 69 43 78 0F 66 6B 06 DD 0C 61 81 3A 0F 51 B3
 9E 96 EC 1F 72 98 4F 01 EF 75 C5 8C 44 B4 B5 3A
 04 57 F4 40 EE 0C D6 0F DF 56 63 65 AB F0 2A A6
 17 9C 8F A8 7D 51 F2 80 A4 AB 21 07 87 AE E2 46
 4E 4A B1 B6 05 70 1A 6D 5B 7E AB A7 F3 9C 21 60
 8D B2 C1 FF E8 41 D1 F4 FB 16 39 56 A7 48 F5 FB
 8C 82 3C 7D 75 72 4E 29 45 95 6B 8A 7C 69 F8 2B
 86 8D 66 B3 A0 0A 3D B6 2B 77 B9 BC F5 90 BF 7F
 E4 A7 B6 5D A6 66 DE 69 52 CD 7C 34 0D 97 FC A5
 BF 8C 3C E7 25 47 F7 5C EA D9 1D 45 BF E3 5A BE
 8C F8 AB DA A9 CD 53 F3 95 25 23 48 25 0D 21 1D
 0C C0 1E CE A1 6E 58 07 21 89 9B FF 18 17 6B B1
 12 AA C0 48 6A CF 6E EA 65 81 49 15 93 7A 05 DD
 28 70 A5 4B 23 27 05 3F 92 11 97 18 68 24 2E 7C
 97 5D 29 5F 45 20 55 46 6E D0 A8 6E D6 50 BE 3D
 3F 35 82 4C D6 95 C1 57 03 6F F9 0B DA 12 7E 1F
 43 4B 8B EC D7 4F 78 91 A3 AE 26 2E 08 01 51 39
 3C 21 C6 A1 2E 82 BA 57 8C 10 03 97 87 7E 36 21
 12 4C 0A B3 90 5C D4 8F 7D 5E 7B E9 FA 0C C5 16
 D2 55 7F 89 68 15 0C E0 B4 FC 70 27 8F A0 96 F1
 B5 BA 54 FE 56 DF 13 43 20 A4 91 03 48 34 D7 32
 27 FA 95 6A 7B AD 3A D7 44 CA EF 4E C0 40 A3 C7
 4C E6 23 BA 1F 88 DD F8 9D C7 91 EF 58 DC 1D B8
 6B A6 5C C8 D6 15 3C C3 8C 7B 18 CC 25 1C 5B 73
 50 F7 71 F3 AA 79 EF 80 5C 0F 42 2A 0C F9 7A E3
 47 57 09 3E 02 E5 39 6F 9B 10 21 68 14 C1 28 3D
 C7 B8 D6 BD 61 6E 85 8B F0 6D 44 91 10 D3 1D 62
 53 87 5D FF EB 66 CE 3F E4 79 57 53 EA B6 BE 7C
 CD 0F EA A6 09 06 C5 9F A0 0D 2C EE DB 46 A9 5C
 B9 B0 B6 A6 0B 91 48 D7 7E 89 53 90 E5 F9 B0 F3
 CB 6D 68 61 A4 C6 76 AD BF B2 62 B4 AC 1F 11 F4
 3B F0 8C AF 68 24 F5 7B 5A 1B 05 AD 6A 3A C4 E2
 2C CA ED 87 E9 77 CF 81 08 26 1D BF 16 B5 3C 48
 B6 50 04 73 C4 80 61 9A C6 BE 99 CA A5 77 FE F4
 49 AD A8 2B 98 01 8A 25 0B 68 E0 68 49 D6 B1 9B
 8C 4B FC 48 C8 A7 47 1C 47 3A 24 9C 16 BA F0 E3
 3E 72 BF 99 BB EC F9 1D 13 48 25 6E 61 3C 71 6A
 09 6D 37 C6 D8 C2 B8 39 DD AF 58 A7 3F 20 35 3B
 D7 EE 5A 7C 67 21 C5 DE 7F 9D 05 2D 60 7F 7D DA
 97 FF F3 BA 9C 55 8E C6 5A F5 1E AF AD 8F BE 68
 98 91 0C AB 9B A0 02 C8 FE 4C A1 3E 75 6B 0C 88
 09 7A 85 F9 2B 1C 5A 8E C7 57 6A 5C FF 9C E9 9B
 31 1D 2E 14 A9 41 08 4D 46 B4 A8 9D 08 48 C3 09
 4A 3D 3C 1E 40 1F B0 F6 FE A5 71 18 6C 81 F9 7F
 82 68 46 40 A5 C0 2F D7 7D BF B3 23 9E BF 14 96
 8D E0 92 CC B8 75 CE 13 27 62 07 51 F3 1E C4 DA
 3C 99 54 30 2F 76 9F 90 20 73 B2 FA 0E 35 EE 2E
 9F 9B 47 F7 C0 0B 0E BC 44 57 30 05 83 1F D3 D5
 3A B7 49 3D 95 0C 68 0F BD 9C 91 FC 4D 68 66 9D
 31 69 94 36 70 40 FA 5E 8D 45 20 08 FC 67 B8 4F
 E2 27 A3 E4 D7 DD 63 F7 EF 93 22 05 C7 3A 40 0D
 9F 94 81 41 CC E6 20 09 3F FE 4E 39 04 9D 75 4D
 82 D8 8F 80 3A 4F 82 59 9E C7 81 F6 96 ED 8C C2
 D9 22 6C 1A 91 4F E1 52 50 A0 52 96 E8 5F A8 3F
 7C 84 43 BB 08 C5 35 AF A0 F1 44 92 42 8F D8 80
 33 3E 70 5F BD 1A 3A 9C 18 A7 AC 4B D9 40 27 57
 7F 38 79 81 CA 4E DC 24 6C 76 B1 AC 91 E7 15 1D
 A0 A1 2A C9 14 95 0C 67 FD 26 D2 29 D0 8B 8F A1
 A1 B1 53 3B 8E 3C CF 63 F1 20 37 04 7C 52 21 BD
 65 E8 CC 38 08 67 79 29 1D DC 10 A1 10 A1 2F 8E
 B5 5D 94 FA 01 6D 9C 75 7A 43 D2 DD EB BF 3F FC
 06 C2 14 1F 4E 41 44 71 28 95 10 87 E6 2D F9 4C
 41 0C D0 67 D0 5F A3 E7 E8 A0 46 1A A8 3C 55 3B
 39 1E 55 9A 0C 73 8F F1 3A CF D4 86 BA D1 37 20
 2F DF 4B 1C ED 41 13 7E 22 A6 C6 15 17 FE B9 88
 3F E8 2C 6B AE 4B 62 D5 5F 66 D1 77 37 B3 7E 46
 92 A3 5C 7D A8 01 72 EF E5 2B 39 6B 00 B0 81 22
 D9 3F B2 7F 58 9A 90 E2 6D 3B 95 9C 86 F6 36 F9
 E5 E9 E6 79 E9 C0 5C 23 68 4C F3 36 2A 27 57 8C
 96 71 AE 48 55 7D 23 44 BF 3E 10 DB F5 7A AA 7C
 FC 31 00 5F C2 C1 A4 71 C3 C0 F3 4A 3A 46 51 57
 B5 2D FC 32 2B 10 C0 F7 F6 CE 04 A4 93 C6 57 3A
 E2 0F 45 C0 A1 54 3E 08 AF 51 E1 3F B8 A8 E2 39
 10 D8 00 F6 FC 90 8E 30 1A 7A DC FB B6 9B 61 B8
 E6 F3 91 FF 01 D4 51 17 38 44 5E 28 E9 33 02 C2
 1D A9 C4 4F 82 7B B4 44 14 2B CE B7 66 E2 AB 73
 1B 8E 21 C6 17 11 01 1E 42 DC 62 37 B3 EF E4 78
 6C 12 54 71 37 E9 82 64 9F CA AC E8 BE 83 AA 15
 78 8E 0B 28 43 81 5C BF BE B8 BF 2E 90 09 B3 EF
 B1 A9 7D 02 78 E0 E5 C2 8F F1 66 E3 08 03 97 90
 60 94 0A 14 93 1C 77 A0 C9 05 ED B2 BB 91 1B CC
 B4 2C 06 EF AF F2 87 E3 C7 A9 96 73 28 52 5F 18
 8F C7 F5 E0 02 D0 2F BC 25 D3 AA EB 11 45 75 63
 1E 72 BC E1 EF E4 3A 87 FA C3 E0 F1 EB 8D 58 E6
 D9 AA 7F BE B3 18 99 D8 D5 F2 1C 7C 31 14 D9 02
 6F 0A 86 C5 2C A6 FD D3 35 78 47 02 9E B2 49 CC
 FF 63 91 A5 28 27 36 30 12 AD C2 25 DB 65 AE 81
 69 6D F3 E7 DC E1 3E 47 08 DB FD B9 EF 71 D0 E3
 8F 09 31 83 38 07 5A 38 35 49 82 5F F4 05 4C 01
 98 CF 0F 47 E8 31 A6 BB 4F 56 49 92 9A 8B 15 A0
 9B B8 C4 0C 22 0C 51 8C 3E FA F3 8D 6C FB 00 FC
 E2 DC 96 8B 7D 76 6C 08 BA 32 8A BF 3A EF 5A EE
 5B 89 5C 44 AB A6 C0 76 11 EB 36 CF 5A CF D4 03
 93 70 07 A5 16 C7 89 D4 73 A9 32 0D 53 94 F3 7A
 20 7F 4F D6 17 FA 0A B7 CA C8 20 CB CA 62 63 0D
 F9 BE 68 16 79 1B B5 44 E6 3A DB 4C C1 2D 3A 71
 5E 8E 3B 7E 78 11 92 BC 96 7F 6D 62 6B DB D1 27
 34 C9 B7 A3 52 A9 53 A1 D6 80 10 72 59 2F BD D1
 F9 7D 9D 0B 92 04 B7 F9 61 40 73 1F 58 C6 00 4F
 71 24 10 43 15 01 B1 F9 A3 98 A8 87 7F D7 2D 01
 71 6B 86 12 F4 4E AE 46 75 2D 3E 21 44 36 04 A0
 9E F6 84 46 0D C6 AF 06 F9 9C 67 BC 2E 28 F1 C3
 E2 8D 75 4D E8 E7 91 54 5F 99 1F 42 32 C9 04 D1
 9C 47 44 C1 45 34 5E 35 A3 3A 2C 98 45 8E 2F BC
 48 92 6F D5 75 09 A7 A7 BB 3D 7E F8 72 62 1D 4A
 C5 E4 46 C5 FD 6E 24 88 A4 34 B1 C8 9A A4 FC 55
 92 D3 E0 65 8E 4A 67 21 CB 4A 2C 8B DA A3 65 92
 30 AC A3 60 63 2A F5 AE B6 A3 C3 41 FB 72 F0 F0
 83 70 29 0A 4E 0D AF 19 7B 9B 7F EB FD 3F C4 11
 2B 69 D5 D3 13 A8 BE 56 F4 A7 FE 0B E7 77 A8 34
 AA FF 7F 2A 19 E1 0D 0B 5B FE 80 03 A6 DC B8 A3
 A2 52 4F 02 E5 18 44 70 60 B2 1E F8 4B 44 B4 ED
 61 15 08 2B 20 F4 E6 57 6B FC DC 16 C3 6C 1D A6
 B3 9D 4E 0E 3B 7C E0 C4 FD 97 FF 65 A2 5B 7C 42
 4C 03 97 AD E5 83 24 56 AD 7F 84 7C 55 43 44 3F
 9A C3 74 8A B2 73 98 78 E9 41 40 AE F9 26 43 C5
 65 D9 78 A3 45 49 76 03 3C 44 0B 2B B6 39 64 D9
 50 35 C5 7B 2B 24 1A 35 5D 31 5A 70 C6 59 CD A6
 39 FE EE 67 70 8D 87 7F 33 54 28 DE 90 D7 CB 20
 D9 C2 67 BC A5 96 98 70 36 DF 4A 8E 53 63 BE 2E
 70 B5 FC 50 F1 43 DF 33 A3 7F 93 FF 21 FC F8 91
 1B 66 98 DD BE 22 EF A2 01 E7 BB 64 89 E4 21 C5
 E0 71 F4 82 7D 01 65 A9 81 22 73 1F 27 AC D8 6C
 BE 5E C4 C1 59 3B 82 EC 06 CF 45 CF E1 B8 7F 4D
 24 69 E5 E9 7C 29 F6 9C 3B 35 7A 47 E1 0C DE 0A
 1A 31 D5 D5 76 2C D3 5D 29 DA 55 98 F1 5B C9 AC
 96 57 52 BC 02 7F D9 89 13 B1 E6 B8 5C 4D D1 C8
 BA 47 D7 E5 41 5E 7C 94 33 63 6F E7 1A F6 E3 7F
 11 BE 9A C5 8B BA B0 96 BD FE B9 F6 2F FF 53 6D
 2F DA 1B A8 AC 5E C0 B7 32 A0 79 97 1C 8F 84 CD
 5E 0C 8D D0 7B 44 7C A8 B1 5E D2 9D 28 08 42 C2
 7F 07 94 93 4D 71 07 5B 7B 44 C6 44 28 26 F9 52
 87 80 1D 1A 64 E4 1E 95 65 37 06 60 BB 4C 24 3F
 96 F1 CD 98 3D 96 91 65 72 E7 5F DE ED 00 13 2D
 3C B4 5A A1 75 3B 1F 81 B9 26 9A CB 5C 04 2A 9F
 36 F5 CA 5F 11 77 47 CF 82 54 7F 5D C1 88 A5 80
 69 86 A5 D9 C0 D5 22 E3 20 62 FF 1B 9E 87 E6 BB
 96 B2 BD B0 BF 67 8B 4D 54 E7 00 11 5D 5A 5A 98
 AA 54 BE 5E F0 D7 10 75 8B 41 9D B0 23 57 ED 08
 E7 31 7B 44 80 C1 66 75 2A 30 45 29 82 9E 21 6B
 49 38 43 65 9E 68 7E 4E CA F3 5D 04 2D D2 45 92
 A3 C7 DA 32 50 EA 62 34 04 31 2D 5C 81 EF E5 64
 8B 4B 36 D1 D8 AB 3D E0 D3 13 E3 A6 56 72 21 FB
 9E 97 0A 9F 9E 99 6D CC FD EE 17 DF 73 7D 56 5B
 CB DF B8 89 0E 8E E6 75 EF B2 D3 A0 AF F3 EE E7
 58 0C D0 05 9B EB 17 72 15 E6 73 20 9F D7 04 FC
 92 1F AB 4B 1A 8C 68 13 8D 41 EF 66 2A AC 0B B5
 6E D1 FA 87 15 A4 EC 90 8E 7D 3C 24 BC 77 59 BC
 02 64 AC A0 CB 17 73 BE E0 0B 42 80 CE 69 00 EE
 21 4E 39 85 21 51 47 E7 40 D8 F7 7D EE 68 78 A2
 CD 83 19 1E 95 05 E6 2D ED 5C 08 4E 44 B3 6E 07
 77 4E 92 BD C4 AB 07 B9 78 BF 0F 76 13 5D 75 61
 96 ED 2D F6 45 CA 5D C6 A1 92 49 F6 DA 29 F8 F7
 60 A3 04 E2 42 72 C8 B2 25 7F ED 27 9D 31 4E 85
 FE 50 CE AF FE 7A C2 49 03 78 05 61 44 DC 95 87
 E4 4F FC DB CC 20 49 E5 C1 48 CD D8 DA 1B 78 C5
 D5 72 09 1C B0 AC C5 EF 90 18 7D AC 2C FF D2 F6
 CB 83 0B 27 CC B8 62 F9 D3 15 67 F2 DA 7B 67 6A
 CA E3 DC 1A 0E 31 CC A9 31 67 CA 7C 7B E8 24 5E
 58 80 ED 08 56 87 47 C1 52 12 FB 12 09 8E C2 16
 23 25 22 93 B6 56 55 8A 57 73 F5 42 2B F6 11 E8
 B6 08 4E CD 7D AB F8 50 D9 8D 68 45 3A C4 B1 CB
 85 80 8A 5A 34 33 77 7D DB 98 91 E2 C0 E1 A4 D5
 43 E0 A7 F6 12 D0 A9 92 BE 50 C5 F6 BA 52 5C 73
 4C 6B 48 F2 79 D5 62 0C A2 1A 35 5E DF 69 47 B6
 9C D4 EC 76 B9 7F A4 2B A3 E3 53 75 AC 00 90 86
 A7 2A 3F 75 0F 56 EB D4 E8 A3 CD 31 D0 A0 7B A5
 17 9B 53 C6 01 6C 07 AA B5 09 8A 57 FF 85 4F 07
 16 31 AC 3F 82 67 16 8E D7 DE 63 4D 0B B6 1D 8E
 A5 28 F4 B2 44 07 1D 9C C7 A1 B6 7D E5 61 43 12
 4B B9 61 BA 7F ED A9 EF A2 7B 68 B3 FA E5 A3 86
 10 14 16 FE 41 56 78 02 46 94 57 60 7C 16 8C 90
 F1 8C C5 8E 02 FB 20 B0 52 C8 C8 A6 38 74 7D 6D
 F2 FF 9F A9 D2 85 01 C9 E0 01 36 CD 2B 7B A7 C6
 F2 FE 3E 6F 83 70 6E 1C 8C 73 AB 4C 4E 76 F9 18
 54 69 94 39 A4 D7 88 71 EB 30 4D 12 74 BA 8C E2
 20 F5 29 68 01 C4 FB 6A B1 7E B1 DA A6 77 1C 97
 73 5B 09 AB 54 27 1E 53 C7 3B D7 DC 51 D9 CC 93
 07 30 C8 75 87 03 01 AE 63 F6 43 CB 3E 6C 09 B0
 2A 0F C3 34 63 D4 7A DF A6 3D B4 E3 6D 39 05 DE
 EE 90 D7 41 54 D4 3A 46 1A 5A 2A 37 3D 6A F6 01
 72 EC 2C 06 B3 7F 71 D0 9C 14 DE 5A 85 FB 93 5D
 E1 3B CC E5 51 22 ED 0F AA 2E 11 E9 70 3E 56 B2
 13 CE 5B 59 02 ED B0 A1 1F D5 8C A6 A1 28 10 3A
 3A 82 67 4B 38 E9 77 31 EB 3A B1 F5 8C 6D 08 4F
 38 63 E3 02 B3 BE 38 83 90 7C 22 40 0D 11 86 A8
 F5 A5 A3 D3 E4 21 03 E4 19 4B 99 C3 01 37 64 92
 95 4E 82 F5 6B 4E DB 41 E8 E8 D5 C9 10 38 7F 4E
 B5 D9 CF 43 6F 11 57 6F B5 D8 58 6F E9 FC 64 F1
 85 91 B7 A4 5A 27 A0 5D 35 B2 D1 A7 31 DB 15 3C
 10 E3 34 23 02 0B 2A 61 2F 9A D7 08 DC 13 03 87
 78 21 32 38 74 35 B6 5E 3E 69 B1 20 32 D6 E2 C2
 4A 25 47 32 51 F5 80 0D BD B4 31 A5 A5 58 04 B4
 D7 F1 7B CB EF DD 2B B4 58 40 5F 5A 51 5B 7F 07
 A6 B0 9B 7B AF 8B 85 6C C1 F8 3A 04 91 05 42 F5
 5C 58 EF 45 74 E5 F3 4A E3 0C A0 C8 97 2F 7D AC
 D3 A0 3A 00 24 AE 51 93 E7 AA 6E 8E 59 BA 16 9A
 D5 27 2F 22 89 35 6B F8 13 2D 6A 85 36 3C 07 8B
 8F 2D 75 D4 1C 2B CD CE 8D C1 D2 25 54 48 E5 68
 A6 A5 FA F6 2D 1F 94 E9 26 38 FF 71 44 39 EC 8F
 09 C1 2B 05 09 0C 00 E2 D6 59 6C C6 A2 02 77 E6
 76 78 12 A6 28 B3 1F 54 1F 32 A1 D7 61 4D 79 72
 AF 53 A4 80 E4 8A DF 99 42 75 00 11 A3 A4 01 54
 8C 43 27 0B 78 C9 78 DB A6 DA 53 B5 17 DF 2A 7D
 24 EF 35 6B 53 BD FF 19 D4 66 0E 7D F6 77 EB 03
 7E B1 6D F1 87 C7 27 E1 A8 4E CF B8 1E DC FF 89
 52 B8 68 4A 31 EC 03 8B E5 B5 45 35 F2 E8 C4 D1
 C8 2E 75 32 DA 79 7B 56 43 19 A0 68 C8 21 61 06
 1D B4 B6 69 01 7E AC 21 80 48 A3 07 02 EF CC 99
 EC 2C 89 1E 06 3D B0 5B 4B 4B A5 EC 93 5E 85 30
 28 64 1F E2 F5 CE 23 5A 5A 21 43 2A 3E 62 EA 83
 B7 B8 53 16 26 8D AF 9A 1E 40 B9 95 F7 D8 23 09
 96 51 A3 50 DB B3 AA A6 76 AA EA A4 03 BF 9B 4B
 9E B6 66 74 16 62 FC 9C 81 86 82 49 2C C9 76 9C
 C8 94 05 58 99 F9 D4 50 37 8A 2A E8 39 DF 17 26
 20 24 29 B6 CE 12 76 6F 39 DD 8D 82 DE A6 5C 86
 C2 53 71 C8 77 7D 57 67 34 2A E5 A8 AD 88 17 0B
 C6 2A BD D7 F0 67 1D 0A 10 69 08 B6 E7 C4 8B DA
 CE 13 D0 35 FE A2 FA 7E AB 0B 31 57 A0 12 D8 B1
 CC 0A 6B 93 41 B0 7A 1C 29 39 D8 10 7B D8 9E 0A
 5B A1 79 1A 80 B8 33 BB 7F 41 22 B2 08 A6 03 28
 7D 7B 32 E7 4C 61 79 A8 6D FE 56 F4 10 C1 24 C4
 41 A0 52 F4 E7 4A 27 1E 33 C5 B0 92 81 5E 05 72
 25 B1 BF 52 58 33 F0 7B D7 A9 07 7A FC 6E EB 70
 E4 B2 E3 E1 9B AC 14 D7 4F 95 09 89 4D E7 C6 A9
 A6 01 AC DB 63 04 8C F0 90 1F F7 C0 BB A8 A0 84
 36 5E 65 0C 81 8D D4 D1 52 9C 08 D2 32 43 4C B8
 81 DD 74 6A EB E1 5B DD A5 32 68 3F CA 1B B2 47
 1E 1E DE 93 28 DA 5C EA 5E 7F 48 14 F8 99 33 45
 61 09 CC 77 30 B3 44 01 52 62 20 DA F5 D5 5A E4
 C1 52 80 39 E2 7A DB 59 F9 56 A5 61 BB 39 D2 07
 E6 99 98 26 BB 43 54 3F 2D D7 07 0E 48 B2 4D BD
 53 85 F7 FB 50 C6 17 07 01 3E 6B 23 3D 77 07 5B
 38 23 28 9E 96 BD 3A DF 10 EA 0D FD 18 8A 57 7C
 EC 31 22 11 1C 13 C4 56 D6 46 77 57 F6 1C 9B 23
 52 09 91 79 34 D3 25 98 EF 88 9F BF A8 83 0D 48
 34 06 5D 21 66 EA 49 5F AA 09 3E A9 DA 3F D7 65
 2F F1 AF CA F2 42 F3 1E C4 7A 8E AD 51 A0 C8 C7
 94 C4 C8 6D 63 EF E0 AE D9 38 8B 8C 61 27 61 92
 A8 BE C7 C1 B6 DD 4B 10 5F E5 28 AC 9F EB 04 34
 DB B9 7F 45 7D 49 6E 75 A4 FD 46 BD D3 37 10 37
 F5 70 1C 38 4F 37 36 39 8F 81 5B 5B 7F D7 C2 41
 F3 E4 4B 4C 5F CE F8 5B 27 8B BF 38 33 5F 6D 69
 2F 1F 96 71 C7 C7 37 7A 74 16 75 1C 48 02 FA 89
 C3 66 70 42 50 09 4B 25 07 DC A0 7B 16 4B ED C7
 81 F0 A0 43 F7 AD 26 BA B4 DB E7 74 95 3E 2F 3A
 8A 8A 7E C5 EF 01 DD F9 F0 F0 81 EA A7 19 07 97
 54 73 28 23 EA CD B0 64 30 18 2E 69 AE F4 8D 27
 FB 3D 11 76 CB 88 EE 6F C7 34 3D 41 A0 94 D3 A1
 C4 59 EB 0A 0E 81 87 A2 9E 82 80 4D CF 82 4D 2E
 D0 09 D7 05 65 A0 51 B2 55 7F 92 EA B7 DB 58 E0
 B1 63 C3 E5 1F D8 83 41 F6 2C 70 2D CA 8A 63 AA
 0B 96 65 9B 8F 4C 58 19 62 02 82 2E 00 87 9D A8
 4A 67 41 85 02 43 EB 75 67 EF 63 B8 41 B8 1C 38
 66 9A BA 43 5B 4F FB 85 7D 2E 36 50 D9 85 48 B5
 C2 C7 38 FC 6F CB 16 67 DF 30 E4 88 33 E1 0B A6
 48 63 E9 19 A6 C4 29 5F 3E 70 E1 A4 2A F8 C9 92
 E8 42 AC A7 AD 16 DF 32 E3 DB 8C EC F6 4B D6 84
 40 3D DC 2C CD F3 96 54 EE E5 F9 F8 15 45 CD 7D
 F3 87 AC 1F 09 5D 3D 46 54 64 A0 20 BC 6D 8E 51
 3C FB 81 E2 E8 B5 08 5B 62 0A AE A8 9D 9F 3F 0D
 B5 EB 44 16 A6 B4 08 D1 CA CF 65 28 87 92 40 1A
 54 73 0A 7F BE AB 37 68 E5 D2 60 8E 55 03 F3 CE
 C0 89 AD 67 BA 5B 78 25 0B 57 BB 1D BD 51 4F 5A
 93 FC A9 4F 6B 74 3C 65 6B 43 D9 4B 5F E9 75 CE
 E3 C8 C6 61 E6 AF 52 E2 31 E1 A6 CC DE 7E 3A 9C
 AB 31 EA 56 ED 48 99 F0 69 32 43 B6 00 97 4F 86
 33 57 58 33 71 35 E7 99 C5 52 81 45 4F 60 D1 DA
 F5 D1 A9 61 74 E0 6E 64 3C 27 2E 08 15 6D E2 E3
 80 4E 89 8C 2D 5C 3A DB 1D 4C C1 BD F4 F0 54 5E
 99 4D 84 D3 FF 59 47 8A 3D 9B 34 5A D4 EC 25 E9
 DF E8 81 EC 86 A0 E3 D2 B9 E7 FF F1 C7 8F 04 0A
 E1 14 73 85 A6 BF 0C 72 84 3E A0 4D A3 81 A2 19
 C6 FF A1 BE 63 2D B4 A4 2D E6 C1 99 3B 60 93 CB
 68 10 BC BB 5F 38 61 20 D6 67 53 F5 1D A4 5F 3D
 A6 D8 41 26 50 FE C8 9E 97 78 46 7C 3B 63 E8 99
 1B 8B DD C6 B9 FC FD 61 11 79 9F 35 44 2E 4F D0
 50 41 A2 82 9D BE 91 FC F1 E0 E1 C8 47 E2 73 98
 A7 F0 C2 AE 7F 8F 08 AA C1 50 C6 3F 5F F1 6F DF
 E6 1A 0E 51 0B B6 3A 94 D5 03 86 B3 5C 3D D0 D2
 C5 4C 6C 8B DD 05 F2 C2 F3 40 FE 21 48 7A 32 5B
 70 AD D3 B1 CF 43 59 23 FB DA C4 E0 E3 F9 93 CA
 83 09 E4 48 08 F7 CD 6F 47 F9 F4 25 2D 20 75 BD
 0F 27 1F 38 61 13 DF 7F 49 B8 62 61 78 44 5E 15
 45 DD 2D D6 F8 4A E6 4D 60 3C DD 82 46 30 D2 3E
 68 3C 4B 19 7C AD 44 B5 D4 00 36 00 71 AA DE FA
 9C 56 6C 27 1D 0B 7F E3 36 F8 DE CC 46 3F 1A 8A
 46 9C 00 BB 00 83 AF 2B F3 C5 23 40 C0 66 9E 06
 C9 D0 3E E8 36 B0 57 D6 87 74 72 29 D2 78 79 55
 98 46 BE 3F D2 BC 98 FB D0 7A A8 F6 FB 7C 1F AE
 9A 6F 3F D5 B4 F3 95 7D B0 B4 AF 74 F5 19 45 55
 7C 3A 5C E5 6D 99 0B 90 97 BF D6 58 41 08 4B DA
 06 E6 19 2C 98 CA 7A 8A 40 09 93 78 57 7E 5D A3
 CE 8C 72 92 3C AB 54 92 FD 88 E2 A6 C5 E0 70 AA
 0E C7 2E D3 88 DB D5 17 A7 38 B5 69 38 37 2A F4
 9F DE 96 56 B4 07 54 FA 9D 61 C3 1D 8F 72 33 69
 57 63 95 2D 41 1D 96 A6 E3 E0 32 77 F8 D7 3E B3
 D0 B5 28 68 6F D6 FF 6C 63 20 80 E7 DD 78 D3 FF
 B0 81 A9 E9 38 11 F6 E9 B0 6C 5D 83 23 50 BA 52
 EF 56 C2 5C D0 1A AB A6 FF 2C 4F ED A8 4E DD D3
 4E C7 93 F6 26 31 65 26 7A 89 52 EC 3D B0 30 3F
 C3 59 4F 1D 5A 9C 90 DC 50 B8 89 F1 B1 D7 95 2B
 4A B2 D7 6B 26 CA 64 9B 85 76 2E 2B 7A BA BB BD
 EB 0C 72 F4 D4 2F 38 64 57 FD B2 F2 4D 1E 60 12
 95 05 45 EA AC 6C 8A 1D 79 81 52 1C FF CD E5 B8
 60 5D 03 63 F2 BA 28 F0 4B 10 77 85 DD 3D 42 4E
 62 2F AA F9 30 8B 96 25 2D 54 2C E6 AA 98 EE 1D
 41 BA F8 58 72 AC 43 E5 F4 1D CD B6 F9 BD B2 C0
 C8 27 0D 55 53 81 21 FE 74 9B A9 88 8B BA 3D E6
 FE 26 1F 40 56 63 DE 05 C1 05 84 5E AA DA 52 07
 CA B5 35 F6 EA 16 8D 99 A6 AA AD 35 19 D5 84 5C
 7C B3 45 A3 ED 39 80 19 4C FF 8B 23 1F 07 9B B7
 FB F0 8F D6 64 CA B2 AC 87 AD 16 47 94 6C E1 9E
 73 C8 7D A1 7F 9C C2 56 EF E3 75 FC FB FC 91 4B
 2B 80 59 25 18 FA 8B B0 38 BF 05 C0 E1 C0 F7 9C
 40 74 48 6F 4F 7D 0B 52 4D B4 7F 4B 29 EA 9D B4
 42 97 E5 58 ED 1F C0 89 40 2F D3 17 C2 2A 58 E3
 2F 43 20 97 00 AE 19 63 77 0A 04 81 88 06 70 D8
 50 DA AA 8B 0F 77 C1 C1 30 15 F2 BD 23 90 74 AE
 B4 98 74 54 00 1D 30 6B 05 4D 8C B5 21 DF 1D 37
 98 B7 89 09 D7 92 40 C9 2B A3 DD ED D7 66 2F 5B
 55 7B DA E1 1E 92 0A 2A 42 75 EE F8 F3 88 AD 27
 3A 78 69 2C 83 D2 B3 45 37 EC 63 AD 40 22 91 6A
 A5 26 C3 4E EF CD 43 DA 4C 5C 9E FB 5C 89 4B 8F
 4B 60 0F 4C 1D 5F 28 83 71 7A B5 36 AE 11 60 67
 94 70 6A 42 68 D5 8B 22 48 26 E0 1A 97 3C 6E 67
 F3 55 7E 42 4B E1 91 E8 1F 61 24 46 B2 50 E4 DC
 47 4B C6 34 C2 39 B2 48 72 1C 3E 80 03 AD B3 3E
 18 84 DF A6 06 D6 BA BD 47 07 3C 2E A3 A3 62 F0
 10 66 FF E4 70 EA 3A D8 4E 1E 88 0F D5 10 48 6F
 08 2A 0C 4E 3E D3 95 8D 59 57 D8 50 6A D2 D1 F5
 A7 CF 11 C4 D1 96 E7 B7 1F 8E CE E8 10 C0 B1 D3
 2E 29 4E 2A 37 BD 77 55 4B 87 45 4E DB 90 60 64
 9E A8 44 D4 A4 E6 88 F7 80 11 80 FA DE 4A 41 7A
 63 B1 20 6C 16 9C 19 EF 78 85 F3 A9 65 56 2D 6B
 7E B1 5B AB 3D 52 1F 79 D2 4D E1 F9 19 2A 2D 70
 9E 2A E0 5D 31 8F DA 21 92 21 61 F7 47 3B C5 BF
 D7 7C E9 9B 35 74 E8 84 17 6D 32 14 78 51 C3 CB
 C2 21 01 2A A9 86 C7 5B 77 A8 25 7D BA B5 BC 1E
 B1 70 49 B1 0B 75 52 8D B3 9E 03 72 5E E0 19 50
 C0 69 F9 57 C0 96 F1 20 32 7A 8D C9 D6 0D 11 C5
 7B F3 A7 5E 40 B7 4A EB A8 10 BB 63 61 B8 5A 8B
 B3 FB E6 BB AC 45 0D 93 25 A7 39 1E 1F 56 25 05
 51 F8 CF EB 34 0D 83 AD D5 2B 15 EA 13 5D 2E 68
 96 05 32 7B 1E 10 B6 93 9A 66 F1 97 76 B3 66 5A
 61 9D D4 C7 51 F8 EC 73 E7 05 7F 8A 08 05 86 2E
 5E D9 BB 2C ED DF C5 FF 60 4B FE C8 77 9F C0 07
 92 BF 2A 37 BB 4F 74 5D C4 B3 C3 74 72 ED F0 2C
 84 10 AA 6E E4 DA 40 E0 76 B0 57 B2 8D 34 EA DB
 4F D1 2C 6A 92 0E 1A D5 86 A2 3D 58 B6 BB 8A DC
 6F 6C 1D 25 FE A4 89 46 86 38 2B 67 9C AF C0 46
 F5 4F 51 2E 14 9F 9B 4D 8A BA 9D 14 83 31 C2 8A
 31 6A D0 40 65 1F A5 9E E1 84 A2 06 6E FC FE D2
 82 D9 5A 35 F9 0F 36 8F 7B 2C AB 58 09 E0 64 51
 D5 32 6D A5 64 A8 A5 22 E8 C7 0F 46 CF 82 EF 61
 D7 82 61 C0 45 F4 5E CA 42 27 4F E3 F1 48 75 A6
 36 D4 89 42 08 E0 C4 DE 35 35 45 AC 2A BC DE 8E
 CA 67 F3 5E 78 28 F6 7F 6F 38 2C F4 96 5E 2E 1A
 15 5C D7 2C E6 A1 79 DB 74 2C CC DD 8F 4E A0 E5
 B9 5B F6 1D C8 BC D0 68 D7 10 3E 33 9C D9 E6 3B
 D2 84 C0 97 23 E3 6D C7 F1 FC 6F DB 2A DC 74 2C
 05 AF 7C 5E E2 DD C9 21 D4 02 42 09 02 0F 89 58
 AC E5 7D 61 60 D1 FC DC E3 3F 5C 5B D7 86 42 F2
 6D 44 FA 8A 56 10 17 C0 5E 8A BE 76 87 11 30 87
 58 14 2E A8 A7 25 19 34 D4 9D BB 42 FB BC F9 E5
 0C D5 C5 B8 08 BE 2F BE 76 07 74 33 6C CE E6 59
 F1 BC B7 A0 83 F9 85 9F 12 DF A4 D0 EE F6 DC 28
 AF 6C AF 3C AD A9 A2 7A 3E D8 8B 4C 10 FC 9C F3
 88 47 43 C9 60 FF 3A F0 FD 8F A4 C0 1F E6 0E 32
 17 2D 81 D2 A1 34 91 CA 8F 67 7C 6A E8 87 03 A2
 2A 54 A5 A0 09 16 7F 6C 3D D4 8C 17 DE E1 DE 43
 89 E9 98 31 A4 31 A8 47 4F 2A D2 EB B9 00 33 2E
 5D FD FE 69 61 7F 2A 8B 56 A1 A7 85 95 E9 F3 E9
 F0 66 8B C9 88 CF A6 10 24 3A A1 0D E5 CF D0 F4
 B8 72 3E 49 13 0D DC 07 3C F2 EC 3E 78 63 ED BB
 AB A6 F1 11 CD 01 1B A8 00 B6 12 AB 50 98 0D 61
 5B C5 C2 7B A7 AC C0 9F 71 1C 1D 5E 0A A5 F6 C8
 0A 75 BC 3D 17 08 24 1A 37 EC 6B B6 02 BE F1 7D
 01 43 32 4A 71 B8 D3 C0 21 BD A9 2B 97 7C 41 D8
 84 15 17 44 BE A9 F4 1C F3 CC AF 84 56 3E 10 D8
 15 C3 D1 0D D8 55 C5 58 7E C7 66 C6 35 82 E7 6B
 A7 3C 22 CB 66 BC 6B 95 FC 53 13 47 65 4F 6A 1F
 D0 39 D4 C6 AA 27 33 E0 77 97 38 B9 18 48 34 31
 58 CB FF 22 5E B2 A9 6D 64 E5 23 C2 2E 6C 0A 46
 05 F4 FE 9D 9B 27 EE 55 58 86 62 E2 D1 94 E2 9D
 12 25 A1 17 1B 0B 76 C9 F9 2B 00 5A 80 D6 74 A7
 16 5F 66 4B 22 7F E3 60 4A 32 42 B4 11 52 FD 05
 02 CB AA 94 35 AA 22 8F 40 F9 AD 40 D2 60 39 BE
 FB 7A 02 D1 53 20 37 19 5C 63 61 BA 26 AA 58 CA
 B6 95 DA 58 1D 75 BA FD 7C 65 6F 5C C6 9F DD A8
 5D 3C D9 AC 1D C9 53 50 F1 BF 5A 19 F4 CB 24 8B
 BA 78 39 04 3B 48 A9 15 7E 8B C8 39 63 19 F6 07
 D7 65 7F FC 64 EB DD B4 3E 0C 24 19 76 1A AA BD
 04 9B E5 36 C2 DB AD AB 44 79 FC 33 A9 D3 42 0F
 DB C7 CD EA 14 4A 2D 27 4D BB 7B 3D 9E 54 06 D8
 E4 C4 8E BE CF AC 0A BA 8F 2E 89 CF 11 EB A5 5B
 5B D7 C6 CF 85 1B D7 15 32 2F B2 40 DD 6E EB 60
 F2 83 15 09 59 50 59 0E 58 25 BA 7C B4 77 E1 3E
 56 D8 EB 6B EC 23 4D BD 1B 08 A2 1D A3 9F 19 DE
 FE 6C AE E1 DB E5 F7 DB 74 D0 D0 38 BC 25 8C B1
 14 0C 6B 12 E0 60 28 05 15 71 DF 8F A2 82 94 EC
 E6 7D 9A 74 62 00 17 7F EA 6C AA 66 B4 B3 A5 9A
 CA E2 B4 F3 E8 F0 0C 36 12 3B C2 CB D3 0F E4 1B
 ED 93 F1 C8 06 35 40 89 FF 20 43 5D 59 99 31 50
 33 7D 20 06 39 09 04 0A 81 21 17 64 54 DB 86 41
 F5 54 FE D1 D6 47 92 DC 04 04 AD C0 08 FB 73 FB
 D6 B3 94 23 09 1A 92 18 EF 44 38 53 CA 5F 49 5A
 EE E3 22 06 5F BA AA EB B3 AF 5D 2C DC D1 2C 3F
 F1 1B 60 FC DD 30 0F D0 1F 0F A0 AF C3 98 2B 86
 C6 08 C2 5F 1B 7B 3C 84 2B CB CA 61 80 CD 6C 8C
 F7 69 C5 6D 05 5C 41 4C AA C8 B9 E5 C7 FD 39 47
 E9 D4 4A 58 A8 59 F8 AF 5F 32 35 07 A0 BE EE 31
 1F 3E DD B8 F4 3A C9 9B 53 66 C0 BD 89 33 B2 98
 3F 48 CC 03 F5 67 A0 01 2D 4D 3E 41 2B 33 91 20
 9E 62 A2 16 99 D9 6E 42 66 04 F8 9D CE 57 D3 53
 BF 11 D9 E9 4C C7 F0 EA C3 44 F8 13 83 D1 4A 51
 3A 71 8A F9 AA E8 B5 13 59 41 D7 C5 DE 59 3C 22
 05 1B BF 92 0D 1B F4 42 70 63 F8 3D DA 4B 54 42
 0F A3 9D 81 E8 AB 51 3B 0A A7 60 11 8C 2E 3A A5
 E0 48 1A 7B 2C 7D F9 72 18 7F E2 13 CE 3E 7F 1A
 3F A2 72 C3 D2 A0 DA 3F FB 3D BB 02 CF EE 6A C1
 1B 72 F2 10 05 C6 3A 96 31 07 36 E8 DE A3 8D EE
 40 6E 3C 38 B2 FA 41 44 D9 2B EB 36 33 D9 08 2B
 0A B6 DB 37 EF 71 49 36 FB 05 8E 3D A5 89 A2 41
 C3 31 4D 94 3D 8F BB 84 22 64 E3 66 AD 21 34 B7
 63 CA 04 22 5C 6C 6A 57 AC 2D BF A9 ED 5D 52 B0
 22 8F C9 0F 5E 6D 61 1B FC 49 0E A9 92 BF 24 76
 B9 82 D2 FD AA 10 3C C3 01 57 3A 02 A2 8C 03 7B
 5C E5 87 CE 1F 51 CB A4 17 E9 9D CA F5 48 80 EB
 4C 4E 4E E8 C5 26 42 CE 57 B9 AE EC A5 AD 80 EC
 C9 C4 08 E9 83 D2 2F FD B8 24 A7 0C A4 8A B6 FB
 1B AF 8A CB F5 81 98 17 AD 30 4F FA 48 02 E6 2C
 4E 46 64 7C 20 02 9C 41 87 A7 9D 2D 85 22 14 73
 A3 5D 22 99 08 3E CE 7B 54 1A C0 1C 0D 43 73 F0
 04 A1 9D 07 FE B7 9D F3 46 45 55 E0 00 35 76 3A
 F5 B8 23 C5 27 37 CE 0A 4B 6E FF 61 9D A1 23 95
 B1 63 FB 6D BE 01 9D B1 66 B7 36 62 BB DE 70 D1
 8D F3 3B 64 76 FC 41 B6 59 5C FB 09 C3 36 2C B2
 E8 F7 23 3E A0 B3 23 A1 C4 E7 1D B7 11 54 8D EA
 AD 23 71 5B 3F A4 EA 77 68 42 D8 61 8F AD 93 8D
 C2 09 52 26 FB 44 88 93 41 36 FA AC FE F1 35 46
 9A 23 14 C4 4C 3A F9 34 3B B8 63 8C 01 F0 D7 EB
 5A B0 DB 96 F2 75 87 F9 28 FE C2 52 58 62 94 54
 16 2D 63 44 48 CB A2 F8 03 0B C8 44 6C 45 24 6F
 ED 42 2E 62 1D 3A E8 68 54 B7 F5 29 74 C7 BF CA
 EE CC BA 68 B4 19 71 9E 79 A5 26 3F C4 0E 08 BA
 0D 90 70 E4 A6 4A E7 21 6D 18 49 0A B2 AF 55 3D
 B4 AD C0 1C 05 AB 29 79 90 84 E8 FC C3 ED 10 DA
 B9 4D 80 E5 27 10 4B FB 26 C8 1F 8B 2F 44 C8 E8
 E0 68 FC FC A7 AE F1 ED 37 F9 07 E1 05 FE 4A FF
 E8 E9 30 0F 60 9D B3 E6 FF 28 86 1B 88 14 F9 53
 8E 3A 9B 2B D3 0B BA 97 51 0D BA 18 53 D9 E7 44
 3A 92 35 C7 12 CD FC FF 06 31 37 3D 9F 44 D4 ED
 5F 24 3E F9 6F 1C B1 5F 32 35 F0 E2 AF 8F C1 28
 13 D1 6B 62 CB 08 DF 00 F4 27 DC 7B 06 7C 10 CF
 11 E8 8D F0 78 DD 02 74 30 C8 E5 E6 32 43 F2 4B
 A6 88 E3 91 71 C2 6F 8C 41 C8 62 46 B6 43 B4 9A
 D1 22 63 64 92 65 E8 2F 47 59 27 4A B1 FC B8 6F
 94 81 5B 3C 06 20 1C 3D 44 A0 C1 0C CA CA FC 10
 65 AB F9 85 FE 27 12 4B DE 7E 2C 42 37 D0 FC 7F
 DB 32 39 0F 14 EC 43 9A 6A 9C 3B 38 01 40 AC F9
 5C DE 34 DD 2E 9C A6 90 27 26 1F 13 53 92 DB 16
 96 4C AD 7B F0 34 9F 8D C0 5B A9 7C EE 94 0C 3B
 B2 A6 F9 27 4A 92 32 00 16 2A 14 41 7B D8 86 D2
 64 06 7C 49 E3 A4 85 C9 A2 70 6D F2 F7 90 F2 86
 B6 AB 2F 63 A2 99 1B 04 FD 48 72 1A D3 22 0D CD
 2A 41 BD 5B 68 34 F4 14 E0 57 DB 15 3A 17 15 18
 5D A5 3D 33 C5 B8 9C F6 30 73 89 E7 C6 D5 59 FF
 17 04 DE 2E 33 8E 5C 39 0C 90 07 43 6F 20 F2 FB
 9E 52 92 5C 00 3E 15 DF 86 A4 B8 81 00 10 FF 65
 85 4C E3 B7 FE 1D 61 51 83 3C 24 F3 02 F4 B4 D0
 9C 56 91 7C 8F 86 0F D9 BE E5 35 39 C8 20 A7 1F
 B4 27 D4 0B 8A D5 09 8D 35 4B B5 1A 62 B0 D6 0D
 F2 97 93 82 1F F8 D7 80 4E DA 2D 40 32 D4 E8 E7
 7E A9 C2 6E 2A BB 5A 4A DE CB D8 B6 FC 01 EC 6B
 3A BB 54 7D AA CE 63 A0 AC 2F CE 6D ED 3D A3 31
 5A CF C5 BD 1C 94 C7 D9 F4 85 56 66 56 00 12 A1
 C4 FF 49 D7 B6 BF F4 3C 7A 11 2B 5A 9E D1 90 90
 0F D8 B9 4C 7E 04 EE 0E D7 41 DA 0E 01 8B 61 AB
 13 4A 10 F7 C4 D8 98 CF 42 D2 03 87 5F 7C B5 38
 0A FD 8B 37 6A C1 56 CE B6 45 F2 00 20 52 0B 36
 26 7B 96 D7 7B FD 3D 22 C2 4E 49 4E AD 6C 09 8E
 D8 9C B7 6C 23 AE 05 71 35 18 09 A8 AA 9F 6F 11
 C6 12 D0 71 4A AE 95 5F 6C CD 78 C7 25 F5 AC 41
 F5 9B 2E 27 66 45 A0 3D A0 E3 4A 43 D4 36 81 25
 48 C7 C2 64 9B A3 E2 27 35 73 91 EB E8 9C A5 4F
 B6 51 A8 4E 55 FA F8 0C 93 C2 34 CF 46 49 C2 77
 26 11 0F 4A 22 10 D7 AB 9B 55 B5 B9 DB 63 38 A9
 C1 3C 76 0A CF 30 3E A3 83 74 E8 58 E7 DA FF 92
 2D F7 B4 31 26 B8 26 96 AB 52 EC C3 92 66 1B 71
 B8 87 26 8F 84 3B D4 EA 9B A9 79 04 46 B5 40 98
 A8 FB 9F F5 1E 2D 2B FB 00 C9 1C 1B E8 4A FF 41
 2A 90 F8 49 58 63 04 45 41 26 B0 83 44 68 5E 48
 98 FA 4C 19 FE C6 D3 5B E3 48 A1 D9 6E BA A6 36
 77 53 22 C7 98 F4 4D 0B 1C B7 AD 6A 78 2B 89 86
 B5 24 80 69 97 DE 8B AD D5 27 AC 49 05 0E B8 76
 10 F8 9C 5C 61 D7 F4 BB F8 34 BE 10 4C FB 9C 6D
 0A 05 EB AD 0E 85 E4 05 AC EF E8 12 14 54 56 E3
 98 CE 5C 63 D1 4F A0 C7 F2 95 F5 91 04 39 34 FE
 54 62 C0 16 D2 AD 47 43 22 54 19 1A 89 F7 75 63
 E8 C2 78 42 AC 4E 8C BD 8B 58 B4 1D BF 01 DC 66
 4C 3E D7 E7 3E A5 A3 11 27 BE CF 8B 59 4A CC 6F
 D7 7A B9 04 F8 7E 66 5A 90 FA 28 8E CD 64 E2 09
 AE 88 D9 C3 19 13 52 69 1B 21 36 B5 8E 6A F3 CC
 0D 0C AF 4C 6C 74 12 FB 27 D7 81 7F 2B A4 28 45
 79 1E 08 75 37 10 2C 1D 27 2E A4 7C B3 7F 04 4B
 E3 39 20 D6 75 85 98 C0 73 DF 1A BE B7 6F 31 4F
 EC 84 86 11 59 9F 11 C2 E2 DC AF 2C E2 E1 7A 3C
 30 7F 1A 17 4A EF 57 51 FB 38 BD E2 00 36 BC 82
 8D 36 73 E5 5E E9 94 6D 9B 8F 93 35 C7 F2 80 B1
 32 E9 AE 0C F9 E8 FC 3A 2F 24 90 D1 CC DC BD 40
 0A 71 85 2C F2 47 25 CE 6E 2D AC DC 37 DC 03 B9
 94 CD FD 57 CB 99 F0 4B F8 38 21 50 9A 04 81 9F
 24 B6 12 CE 2E D8 44 FE AF 38 A8 97 03 26 66 85
 72 F6 A5 72 76 45 7A 7B CF 4D CA 6F 01 0F E3 BA
 9D 70 70 AE 17 F7 DD A2 6B DA D2 55 BA B2 99 98
 FD DA F9 33 CF F2 BF 55 91 4D E5 D3 11 FE C8 6F
 E7 CD 38 F8 A6 27 DC CF 03 44 32 F3 84 E9 8F 0C
 57 8E F2 40 1D 94 38 E6 35 0F E1 96 77 34 37 1E
 29 BF 62 17 89 54 33 81 1C 53 05 C0 5F C9 18 37
 86 2F EE 63 C3 F6 39 EC 8F 86 82 50 B1 CC 3D F1
 D0 D8 A8 1C D0 16 6A 67 F2 FB 7B 46 F7 6F D1 A0
 98 83 DA A7 0F 9D DC 89 99 17 A9 B8 83 E3 E3 AE
 39 9D 94 84 11 A9 E1 2B B6 91 41 AB 56 4A 3F BC
 08 1B 8D 3C 68 A6 7E 7C 9C 86 44 32 57 92 81 62
 9B A2 39 9D 12 BC BA F8 EB 24 AF DC 44 22 39 6F
 33 7F 30 36 22 73 28 25 3C 5D FD 59 1E 3A 9D 78
 5E 3E 0B 0A BE F8 E8 9C DE 69 5E A0 82 29 55 C6
 AA 15 02 6F 78 C3 92 B0 6C 17 F5 77 45 00 65 FF
 8B 2E BA 2A 51 50 C4 44 59 05 B4 26 80 EA E2 57
 81 C9 47 D2 57 A8 3D CB 2E 9F 8D 52 AA 2A 92 B5
 06 B0 D0 C2 4B FD 55 11 1A 07 FB 72 E7 74 63 2A
 99 3A 2C E2 56 EE 87 78 AE 5F 9C 01 C3 A7 E7 50
 EC EE EF CC BF 0E 4C 69 FB EB D9 3C 84 F4 C7 3E
 9D 1C BA 25 FE E7 EE 24 87 75 5D 79 53 36 AD 09
 4C 28 7A C9 2F 28 48 28 D8 1F B5 76 80 11 7D A1
 2E 1E 02 35 21 8E 49 25 E3 54 11 17 D0 CF A5 29
 53 4D 21 7E B3 13 54 42 D3 6C 99 B6 1E AD 44 D2
 37 82 62 45 BC A0 E6 75 AC B5 93 A9 46 CD 37 60
 5E D2 58 F2 93 38 BA A7 47 8A F3 F0 D0 00 EF 8B
 15 FC 6C 31 67 DA B1 F7 B9 ED 31 40 46 3B 90 32
 CD 15 A7 C5 A4 CF F2 51 91 75 16 85 D7 D1 08 5C
 EC 80 1C 74 DE 42 80 78 95 4B 3C A1 83 95 D7 C0
 23 2E 5D 7E 46 A8 ED C4 52 0A B0 A0 15 F9 49 C5
 DA 42 B4 4F 97 5B B1 E8 BE B9 19 B8 D9 50 8E C5
 E0 A0 0E 6A CA 07 F0 72 55 DA DB 15 C0 F5 81 DA
 3E 10 89 2A 7C 71 45 52 47 BA 42 F6 4C 05 F1 F5
 09 18 91 85 43 85 EE DA 3D 6B 11 8D FD 59 05 6D
 4E D2 A0 53 8F B8 AD 35 26 05 3D 83 DF 5B E5 A8
 90 83 DD D3 AE 66 68 97 61 57 AA 13 9C FE 31 3F
 60 54 18 D0 89 F2 3F 6B 3C E7 FC 16 63 18 31 4C
 F1 CE 97 12 AE 07 6F 49 4D 97 53 3F 77 7F 8E 03
 BF FF 1B 09 B6 DC 4B 3D 85 BA DA EF 60 61 BE A7
 1B 00 AE 6A 6D 05 AB 8F F5 4F FC 03 3F CA 08 92
 A7 3D CE 19 2B 33 2F 75 0F C8 72 E8 40 44 9E 61
 F4 6E 0D 8E 19 EE 36 51 27 30 11 F9 B0 5F 10 1F
 77 42 50 35 EC 83 16 D8 C3 63 C8 43 55 C5 B1 2D
 89 53 04 3B 74 88 A3 F5 B3 D1 3B E7 07 71 24 FA
 18 13 22 F0 92 29 47 AC A3 35 7C 66 79 F2 C7 8E
 11 D5 DE 11 4D 49 35 0C C7 4A 0B A0 CD B7 DF 20
 B1 52 76 64 5B F6 1C 42 29 8B D8 00 F6 8C B2 B2
 92 4A 37 37 59 97 BD 2F A4 47 79 DA DB 1D 02 F7
 F9 A0 78 3C 32 17 34 0F 49 6D 99 F8 EA 26 B1 78
 B5 60 3E E6 51 B1 85 AF BB 57 39 4A 4B AA CC 5A
 2F 82 B2 F2 95 F7 9D CD 18 8B 8C 7C F7 DF ED 81
 46 22 1F 44 2F 7A 32 AE C0 20 03 2C EA C2 F3 0C
 41 F3 6A A5 91 79 32 06 75 BC EE 7C 32 01 4C 26
 BC 29 D0 ED AF A5 2A 1F 3E C6 6D 0D 02 97 52 11
 36 5F AA 48 75 5F EE CB 0D F1 22 18 8D 21 D0 9B
 EB 2B A2 A9 9E 2A CA EB EC 15 2A 29 B0 C2 AB 0C
 D3 DA 8C F4 7D E3 65 A0 F1 0E E6 F5 E0 D3 6F 21
 52 24 F3 44 32 1E 71 59 66 FA 1B 90 E1 F6 D4 85
 D9 BD D5 DC 55 0F 6F 9F D9 FB D6 C6 CC 41 CE 7F
 9C EB B2 39 8A 82 99 AE F4 DD 79 D4 C5 15 89 1F
 2D 64 97 73 AD E7 A1 0A 56 D7 CD 01 E5 62 31 57
 8E 6D 4E 56 6A 05 B7 9C 3A 7E 32 8A AE FD 67 7F
 69 50 EB FB F7 35 E2 01 E6 42 D6 FF 37 E6 8A 9B
 E4 B4 B5 39 26 44 C0 B8 4D 59 C8 AA 63 25 1A 1F
 25 03 93 B8 5C 38 01 21 BF 91 FC AC BD A4 F2 54
 DB 01 D7 0E 0E BE 5F 27 EE A7 0D F7 0A 11 69 9D
 5E 45 93 FD 8D 1C 2F D7 F1 69 1F BE 82 DE 1A 3A
 0C 69 4A 60 46 0E 95 1B B5 13 09 83 C3 93 25 61
 F8 C6 F8 9D 2D 32 92 17 50 EC D9 27 00 61 3E 60
 20 73 8A 81 B9 2A 6D 25 13 5A 07 C8 17 21 6A 6D
 0A 74 2B 5F 76 A4 AF 9F BD 9C B7 46 9C D5 7A C9
 57 25 01 81 BE 06 35 A8 CA 92 8C F3 BB 7D 49 7C
 BC 64 7E 7B 82 9B B9 E5 A2 1B 04 03 BF 7B D1 F4
 63 9F BF DB 60 6F 58 F7 1E FB F7 DC 83 A2 BC 8A
 74 0E 02 92 CE 49 ED A5 D6 6D 70 27 4E 94 49 B1
 CC 78 B1 52 14 8B 47 13 7F 73 27 E4 D7 2F C5 E0
 6A 8E 9D 86 68 20 32 09 C0 2E 81 8D 93 DF 10 60
 A8 E3 79 87 CC 7B 73 AC 2D D2 1A 80 89 8F AE 70
 34 5C 59 88 09 E6 D0 E6 8B E1 68 57 E8 AB 7F 80
 14 6F BE 0B 2F 74 0F E6 18 30 88 7C 8F B9 48 5F
 DE B5 EA 8E 7F 82 13 41 CF C0 7D 9E 4C 46 D6 EC
 E5 43 22 ED 60 7D 6C 64 24 17 62 D2 90 07 01 08
 BC 87 30 55 0F 58 76 A5 97 92 F6 EB 96 63 2E 26
 01 82 B6 48 C4 B0 DF EB DA A4 D3 D4 9E 8D A8 CD
 CC B0 2D C8 6D F5 4B E4 D9 22 67 79 4E DE C7 82
 E3 1E 13 37 C3 73 56 EF 86 F1 8E 3E B9 B0 C4 CC
 1A 47 37 B3 A3 F7 0B 6D 6C 3C 7E 62 59 6C 5B 3C
 9C 42 C5 C5 7A A2 F3 C7 11 1A 14 18 8E 04 FF C4
 74 7D 12 16 16 46 D6 DE 27 66 BD 13 90 04 97 6B
 42 D1 9E A5 39 66 AD F6 A2 7A 54 B9 CD 78 34 39
 5B 7F 63 BD 22 72 55 C2 5C 24 A5 86 F5 39 AE E0
 D4 95 E6 0F EC 29 0F D9 97 3B F2 DC B1 AC 89 7A
 66 4A BA A8 B5 E5 24 22 EF 20 3A 6F 8B DC E1 94
 5E A4 1F 31 3B 98 A4 09 97 C7 E2 B6 65 11 FB B5
 2C 37 B8 9C 0F D1 78 82 02 0A 36 5A 34 EA 86 3A
 8C 1C E1 24 95 5D D5 10 63 B7 00 67 7E 0A D6 2E
 DB A2 4D F5 94 52 67 30 D1 54 63 D2 B3 5A 64 29
 3A 7B 56 01 CA 22 73 D8 F9 C1 D2 C0 8C A6 3D 10
 1E C8 EE F2 16 3B 3F 10 1E 76 AA 34 7E B6 E3 81
 A8 32 73 CB E0 04 34 39 A7 43 BC 3D 52 2D 18 B7
 BA 6D 89 CE 8E 81 65 64 EC E7 5B C1 24 61 1D 36
 4A C8 50 43 77 C7 C5 03 E0 71 B2 91 B5 FC D7 56
 07 D5 9F 9C C0 A5 3E 98 7E F0 0E 7E 5D 13 3E 0B
 B7 EE 30 3A 2B 52 49 C8 BA FD 38 7B 4A 74 75 86
 1E 1B 4B 78 D5 20 0D 69 FB 24 DA B7 3C 6B B8 C1
 5A E1 F6 D0 AA 02 47 E5 C3 8A F6 BC D3 63 15 3D
 F3 23 2D A1 76 73 88 F0 63 E3 88 95 D6 39 98 9A
 F6 06 63 C3 72 DD FE 8D C0 42 93 08 7C 7D 5D F3
 DF 36 6B 9C DF E0 F3 8F 0B D9 80 51 F6 BE D2 6B
 A0 5F 44 78 C6 80 72 81 48 53 51 43 10 06 86 4F
 EC 14 EC C8 E5 84 4F FA 31 CC 92 14 93 F0 B2 03
 C3 7D BF 5E C4 43 B0 0D 8A 5D 41 16 C5 08 30 51
 A4 4C DA 71 52 02 08 72 E1 4F 7D 29 F8 0C 53 DC
 4E C8 37 F3 E6 C8 2A 5B 0C 88 56 9B FE 06 9F 08
 49 97 13 A9 81 D8 6F F5 56 71 40 9A 5E C8 B3 AB
 E0 76 7C CB 63 5E 5D CA F7 25 BF C9 ED A3 18 67
 61 C5 B7 7F 89 AE 71 DF 37 A1 CF 49 E5 36 3E 1F
 C8 E9 B9 18 2B 92 17 18 58 B0 7C EF 4D 5F 2B 7E
 3F 6A 31 6F 23 9C B1 80 72 7D 36 FF 69 6C A1 FE
 35 D5 25 D6 23 3F 70 5B AD 2C 6C 05 8B 11 1E 85
 0C F6 B6 6C 44 C3 C8 00 A1 85 A6 5E F1 A4 9D FF
 E6 8F 89 1E 60 36 A0 0C B7 AD 4F 3D 4C B0 7E 96
 D9 06 9D A2 BA 0F 2A EA B5 3F 09 B9 38 C5 A7 28
 4E 88 26 8C 3F 1A 47 B5 EB 8D 50 6A 54 2E CC 26
 D7 3D 3D FC 71 CD 84 51 97 16 E9 C4 DD C7 47 FF
 6D 3F 92 A5 41 57 53 BA 1C 15 C0 47 48 E1 D2 7D
 59 40 E8 AF 5E 77 12 71 AF 4B C5 0C 9D 46 D5 63
 E0 1F F4 57 C4 D6 48 B8 8C C5 9C F8 52 B3 12 4A
 44 C4 9D 11 73 36 B3 4E 0C DE 21 06 6F 5D F5 BE
 BD E1 EB B6 E8 91 94 6B D3 6F 3A 2A 84 5C CD 03
 C8 BC B5 3D 9D 9B E2 EB B9 F5 6B 62 B8 78 2F 43
 A3 50 3C F4 F7 21 36 C5 BC 23 50 E4 70 11 82 1C
 DB D7 D6 32 E0 9A C6 28 E8 19 96 1B C8 17 46 DD
 91 2C 2D 7D 2E 85 B9 69 4A 53 0F 44 85 FC 5F 75
 70 AA EA DD F3 22 E9 40 43 C8 2B 7C 45 65 B1 76
 1C F4 FF 3F 16 E4 D1 9A F4 32 92 F0 8F 6F 50 CC
 FA D1 F4 94 A1 5D 2E 26 22 24 DA 92 92 67 20 5E
 FC CD DE 9D 45 EA B6 B1 37 11 3B ED 87 A3 8D D0
 62 8F 0D 46 A3 9A B5 2D 5F E9 1C DA CC 58 D3 68
 3F EE B9 6D 24 EE C8 04 51 19 3A 8D C1 C2 F0 FD
 63 AF C7 FD 04 76 38 75 62 DD FD 0C 85 9B 51 EB
 AB 69 30 74 C3 27 EA C2 68 7B F3 DE 05 DB EE 9D
 D9 62 D3 2D 5D E2 DC 02 65 8B 97 DE A7 9E B6 A0
 F4 67 BA C9 E9 45 6D 3F 5C A4 47 E3 28 7F 3D D4
 70 3A E6 79 FE EF 89 E9 43 64 EF 04 25 FB 1B 77
 14 6A 76 61 A2 2A 54 98 52 B4 90 60 E5 9C 6C 04
 57 CF AD 23 25 69 A9 A9 53 87 67 FC BD 53 5A C0
 82 50 D1 4F 6A 42 F3 BC 82 84 54 B2 18 BA 3F DA
 B8 5E 42 17 58 81 DA C0 9B 46 19 40 CC 4F 6D AD
 8B BD 02 A6 40 7C 08 1D 3D E5 94 57 D9 69 F2 C7
 B7 21 6A D7 E0 05 66 22 23 28 B5 34 C8 08 19 18
 47 42 59 B5 8C E6 0D A1 AD CF 2E 3E 5F 2C AA 6E
 1A 98 48 C8 AE 92 EF F0 6A E4 B0 F7 85 09 5D 08
 FD 80 A4 E5 27 D4 2E 6B 0B BD 0E 72 8E 05 DB 0F
 A1 E3 36 9F 1A 0B 63 F2 4E F3 49 A7 4E 39 B3 57
 49 76 F0 57 10 16 DE 5F 63 AA DA B9 37 A0 49 7F
 BB 79 EE 0F F7 DF 6B E9 C4 84 D0 32 E8 8C 09 BF
 2A 1B AC 36 46 5F 11 42 0F DD AF D2 63 A3 78 C4
 AE E7 9A 46 86 2E 2A 00 F5 2D 24 9B 65 51 B2 91
 BD 61 3E 31 ED A1 85 AC 71 CC 83 49 DA 11 8E 56
 FA 92 68 AC 5D A4 D9 1C 1F B1 FF 7C 2D 93 A0 AF
 AF 53 F6 61 CB C2 27 DA 15 0C AC 43 13 D5 6E A3
 ED CE 88 4E 98 73 65 18 B4 CE F4 D6 19 C5 49 D7
 94 CF CE B5 85 49 5A 2D 98 02 C3 9B 57 24 CF 7B
 87 33 F7 F3 C6 5A C4 08 DE 34 76 18 A4 2A 40 E7
 C5 3A 6D 10 54 B3 80 55 C0 85 92 A8 CC BF 4F DB
 50 9B A4 22 D6 65 91 0E 9D DF 63 04 1A 67 C3 A9
 A0 E3 59 48 FE 2B D7 92 C5 6F 7A 45 D9 E4 53 92
 A3 17 B8 D4 D1 62 97 E2 E6 A3 7A 87 76 3E 61 36
 4D D3 BC E2 CE 44 41 85 AC C5 D4 87 DE B0 C2 63
 98 60 6F 8C E3 90 3A 1D A6 A8 E1 B4 7E 77 58 D2
 96 E4 F4 82 1D A7 7C 16 EF 3A C0 40 A6 D9 B7 90
 DA 37 0A 7E ED C1 89 3D DD 5A 08 F6 9A 15 72 53
 25 36 98 4D A4 62 B7 3F 00 33 B0 59 4E C6 1A B8
 B7 67 19 32 A0 3A 8C 26 DE CD 51 3C 1B 7F 59 F1
 84 28 1F CE AC CB ED 17 40 A3 EA C4 12 7C 03 87
 5C 0C 58 FC 0C D3 15 B7 32 1F C9 0F EC B1 B0 79
 33 5F F9 7F F4 0E 79 F8 F4 07 B7 7D 80 AE 18 E2
 EA 53 43 AB 23 93 88 CB 8B 5C 93 D6 89 71 60 38
 81 EE 01 CA 1E E1 EC BE 3E BE 21 7A 10 2D BF 21
 68 DF 47 B3 0D 95 90 B4 B8 50 60 E4 08 D8 18 9C
 3C 3E B7 BD 71 21 27 9C CF BC 93 FF 2B 96 AC C3
 CC 56 4D E3 AF 61 1F 57 7B 53 45 F2 5F C6 5F 09
 70 FF 63 B6 3F 46 D7 13 D3 22 92 1C C1 80 7E 9F
 42 FD 24 41 1D 0D 50 63 A8 4C B4 4D 91 EB E7 2B
 C4 32 26 72 07 76 07 8F C7 9B BB CC 93 7A A8 89
 38 60 6E 6C B5 88 49 41 91 23 F7 15 83 A9 7A 3E
 A7 B7 83 75 75 84 D6 25 E1 25 C0 C6 14 A4 BB A0
 B2 F1 37 0A 77 47 94 76 05 87 B7 31 91 B6 8C 5A
 11 C6 6D A1 84 78 0E 95 DB D2 79 3D DF 8D 3E 43
 20 FC 47 36 00 2A 04 55 C6 B3 96 D5 F5 CD C8 96
 FF FF 1A 0E 89 F3 6E 75 24 87 A1 BF 1A 1B DC 49
 52 98 85 CC 27 BB E8 D0 F4 B1 69 9E 7D B3 CB 66
 40 B6 58 30 1A E4 C6 16 86 DA E3 EC D5 77 09 6C
 14 15 31 01 E6 A6 AE E7 8B 46 65 0C C3 CA 16 C3
 E6 B8 F5 C4 D8 15 33 10 AB 5F 44 4A 45 DB E6 23
 75 62 6A 0E 8A E7 06 F7 95 5F 18 81 14 A4 77 2A
 15 7F 01 24 5B 5D 1F 86 A5 FE 4E 0A 62 A0 9B 14
 3C 22 FF 5E AD 88 2E 68 C3 4B A1 26 CC C5 F4 56
 6E 19 0D 72 0D DE 91 3F D0 2A EB A9 D3 2A 52 E9
 56 23 1C 51 72 9E 51 D8 3F E6 CD 91 63 F4 59 84
 C8 F0 53 9D 74 90 06 1A 04 42 49 46 80 AF 90 C9
 DE 0C CD 42 83 46 B6 64 EC 01 68 A4 C4 B2 03 43
 EF D4 69 CB 29 85 C8 15 F7 DA B5 F1 AD D6 53 E2
 23 38 3F 85 4E F1 1C FD C1 3B 25 ED D2 46 9E 42
 1E 4E 0A 46 33 68 20 62 03 45 88 73 35 EA 22 A5
 97 97 2F 7C AC 90 B7 2D F8 0F 60 26 23 69 50 A0
 ED 2B 46 03 CA 37 BE 8C 1E 5F B0 D8 23 73 FF DE
 FB 01 49 EA 31 04 57 ED 54 F9 53 8F CA 10 AA AD
 70 F9 4B B4 5D 2A 45 A9 F3 1F 74 79 B8 26 85 D1
 97 96 C5 54 E3 AF 02 B0 73 0E 4C F4 8D 64 E9 D1
 C1 C6 DB 86 39 DF 5A 48 BB 4D D0 03 37 FC DF 47
 45 E0 E8 9D 44 41 C0 72 11 EA DE 21 7E 27 E4 F4
 51 15 B3 67 52 13 6E 36 AD D5 F1 DE D9 6D 40 03
 4E 0D 75 22 7A FA C0 5C 3E 1C EF 79 DE D7 C6 85
 B2 EC AD D8 5E 37 42 91 3B D5 AE D1 2E C6 5A 7F
 4B 4B AF EF 22 E2 4D 51 FC C5 A6 24 06 17 34 21
 0C 62 C7 F2 D1 9B FE 45 0C FE E1 50 38 A0 88 DE
 85 4F 5C 22 18 B1 C1 C3 EA E7 EF 49 16 83 64 65
 BC 45 9E 64 22 24 A3 49 7B EC 5A D3 4D 5C 27 8B
 7A F2 19 D3 81 5F 4A 18 2E 93 4B E7 1B B1 BC 99
 0A 0D E9 F0 00 FF FC FE DA 9A 72 E9 3A 1A BA 3E
 63 AE 71 3E 28 02 5E D5 05 E0 0A 19 36 F9 AE 9F
 98 46 0E 75 AA 75 ED 0F CA CE 60 CC B7 27 20 F7
 B6 9F 8A B6 51 5E C6 9B 3A 40 03 87 F0 E9 F0 78
 23 DC 9F 90 48 D7 41 72 D9 DC 9B 5B DA E3 46 6A
 A8 95 A7 0F C5 27 71 4F AD A2 66 4C F9 55 55 AD
 FC 69 07 DD 39 86 83 0C 74 D5 3E B4 73 4F F3 FB
 85 48 14 6A 6A 9C 7D 60 42 A0 08 70 32 03 0D 7B
 CD D6 B6 24 95 71 A2 B6 F2 E7 33 BE FC 98 C6 E8
 E9 88 9C 8C C4 11 AD 1B 29 C6 86 12 E4 55 9D 3C
 80 72 A8 02 98 92 3A 10 A0 B0 A9 C0 04 25 EB CC
 F3 CE E9 CB FD F6 20 F3 E7 07 61 AE 15 FC A1 E0
 70 BD 79 2F 3D 91 99 4B DD 7D 6B 03 16 EE 51 67
 8A 6C F9 42 1C BB 0C DC 3D 62 A1 AE 85 63 5F 30
 B6 EF 81 C8 AC BA 70 1E 26 AF 59 CB 14 70 E1 C8
 1B C6 F9 C2 FA 6F 91 B5 4E 32 F6 C3 3A A0 B5 6F
 87 21 26 73 C2 78 5D E4 E7 2B 74 1E D4 83 2D E5
 32 86 3D 0B 18 34 20 31 93 97 25 05 61 9F BA 69
 72 D7 36 23 31 F4 99 C9 0C 4A 4C 18 97 77 D9 C7
 1E 38 F3 9A B2 2C D8 2F ED CB 6A 8E BA DB BE F8
 9D 3B 4E 1A 99 08 F6 E6 9E 4A F0 D4 87 60 4C 67
 22 44 64 79 D9 EE 1D 71 21 D9 90 94 48 31 9C DD
 B2 56 66 78 B3 C5 BD 50 8B 5A D5 B3 3B 83 9E E2
 72 B5 16 3A 96 09 0A 1F 87 CD B1 97 54 C5 DF EB
 19 71 EA E7 26 E5 03 FE ED 5C F8 54 5F 89 27 EF
 CC 70 C0 00 D2 6A 43 C5 5E D6 59 1B 16 B8 91 2B
 ED 20 7B 6A 61 17 42 56 F1 AB D7 5B CD BF 61 0C
 03 54 F1 C5 8F 64 7C A5 4C C4 64 45 C4 3C AA E4
 68 97 73 1B C2 F7 46 72 E1 16 61 9B CA EC 85 25
 53 EF 4D 90 54 B9 82 30 ED 67 EB 71 E2 C9 AA B9
 DD 26 70 B2 D0 4D B1 C7 4D 9C FD 50 AA 17 A5 91
 7F 27 E0 53 5C 24 A4 AC C6 04 3F C9 68 4A B7 6B
 FA 61 98 D8 CC 88 6A 9E B6 95 05 2E E3 B6 0C 8E
 95 26 A3 5C 6A 36 39 98 DE 6F 96 9F BF 43 74 27
 A3 6C 2E 0B 79 1D 99 49 E0 27 81 B4 C4 1E 36 0C
 80 83 63 DB CD C5 ED A8 8F C0 DB F5 26 A4 74 E8
 EA D9 F3 82 BF C0 AA 9B 9B 06 A3 BA 0A EE B3 09
 2A F3 9B 07 B6 C5 DB A1 82 D0 36 DC 8D 08 3A A6
 FF E4 FB 9D BC 82 78 7E E4 BF 76 8F 70 E9 4F 61
 C7 72 71 5F 23 4C D8 86 20 EE 58 4A D8 54 C9 11
 EE 0C D9 D1 16 AD 01 F2 CF 5B 4F EC 62 B5 4F 1C
 95 82 76 C0 FB 25 EF F7 B9 4F E0 F0 47 33 A5 98
 68 93 4C 72 DC EF 9B 9C C6 9C 9B 26 AB F1 41 06
 15 B7 2D FA 18 0D 29 5F 6E C4 31 A4 D9 70 DC D2
 0F 60 C3 11 08 D1 C2 36 B3 15 93 D0 CF CA E1 9C
 EF 17 BF 8C 13 FA 46 99 58 14 0E 7A 84 93 A6 57
 60 1E 4E 7A 93 61 EB 72 8B 68 10 A2 77 7C A9 A5
 ED 2C 91 C1 70 33 4B F0 0A 4B 6B FE 1B 7A 17 0B
 0D F0 8A 97 8E 33 39 33 D3 99 16 05 09 13 FF AD
 D2 83 8B D5 C9 15 B7 F4 71 DA 22 7F BB 16 0D 32
 BF 51 A5 A0 60 BB 3A 57 9C 42 DC 2C 8D 33 75 6D
 FC 17 96 54 9F 76 CE 07 36 A3 2F AE 2D 46 37 27
 D8 C3 74 75 8A 19 1F 00 FD 39 09 E1 6C F8 D7 03
 C3 D9 3F 49 6F 80 EB 43 D7 A6 9C CE 05 22 6C 3C
 3E 90 A6 E9 87 A9 E6 CC C3 1E 6D 14 7F FB 1D EF
 DE 1B 49 B0 58 B5 69 9A 98 FE EA 5A 35 55 A3 59
 C5 70 17 44 8D CE 7B B1 EE 35 C4 6C 85 BF 3D 60
 E0 7E 57 42 BF E9 D2 AA 3F 9E 4B 64 C3 16 12 DB
 F6 33 FA B4 3A 07 9E DF C3 E6 46 06 AA 25 73 D3
 B0 E3 03 E4 42 2F 61 A3 A9 26 6A 27 BF 50 31 F0
 C3 6F 10 DE 00 B0 50 BD 51 D9 2B 84 CF 35 20 4A
 F6 79 A2 13 86 56 99 A7 B9 B2 91 90 A4 C4 DC F8
 51 AD 55 07 4A 0E 69 7F 15 9D FE 81 75 7C B8 1E
 9C 4A 1D A0 92 32 AD E9 95 E8 00 E4 C2 A1 7C 7C
 28 80 DA 3E CD CC 73 43 AC 93 D5 88 F9 27 C1 D9
 A6 97 B3 31 4E 8F F4 08 0A 17 10 E4 04 A4 89 48
 B8 48 68 B9 AC 70 B7 52 EA 11 AD 55 2A CF 0D FF
 B0 86 B0 D4 71 86 D0 A1 F5 81 85 A1 53 9B 83 96
 C3 8A 20 24 2C 30 8C DF 40 E1 FD 22 BE 13 35 6D
 7E F4 49 65 CB EA 54 1F 7C 3C CB 57 E3 B5 DE D2
 45 EA C4 C2 A6 59 36 BE E9 D7 A5 20 F4 FE EC 19
 48 A7 F4 D9 75 48 59 65 CA A8 CA 97 25 82 D3 02
 B3 C9 04 BA BE F9 53 95 C4 14 2E 60 22 11 C8 0E
 BF 30 1A 1D 4E 01 4F FD 26 25 B4 F2 CA BA 77 94
 F1 DE CB 60 2D 06 2C 7B D3 36 18 C9 3C 01 02 45
 D7 9F 8C DC 65 6E 99 59 4A 72 D9 26 61 2D 6D 23
 E3 3A C9 89 4F C0 23 7B B1 BE 82 44 4C 73 49 9B
 16 16 88 C4 FB 93 78 FF CC 7B 9B 7B C4 A3 0B 96
 39 3D 69 77 1F 5F D1 83 FF D1 D8 34 F3 6C C2 C1
 54 5C 08 67 D4 C0 0F 1C 63 88 E5 B6 06 E8 6A 50
 3E B0 46 1D B0 29 65 6E 73 06 B9 E9 44 7E E6 B9
 E3 2F F8 49 EB 3E B4 A8 71 09 FB FB 59 ED CC 7C
 F0 8E 66 E7 7F 60 8A C3 F9 2E DD C2 7D 10 FB 19
 EC 04 2D D3 91 EE E9 6D 73 AB 28 00 95 15 FC 00
 59 B0 36 C9 10 98 9E 44 9E 84 6B 5C 4A 04 2C CB
 17 FF 5F 0C E9 7A 0E 46 DD 7C 68 3B B5 3E 18 45
 E9 02 63 67 BB E9 56 F5 B9 81 45 A9 8D 12 49 7B
 D1 CC 4F 90 CC 82 39 E8 DE 75 0A FB 4D 44 95 C4
 43 DD 6F FF B3 79 B3 6F 7B 0A C0 C6 94 C7 9D 09
 60 56 E3 7C 37 1A B7 31 DD 32 BD F7 45 A9 E8 CB
 7E 37 D0 C2 98 4F 1C A6 EA 01 2D DB 1E 07 5E E1
 37 86 27 EC 91 8E FB 42 AD 63 44 8E 52 02 34 C2
 37 1F 68 7A D2 6E 25 0D 17 93 54 6D 02 21 5C 54
 36 B2 0E 89 CE 69 45 29 C2 B5 02 8E 89 CE 5A A1
 28 2D 65 0B BE F7 03 34 6A 68 E8 9F D7 10 8F 2A
 4D FD 6E B9 28 4D FB F3 E2 F3 93 13 FE 0A E3 A1
 49 AC 53 57 9E 40 ED A0 27 A6 BD E8 A9 64 99 52
 05 85 14 36 79 30 27 3F DB D5 03 38 75 B4 3A F8
 54 CC 4B 04 4A AB C2 44 AD 15 AC 25 BE B9 30 5C
 2A 37 39 2F 8C DD 52 BF 4C D1 1F F0 35 29 25 C6
 E0 F6 7F 91 19 45 96 94 73 D4 1C F2 46 9A 38 25
 60 D1 02 FD 9D EF C4 3A ED 81 8A F8 80 DE 35 61
 D3 2D 5B 36 2B D2 1A 0C 56 DD 32 A3 D9 F0 BE 17
 FE 13 7F 84 DD 42 72 B5 A5 75 D9 6B 2C B3 9B F0
 DE BE 3B 78 3C B2 30 20 5F 80 C3 65 29 5C 2E D9
 34 48 BE 1F 2D 8A 57 08 FF CB 38 80 FF 41 FD 81
 F0 2D 3C DE 95 3E B4 FF 88 5F 24 36 6E 15 35 BE
 ED 81 C1 2B 21 53 BA 56 C0 84 E0 3C 90 CF 2C 39
 2C AD 35 68 BD 20 9B D0 7C 4B 0F C3 76 1F BA EC
 59 BB D0 8D 05 DC 29 79 2D 35 E4 DD 75 23 56 61
 51 C2 1D 12 C5 A3 FF 42 23 19 6C B4 0A 09 67 46
 F1 9A B6 17 E7 0D 32 04 49 5A 2B 50 DF DC 14 20
 EA 15 6C EA 79 E4 D6 9B 3B 85 30 0C F2 87 16 FC
 82 FA 99 11 CA B6 67 DE C6 76 7F AF D8 B3 1E FA
 AA 6F 1F BA 38 97 9B 3F 2E 26 CF 4E 4A C5 51 2A
 43 6F 5F 3D 0D 0A 69 E3 A9 E7 3E 63 7E 8A 56 5C
 4A C2 9C 78 CA 9B F8 BE 15 B9 AD 3D FD BD 35 F5
 79 D9 F9 71 FF 51 DC FC 29 F0 08 84 78 4B 9A E8
 94 4E 6F D3 D9 91 35 64 9D 61 7F 77 23 41 11 96
 FB F5 83 94 CE C0 98 80 95 FF E1 DE 4C 52 82 59
 58 D0 F4 29 13 95 8C 0A AE 1E 27 70 26 21 BD D0
 99 B2 A8 3A D9 D9 8C 77 F1 10 A5 CC 22 B9 FC FA
 80 BE FB 30 3B 37 58 18 BD 6D 5E 82 BA 0F 08 B4
 0D 67 5D 43 76 32 28 60 83 B7 59 96 23 A7 A6 22
 27 5C 69 16 02 56 70 F8 46 03 6B C9 13 A4 BF 90
 61 3E 2D 68 50 02 63 66 82 0F EC 0B D0 38 7D 85
 C7 2E 69 A0 BA 05 CA DC 52 FA 7C 1F D7 7D A6 26
 AC D4 FB 6C D0 1A A0 74 6E 46 FC 5F 94 B5 13 D8
 ED 2F 62 C2 CB E5 C2 60 6D DE 84 AF 76 1F D5 54
 76 C9 B0 0F 6D 96 C4 88 B8 F6 1E 0D E0 EB CD 0F
 65 22 A1 41 FB EB FE 95 4F 0D D5 54 12 3C 43 41
 0C 0D 5E AA FD B3 26 10 13 D6 AA E3 32 10 E5 77
 99 A0 95 9A 41 4B 1A A0 05 A4 5D 76 15 A2 F2 91
 DF A1 8A 2C 5B 7F 98 2E 7D 52 01 18 55 DF 3A E6
 A5 59 FB 93 E7 35 76 67 73 69 48 D6 9C CB AA 53
 B1 24 6A 90 FC D0 1A 62 32 1D 7E 3F 7D FB 4E 83
 A3 B2 2C 03 D6 D3 AE 42 F4 52 F3 D0 0A 46 55 74
 CA D5 45 67 16 20 FA C8 42 93 38 E3 4E 57 F5 DD
 23 AF 42 58 D8 00 43 7A 05 01 FE B0 07 46 54 E1
 ED 8F 70 22 41 19 9B 50 95 27 4E 71 70 6F 26 CF
 CD 51 4A 67 6C F9 77 64 F8 90 EC EE C5 89 0D EF
 4F D0 C2 6A B0 E5 A9 E6 B3 63 32 D9 F6 4E AA CA
 4A D1 5C FA B6 9C 20 8A 99 82 DE 5A DC 6F E1 00
 98 F2 F9 4E 9E 87 42 0C EF 04 7F 2C E7 67 E8 F0
 4B E0 6A 06 20 A8 FB 24 1F 8F B0 9E B3 77 29 73
 6E 88 45 EA 92 78 11 4A FD D1 C6 18 0D 1C C0 22
 57 29 25 B4 11 FD D1 AC 23 3E 5E F4 D7 EE 30 CA
 3F 6F 7B F6 0A ED 2D EA 16 9A 9F 79 8E 0A FE D2
 C9 B6 64 5D 98 CF 02 F5 B7 83 10 ED 46 33 8F C3
 1F 38 D7 F1 D1 60 E6 AB 11 04 D9 4E A1 4B 19 27
 E1 AE 00 04 47 90 5D 00 17 54 DD CF 48 24 DC 3F
 69 5A F8 99 BA 0C DE 48 75 22 B7 65 F8 F2 95 0F
 E5 2D AC 0C 50 FA CC 8C 08 A0 84 31 AB F2 B9 9D
 B5 9A 3A 1C 01 B0 BD BB 8E B8 BD 6D 22 70 49 4D
 B2 D5 EA 06 93 E6 86 43 E6 1D 8E 09 2D C5 F0 3B
 DD 9B 52 C6 AD 58 07 E1 E0 15 BA C1 44 36 DF 4A
 C9 44 2E 53 0A B0 01 50 2F 45 83 58 8B 7A 86 70
 BF 6A E3 C2 2B AB DC 12 91 E3 83 A5 7E D5 EB 40
 75 56 EC 18 3E A8 CA 69 F1 F5 EE EC 68 59 E0 7E
 F0 D4 13 42 32 AC C1 C6 C0 19 78 C7 D6 F4 AE 09
 B5 73 5C 19 D7 CA 4A 55 F6 BD 07 34 1E 78 E4 70
 78 18 EA CE DE A2 9E 31 06 DA 58 57 42 9C 40 D7
 F5 B5 8E 7C 5F D0 60 31 31 12 7E 17 A1 38 2A 5B
 70 F5 81 8F F4 25 48 8C E9 9F 97 EA F3 D5 19 65
 49 FC 69 FB EC D6 74 89 F7 D0 89 70 04 1F E3 1A
 43 75 50 E8 2F 30 E4 0A 44 40 8A 02 48 33 D3 4E
 FC 1A 24 23 E0 06 32 55 0A 50 0A BA 65 FF 19 90
 9F A1 A3 74 1B 82 92 45 48 9F FD FE 19 EE A2 8D
 62 DC 3E EC 69 C2 49 AF 06 1F 9A 5B 2C B6 53 7B
 CA 9F 6C 71 C4 08 23 36 71 EF F8 8E 24 45 A7 83
 4A 65 4E 47 62 E3 B6 19 03 C6 C7 7B 79 9D D0 49
 43 03 26 DC D8 60 72 61 3A 95 86 17 E5 3F 31 F0
 79 57 63 6C 00 16 0E BC 6E 67 B5 A4 E9 3B 7F 30
 EC 79 91 D5 11 D1 0A A6 99 D4 5A D7 8C 1B 99 FE
 C9 3F 58 4F 69 9E 8D EA 24 6A 56 1B 2E DA 81 21
 74 E7 77 A9 E6 CA 98 FB 6F 5E 84 71 29 A0 E4 CC
 51 7E 85 42 3F 44 EB 17 0F 50 2C 18 C7 12 20 61
 6F 72 90 4C 9B 74 67 30 B7 44 EE 8B 61 8A 0A A7
 57 D4 04 8D 22 2E 5A D9 65 56 67 9A A6 EF 15 9E
 13 43 27 C2 D2 73 22 D9 ED 73 D3 8C 1D 1B F8 0E
 C3 B1 C7 C0 CC D7 87 2F 1B 09 26 45 4F E7 8E AE
 B9 30 F9 59 84 8B 9D 1C CE D7 66 E4 C7 F2 E0 4E
 71 BF 71 E6 19 0B 58 0E D3 1B E4 50 7F 0E 3F 97
 9B 5D 89 4E B9 EC 30 EE CC BE 77 A7 1C BF 00 B8
 4B B0 72 8A 30 D2 F8 CA 30 DD 23 84 3B BA BE 0F
 E9 F1 1C 9D AD A1 F2 8B F2 45 8B 6C 6A CA BC 97
 9E 35 F9 71 55 EA A9 63 4A 82 5F 81 DA C6 57 F6
 C0 A6 91 6F 9D DF E1 26 8D 8B 64 C3 01 9B 02 F5
 14 89 78 DC D2 B7 5A 8C 36 47 BD E1 7F 42 E2 B8
 26 52 3E 64 15 15 83 9C 9F 3C 0C 03 93 5B F0 66
 3A 63 BE 10 FB AD 8D 59 D5 D9 F4 C5 76 60 CE C1
 78 9D A6 1A B2 7C 93 0E A2 08 51 DE 75 EE F8 7B
 87 3D 8B 51 42 0B 64 2B 7D 00 6B C9 F7 28 9D 02
 68 93 61 CF A8 73 9D 23 B7 D9 E0 3C A7 DA 0C 26
 67 29 AF 28 E8 90 45 3C 91 A6 BB C7 A9 B8 5F 1F
 10 C9 50 FB D3 0E C0 A1 C1 48 7F DF 07 B4 2E 0E
 C6 26 6E 51 75 25 8A 21 5C 5D BB 33 33 77 8B 36
 7F 84 5B 9B FF AB 4F FD B8 E8 1A 0D 43 3D 6D 05
 45 7F AD E7 27 7D 23 05 FE 8D E2 6C DC BC 14 EF
 12 29 67 64 C9 0E E8 94 2A 0E E8 F1 7A FC 2C C8
 C5 0F 95 5E A4 E3 01 1F E8 6C 45 B5 DE 58 18 1F
 66 62 E7 B5 4D A4 0C B6 15 00 49 AF EF 77 4E 1F
 91 11 AC 68 16 99 82 D8 B9 CA 6B 81 36 D5 C7 8D
 C6 E0 75 61 76 E8 30 82 7F 5E 1A E7 F7 00 07 14
 F6 5E 5A 15 84 10 90 B1 DC 44 7D 90 4C CC AD AA
 E3 8B 4C C3 56 1B 91 9D 20 04 8A 5B B6 95 BF 59
 82 D2 F4 B0 DF D0 B8 83 F3 3C AF FB 6C 1E 7B E5
 E9 D9 99 BD 79 AF 91 45 2F 80 18 E3 87 DC 9E 31
 E5 C3 72 28 1B 18 60 7C E2 EF B0 5F 0A C3 4F A2
 63 2B FF AB 2A C1 AF 3F FB 6F 8B 05 C0 38 84 1B
 60 20 A5 0D D3 B3 8A C0 83 0B 3E 7F BF 22 DE 7E
 1F 22 C0 D3 B8 F4 5F 72 6F CD 4A D2 74 93 33 A1
 E3 B4 4A 38 2C 05 AA 75 5F F2 B3 EA 77 EF CC 6A
 D7 A8 F5 02 34 62 CD E5 5F 21 7B 50 83 BB 46 6A
 86 FF AF 0F 2A 50 D0 EB C1 8A 75 EF 0E 74 AC 95
 4E F6 AC 5A 8D 41 77 13 FA 24 FF 15 9D 0F 94 56
 9F 0A 57 F1 39 FF B5 E2 C9 BD D4 75 39 B1 05 4F
 1A 12 F4 C5 9A 52 79 F1 CC B7 59 B4 56 D6 1E 57
 59 F4 84 62 F9 36 D8 0A A0 2B C3 17 E1 2C 26 CD
 97 FF 5E 63 FA 80 8D 88 2E 47 74 BE DB 0F 3C 37
 E0 B2 90 3C 6D 6C 7E 2C EF 08 FB 9D 4E E3 3A 20
 67 91 00 E7 4C 56 41 F6 61 19 9A 80 B9 9F DB 5D
 21 28 6D 60 05 0E F3 B0 2B 88 35 9E BD 37 91 34
 86 BB 17 A7 94 A3 9B 26 76 99 F3 BA 90 65 D9 ED
 35 E8 1D E8 8E FE F1 03 3C 2E 5B 22 DC FA D1 D0
 70 C1 21 76 96 02 A5 48 6D 7C 4D 32 06 74 9A AB
 1B C6 61 EF 10 8A 99 C6 2E EF 3D B7 E7 EC B1 5D
 F3 A9 FC 6F C9 17 C2 0A 7D 9C 81 EC E6 10 64 A9
 C7 D7 51 FA B7 04 5A EF A1 00 1F A4 6B 55 52 4C
 F5 93 A1 1D C6 25 D5 39 8F B0 29 07 B0 FD F2 D3
 D0 67 A1 7B EB D4 43 7C 22 D6 5E 1B 1B 3E A9 1F
 E0 6C 91 F7 67 4A B6 B6 8C A0 F8 95 D1 36 58 C6
 47 AD 69 EC 37 21 67 BF 10 A3 A2 43 3C A5 28 D7
 42 52 A4 A0 73 6E F1 88 3F 72 36 05 D0 A5 62 13
 75 1B 3F 0E BD 15 65 FC 2E 84 13 51 77 FF DA 3A
 A5 B2 8C A3 F7 BE 7F 64 DD 7F B5 E7 D4 85 3B 37
 84 01 95 E5 9C 4C 3E 93 60 E5 48 56 1F 22 3F DB
 81 81 53 B0 57 D5 7B A9 13 22 1B 8C C9 36 FD DB
 91 18 AA C0 D4 00 9A DA 84 2C 4A A9 A3 C3 A5 40
 BE 1F D7 FA AA 6D 81 7B C8 EC D4 85 C2 A7 A3 B9
 81 A0 09 80 2B 3B 91 84 8C 47 DA A6 E5 0F 4A EA
 56 38 EE 67 26 25 AF 86 BA CE 5A 1A 47 55 43 C6
 80 79 C6 07 00 C7 5B E9 18 43 04 FD D5 DB EC 9B
 81 04 2B 53 60 0A FD 9E F5 58 82 21 61 69 81 16
 C9 6C 10 B5 33 5B 12 2F FE 66 CA CE AE 71 C4 04
 CB 03 9C 23 31 E3 4C 04 39 50 34 A0 BD 74 3D 48
 29 64 21 D8 A8 7B 15 0F 14 F7 6F 67 35 20 85 7B
 E7 5F 84 77 09 08 A2 6D 82 E2 98 2A A0 C5 06 8B
 FB 0A 74 51 80 05 B3 38 E5 4C FF AA 2F B9 52 02
 AC 92 31 03 C7 44 40 7D D1 B5 77 D4 38 AF D7 7E
 7D 37 54 C2 9E 91 64 B3 EA 3D FF 99 86 53 3E 51
 3F FF AD 91 EE 76 C3 65 8E 30 5F FF 36 B1 13 68
 AC 7A E7 73 89 86 88 C3 C7 FD 6E 5C 14 18 51 81
 83 B0 81 C5 D0 35 57 A0 C4 01 D6 48 D2 6D A3 E6
 F8 F4 99 83 1B 65 7C 53 5A 17 7D 9A A2 E3 D7 FC
 8D F2 16 FB CE 70 19 ED 9D 12 3C 98 EC 58 4B 5F
 02 71 6D 5C 65 14 CB 44 DE 1B 11 A5 28 DA 89 A9
 B9 6B 90 B0 EF 9F B0 76 2E D1 D4 7D C6 11 16 68
 EE 6F 58 E0 9C 92 D8 FF 0B 3F 8B FA 08 BE D6 12
 D4 28 41 F1 88 74 A6 0B DB 0C 88 21 43 E7 FE 29
 D7 CE 2C 9B C7 1A BA 1B 05 D6 9F 4C C0 85 7D 9E
 67 F1 AC 87 40 2F C9 A6 96 15 07 0E 4C 2D 0E B8
 0E 2F 17 0A 5F 35 41 34 95 0A 0D 55 68 6B 80 52
 06 1C BA 9E F6 B3 21 22 1E 03 87 23 78 ED E7 F3
 E4 26 15 E0 D0 AF 4E D8 AB 12 34 68 FC 11 7A DB
 66 A5 7F A2 83 53 D1 90 FE 10 C0 C0 AD 00 45 86
 A0 60 88 55 0A A4 26 8D 50 65 77 A0 A7 4E 1F F6
 1E A3 B0 3F 1D EF 50 3F 60 76 E4 61 31 66 D9 A4
 A0 34 C7 CB F0 DB 8C 68 6F 2C A6 2E B6 BF BB 16
 27 49 03 ED 22 EC FA FE BC 01 0C 48 E9 1A 52 74
 01 C7 43 9E 24 E9 2C 56 BE B2 40 60 24 7D 0C FA
 8E BA FA 41 46 F9 48 14 A2 BA 76 AB 52 04 FE 33
 BA D5 E4 BA 0C A6 62 0E 10 B3 AE 6D 5B E4 F9 07
 88 35 A6 A2 33 1B EA 5A 85 78 56 5A 10 39 1F 22
 51 07 BD 3F A4 F9 2E 02 CC 17 A9 6B E2 54 DC F9
 45 D5 B2 7B 41 0B 52 DF 08 44 12 0A 84 A5 CA A3
 E5 35 03 F2 42 49 5F 24 E9 EC C6 C9 F9 D9 F2 2F
 3C 9E EF A6 A8 5B 7E 49 B5 20 CD 18 BD 3F 3B 15
 AB 74 A5 77 3A F0 8D C1 CB 73 45 63 EE 71 C3 F5
 C4 CE 45 E1 37 8D 49 FE B8 59 82 57 50 E0 EF 4B
 B7 FB E2 7E 67 3D E1 6C 9A DA 01 B6 81 C8 A8 9E
 7F 04 7C 6C D8 AC 39 B8 36 1E 73 FC 83 32 DF F8
 61 80 85 58 95 50 14 4C DD FE C6 76 D4 0C 32 4F
 CC 07 87 9A C8 10 4D 0E BD 00 CC 88 F2 6D B3 C0
 83 DB D4 5A 25 CB E1 E3 87 79 FE 71 DB 96 55 42
 A4 80 7F A0 BA 7C C8 A6 8B D8 C5 0C 4B 2E FB 5B
 EA 13 1C 95 A1 34 4D AC 7C 5D DE AC CF DE 9E 1E
 B6 8F 62 F5 05 72 00 D2 56 C7 0F FD AD AF E5 42
 A3 A2 BF 67 CD 75 97 F6 FC 65 3D 5A 15 46 71 8B
 DB FB A2 AB F1 E9 30 75 40 79 54 51 B3 E9 71 01
 22 71 80 54 9C E4 8C DB 14 42 32 83 8D 37 D6 CA
 AF CC 62 68 9B 17 AE 04 F4 12 69 0A 78 CD E7 6A
 DA 68 9D 13 3F 09 32 77 5D 2D 18 AF CD BC 56 7C
 A8 C6 FC BC 22 C8 1E 9A A4 14 87 B2 A0 EC 7B E4
 20 1D 30 25 4A E5 52 26 10 11 A1 85 27 29 55 1A
 86 CF 35 DA 01 32 48 CF 70 7F B4 F9 A2 87 99 78
 0B D7 79 F2 11 91 22 F8 84 F6 54 73 CC 47 5A 1A
 F9 B6 59 EC 15 DB 2F 69 85 E7 5E 38 C0 40 A1 AB
 85 A9 39 A0 C2 3D 82 C7 42 C3 46 9F 5E B5 7D 2A
 5C 52 92 CD FE 64 55 65 C2 16 5A 6D 1A F6 A6 56
 F1 0E 17 01 4E 4C 37 76 74 4B C1 89 A7 BC 40 DB
 9B FB BA 61 54 25 08 C3 1B A2 9E F3 AD D3 9B BC
 3E B4 84 BC D7 81 9B 97 70 69 BA 62 E3 C9 F3 68
 53 A7 39 06 B5 49 6D E9 E0 21 B7 71 45 17 D4 AA
 FF 58 1D 4D EA 73 E7 BF F4 17 39 22 EA DD FD FF
 94 7F 5C 91 1E C6 2D 03 AD 4A 0F EE 2C 9B A2 A7
 A5 E8 5D 21 34 E0 68 21 FF C6 BF 17 16 DA EA BB
 78 AA D4 18 DE 23 BC 17 E2 22 D7 8A 47 F4 8B 6D
 E4 A0 B1 C1 15 F0 32 AF B8 2F 77 B3 A8 4D 6D 59
 9F 0E B8 3E 20 81 D0 B3 5C 74 B5 56 FE A6 46 AC
 3B CC 7B F9 7D 27 14 77 A2 1C D6 A3 88 12 F7 58
 A4 76 74 4D 55 A5 28 4C CE CF 21 1C 87 D2 99 51
 A7 6C F1 98 DC AA 0F 5C D1 05 6A 86 4B 2B 27 73
 EF D0 E6 C6 D8 3F AC 4A FF 96 46 A0 8C F6 76 A4
 47 01 1A 01 02 57 22 B1 24 06 DE 43 E4 0D 4B 84
 B4 4A F9 A1 03 48 85 C7 46 28 91 C7 DF 61 F4 72
 F6 B7 9E 73 13 57 EF 60 09 EC 70 E1 D8 6C B3 B5
 17 06 2C 3B 2E D7 C2 39 CF 3F 0B 10 EB 5F 4B CD
 BC 2C 21 59 93 16 6C 56 B3 D1 C9 8C A1 86 01 DE
 4A C7 8F 95 82 A0 5F 96 86 18 0B 48 33 2A 96 D4
 DC 77 AF DB E9 D6 89 FA 63 D7 3E A0 D2 07 22 A4
 FC F2 C9 3D FF F6 FB BB CA A5 A1 97 AF C3 05 92
 7D 7A B7 F0 96 99 88 D0 4A C2 5C 5C 65 3C 68 4F
 75 8B 0C 16 D6 77 2D 4A 0C B1 15 99 08 B9 BB FA
 BD C4 21 46 52 32 F0 A2 3D DF 8C 59 21 94 FB CB
 62 3C B9 F1 49 9D A8 74 54 66 9C 68 A9 6C FB 1F
 9A 78 32 AC 05 9D 1D 81 85 3C 37 27 FA 1A 44 12
 A5 BA 8F 28 25 93 04 11 6A F0 8E BC 22 FF 49 0B
 88 5E 44 DA 61 E3 E7 FC 09 3E C6 EA 16 BE 93 AC
 E1 51 56 66 FC F0 48 E7 36 5B 52 72 DB 5E 9C A0
 67 EB D4 C4 CC DB 26 A7 65 1E 20 5D 0D E6 05 38
 CC EB 84 11 7C FB E6 01 62 58 AC DD 3C 2F 1B 13
 0A F2 A2 DC E4 40 06 D5 B5 DF 69 31 30 07 49 C6
 29 F3 3F 65 28 5B E1 3F DD 7A 6C 17 45 44 3A F3
 34 80 7F 23 FB 7E BD E5 03 DA 9E 33 A2 A7 01 17
 21 94 10 91 14 FF DB B9 79 71 47 71 1F B6 9B 47
 A8 8E E1 E8 21 2C 89 22 51 3A 16 74 84 AC EB 79
 C8 AA EC A2 B6 6A DB 5A C3 05 E0 95 5F 3F F3 84
 67 8C 8D 71 07 5D 27 2C 0B EC 8A 2C 59 52 27 9D
 90 86 3E 78 B9 0E 38 BF B7 67 42 C4 5A 6C 9A 60
 7F F6 3F 55 15 55 AF 0F 2A 4F 22 7E 0E 0F 10 5B
 A4 EC 28 06 CF 12 3D D1 3C 1F 97 A5 1E 92 9C A6
 01 AB B2 EA AC B0 BF 2C A5 82 37 5E 56 BE 07 3C
 27 0A BE CD C0 EC AE D5 33 07 41 B0 AE 79 32 D8
 9D 6B DE E5 37 30 A3 EB 96 CE 46 11 BB B2 0F 01
 FE 14 6F 02 4A A2 B7 5D 1E 78 86 FC 9F 74 DA F7
 CE C3 4E 1F A4 58 AA D3 FE BB 0B 38 AF 7D 87 F1
 EC 1B 07 FD E3 36 A5 70 60 3E 10 66 B7 CB FC A3
 07 4D EE EA 40 BF 48 15 58 6A A6 05 3F 0D 09 F5
 74 40 E3 08 0B 6F 70 3A E1 E4 A6 EB 24 C7 C5 32
 2F 4D D0 89 7D 3D B9 D5 58 67 C1 36 0F D7 10 E0
 2C 90 4E 00 FE E2 06 7C F6 57 01 09 46 2D 91 5F
 DD 1A 4B A2 48 77 57 AF 64 50 19 4B C6 B3 42 E7
 A5 DC 25 BE B8 5A 23 59 0A 22 CD 58 5C 57 F0 73
 43 7A CB C8 3F C0 5D D0 A7 C9 40 AF 70 05 D0 42
 4D 9E B7 3B 4E 61 E9 55 15 20 6B 2A 5F 68 23 35
 F7 72 23 4D 1B B8 70 D6 B7 56 29 12 4A DA 5E 17
 65 BE 99 D5 55 75 66 9C 1A 5E 95 FB E4 73 B6 8B
 8E 1C 75 E1 B4 EB F7 F2 E1 B2 65 F8 49 BC 3C 70
 BF 3E 7F D7 CB DC 6C C7 CB 2A AF 8E 07 9D 60 49
 7F 1C 48 99 5C 94 3C 56 9C 6B 61 B8 05 80 8D DA
 38 D7 F8 5F 96 F8 7C 88 83 B5 E7 81 18 90 F4 53
 B0 F5 3C 9F A6 7D A4 1C A7 4B F6 78 47 8A CB 92
 37 89 00 62 E2 28 21 27 5F 1D A8 67 E2 F3 C9 6F
 4A 0E F3 2D EE B4 2A 33 4D 54 8D C4 AF FE B1 ED
 AB 1F 9C 61 70 D2 A1 DE 9E 47 F0 BC 30 4F 4B 6F
 68 7F 2A 8B AA 57 CA 91 42 78 41 AF 8A 19 0F FC
 EE EA 73 0F 37 F4 98 77 57 94 7F B4 73 2C B8 05
 93 16 E8 0B 4F 0A 8C 39 B7 C3 F3 2B AF 40 AA 6C
 D4 0F 2B 8F A3 ED 21 78 FD 19 4B AF 12 B3 99 6C
 E7 74 A7 6F 69 92 A9 BE 2C 2A C6 3D F1 46 D8 DC
 6A 4D BD C3 F5 8F 28 80 2F ED 15 3B F1 74 1D A2
 4F 30 4E 83 3D 3D C3 4E BB E2 8D FA 36 F4 C7 B1
 DB 36 2F BC A6 CC 94 A5 BF 13 93 05 1A 37 A1 5A
 55 9A DB 65 3D 00 61 14 A4 13 3F C7 94 E1 B6 15
 B2 D7 59 B4 F2 42 33 14 C7 5B C7 24 6E FF 17 21
 E0 0B C7 56 E6 E9 B7 80 78 E0 B6 16 FD FE CB D1
 42 9B 52 BF 3D 60 85 9C 52 37 0D 36 E6 DC 3C 9E
 8E 32 37 A9 36 82 39 8D B7 61 08 49 CD 1C 40 2B
 21 5A 62 08 2E 17 98 2F 5D 0A 8F F3 B3 5E 0B D0
 7B 7E 18 32 C3 66 69 7F 07 EA 41 06 4B A2 18 66
 B9 DD 64 F7 28 EB C8 3B E2 98 7F 6A 1A 08 26 06
 48 69 8A 0C A5 0D 76 7D E1 4C 18 31 5C EE 2C F3
 74 54 F7 6A 19 03 68 A3 80 DD D2 04 28 53 67 5F
 C1 FF C8 2C 07 1A EA FD C9 08 1A 0D 6E 93 94 E1
 C4 09 18 4A FD 0D A3 CE 76 99 AE BD B9 81 EA FD
 F7 10 9A FE 81 9A 9E E4 AF E7 E0 B0 E7 73 2D 2B
 81 C6 E7 95 52 14 D6 F1 C4 78 6D 91 25 86 A4 70
 F8 47 2B AC 81 0E 16 9E E6 F1 F3 32 3E 09 1A 67
 06 47 A3 DB 72 F8 D6 BC 4F 85 4D 6C 92 CF 99 A7
 05 5C F0 01 87 7E 85 9F F4 39 CD 25 A0 98 83 71
 C6 05 07 94 5A 11 60 49 38 FE AE 1A 9A 27 7B 5B
 8A B1 4B A3 CC F3 CD D3 37 CA 8F 32 C4 75 36 84
 95 FC 3C 8F 6D FC AF B9 36 2E 66 C2 40 D1 BF AA
 E7 E1 95 AB 7B BF E3 35 64 91 D7 4E 72 EE 41 69
 C2 33 32 40 41 80 53 42 8E 99 59 1B EE 95 96 19
 B0 3C 9A 55 38 0C DB 3D 36 A0 63 0A E4 C2 0B C8
 7E C9 47 3F E2 15 D2 40 2E 97 74 5C 79 BF 6B 5D
 E6 42 E0 26 07 11 38 44 F4 1C 34 4A C4 64 C3 37
 36 3C BD 22 CA E7 E4 4A 31 DB 14 EA 05 4A A0 41
 D9 E5 08 7D 83 A8 69 BD 69 01 84 2D 59 EF B3 01
 9A F6 AE 6F 48 74 73 FD F7 E4 F4 36 36 7F DB 82
 43 E7 91 FD 00 B0 D1 8D 2A 9F F6 6C 75 5B 1C B7
 24 CE A2 2D 95 A4 EC 88 CD F4 57 A8 84 1D C6 ED
 4F D5 6E 68 79 70 70 FE 7A 41 7C C3 5D 3B C3 3D
 B4 AB 99 C7 81 0B 53 79 81 99 FD 03 B3 CC 41 1F
 5B B4 49 D4 9A C5 74 5B 6F 3F CC D1 1E 80 71 B5
 B5 A7 7F 78 3B 25 0C 69 5C 4D 85 16 C4 33 D0 93
 AA 79 10 01 33 04 4D 6D EB B1 12 D9 A7 CA 47 05
 E7 36 BB 9D ED 79 12 5E 86 B2 D0 6E 56 29 9C 65
 10 14 B6 B9 D2 A3 A3 0B 10 0A A2 B1 29 A3 AB 95
 37 FE EA 66 A3 1D 16 25 DD 9E 39 1A 49 1F 8B 64
 85 C1 82 46 2A 05 50 7C D8 6B AB 14 BC 28 D9 0F
 2E A1 5D 6C 9F 93 AB 86 0D E6 6B 00 3C 5E 32 A7
 62 AB 25 F4 36 54 28 FF 8A CD BA CD EF 3D 47 2C
 7C 1B 2F F4 BA A5 B0 DD 4B 49 03 E8 F1 5A 41 A6
 44 4E 12 EA E6 3A EB CD 4A C8 38 B3 45 D5 CD 34
 1E FF 75 A6 53 24 2D 17 3C 2C E2 D3 41 3A 82 BB
 01 4B 12 12 FC 3E 59 CD 3B FA 15 F2 80 4A DE BC
 DF 3C 95 9C 32 DE 82 40 F3 CA 9D BE FE 51 06 6E
 7F 42 46 47 BF BE 32 4F F6 03 7A 11 46 76 DF 75
 F9 B7 95 56 B8 C3 96 C8 F9 8E 36 3C 14 A3 ED 77
 BF C0 DA A1 11 0C C8 57 3B 60 A8 E4 48 AC 7D 83
 FB 19 FE E9 0F EC FC 33 6C B6 BE 29 5F 45 59 94
 3C 94 B0 09 13 7C BA 9C 03 82 62 C9 EF F8 32 EF
 B2 1C BC 74 95 E4 23 82 E2 37 8B 26 5B 7B EB 82
 25 BC DE 6B 6E 52 55 8E 7F 22 5C 16 66 A6 CF B0
 60 B5 B3 CC 73 02 63 44 91 54 15 BF 51 95 C9 B3
 76 D7 97 27 15 22 F3 EE BA EC A8 C0 5B 39 8F 0F
 5C 58 FF 11 8E FA 40 58 ED 98 32 EB CB CA 15 4D
 A8 99 E6 FF CD 0D 78 B6 D2 89 01 2A 05 52 69 59
 31 CD 5E D7 CD 40 89 C2 1E A3 12 77 A8 90 56 CB
 FC D8 A4 00 60 DC BA 21 D1 82 15 62 0B 28 72 E2
 20 CA 9E 98 04 A6 D0 EB 7F EF 5A 75 40 29 11 88
 09 EF F6 3E 98 06 4F 28 0E B4 2B CA C4 65 FA 8C
 DC B8 4B AC C0 55 A4 1A 56 76 57 CC 7A 81 C6 83
 CD 67 E2 76 C9 23 95 10 C0 1A 62 C5 2D FF 88 E0
 2F EB AE FA B3 EB 9D BE 83 5C BC 5C 40 0A 97 3C
 A8 96 FA 55 37 23 17 98 EF 5D 68 71 E6 80 6F DA
 02 BB A6 A6 77 C2 EC AE 10 DA 95 B1 73 E5 1B 8D
 CA 49 9B 24 61 B1 E5 76 3E A0 D4 DA DE CA AF CC
 95 D9 9F 5C 87 78 99 0E A7 02 B7 F3 C3 FE 55 50
 7C 47 FE 63 A6 C2 42 83 A3 89 6F 9D 8C 5F A9 D6
 B0 79 76 BD 18 A7 AA 4F B7 25 D4 85 F5 38 90 8F
 F9 DC F3 EF 7D 2C 42 80 EE 7A 05 CF 5D AA 74 B4
 6A 3A E6 4E 7A E4 DC AE 9D 62 48 51 A6 6D BF B9
 8D BD 3F FF CF 24 B5 22 BE 2A EB 02 EB 0C FA A5
 96 E3 F2 7B A2 52 DA DB 08 9A 1C 18 D1 17 A5 68
 4D E4 DB 43 20 AD 67 3E CE DD D8 88 C3 00 F7 0B
 C5 A2 02 86 6A 8E 07 F9 3D 40 44 04 65 40 28 FF
 09 C1 D8 C0 84 C9 95 09 92 88 13 84 CA A1 71 F6
 EC 43 B3 73 0A B6 24 83 1F 89 7C 5F 64 9E 37 72
 06 55 3E DF 0C 53 13 C7 E5 B7 20 8E 73 C2 0F E3
 11 DB 27 6B 93 2E 0F EC B8 3E C3 6B 58 49 0E 74
 BB C2 A5 42 F2 7E D4 67 4C 31 15 9E BD 77 01 26
 CC 6A 02 43 25 98 F8 C4 6C 76 27 28 76 E8 25 4B
 DF 82 AE BC C0 64 F4 9A F7 C6 47 11 33 F5 A6 94
 DF 59 4F B4 B4 8E 02 90 8A 9C 2F 06 F6 30 4A 13
 F5 87 F8 15 3A 9C 1C 77 47 FC 71 04 B1 4F 81 26
 BE 98 15 2B 33 B4 3F 2C 08 01 D6 07 83 41 EF E1
 C1 BA 65 21 6E 5D 46 17 52 CA EF 4A 27 E0 B4 B3
 59 73 BA 96 D8 5B 2A F2 C5 AE D8 62 4D EE 04 03
 DD BE 41 8D 23 09 47 9D 6A E9 F9 E8 8F 88 BE C0
 52 78 E3 03 D3 A5 C9 B7 D6 38 AF 5E 75 32 0B 3A
 C3 03 AF 58 61 2C 66 40 88 E1 D7 0E 33 8D 1B 8F
 60 59 80 F0 D7 A7 26 7E 56 81 C0 A0 55 D5 66 4D
 FA 10 24 F7 3A DE 0F 97 3B AF E6 DA 05 62 CA 3F
 86 C7 A6 8F B7 2D 53 12 A0 05 2A E2 2F 17 53 DF
 FF 1D C5 EA 99 0F BC FB 4A 95 65 5F 2E 14 D8 E4
 F7 76 B4 ED A8 BD 4C 5D 12 06 C1 FF 23 B6 83 48
 1E A7 4A EB 07 2A 7E 13 88 DE F9 C4 63 94 BA 27
 33 F5 20 17 CB 5F 86 97 A4 07 22 7B F1 64 2C BC
 22 6E F6 62 BF E7 CB 9E AA EB 2B 1E 59 05 4E CD
 46 6E CD 44 BC 11 9B 2B BE 9B 6E BB 34 DD 42 80
 22 84 33 98 B2 C8 75 A9 A8 BF 13 06 A8 A1 9E F1
 B0 EC 09 20 DD 8C BC 64 0B C4 38 87 DB FC 61 44
 87 BD D6 66 32 AB A0 9D E5 96 9C C4 C2 2D 6D F7
 14 AD BE 05 68 23 2B 9B A8 86 C7 A0 9D D2 EA 84
 87 05 9D 21 C1 C2 D8 16 43 5A 05 E7 96 14 A1 FC
 BF B3 27 09 2B CC B8 70 D1 92 34 00 F4 8A 30 0B
 5E 9B AF 8A 42 C6 34 D3 8D 43 70 BE 03 6F C8 09
 A4 9A BB DC 02 C9 07 34 C8 C9 D2 DF 80 CB C4 1C
 48 69 AC 76 8F 7A 7A 84 02 F6 19 E0 20 4D 16 17
 89 ED 62 4C BE 41 F3 B5 89 50 41 37 B9 AD 60 34
 AE BB 86 E9 D1 A1 9C F5 83 66 D6 6E 94 D9 39 4B
 A8 F7 17 1C 77 FD E1 F3 76 EB 88 24 4C 88 A6 20
 64 41 61 FC E2 C2 82 88 C2 58 81 D2 63 E4 B2 47
 25 1B 03 1E 52 B9 F3 A6 1F C8 A7 42 38 C5 78 39
 3B 93 3E 7E 7F 35 7C B3 ED 75 29 E2 12 6E 1C D5
 EC 4A C2 5C 3E FC C3 2A 3D CA 93 50 21 4D 06 12
 93 BB 01 E8 30 3E 5C AD 78 A9 5F B1 4D 11 5E 74
 18 24 26 B5 09 58 4F 06 5E 07 0B 7F 95 81 B1 C0
 A9 A4 ED 75 6A 05 8C B1 E3 B3 7E 89 A1 1E FA 87
 B5 5C 06 6F 9B FD 01 D1 C4 11 46 4D 84 79 1C 94
 42 22 56 16 F4 91 D1 1C 3B 56 F7 AD E2 BF FC FA
 76 EA 0E 42 2D C7 57 EC D2 9C 38 47 D7 5B F7 80
 BF E1 E9 CA B1 C2 74 37 AB 69 05 89 97 82 3B 1E
 67 30 63 D4 FB 0F DB D3 86 DF C2 2D AC 51 46 88
 15 52 7D 9E E3 DF 88 D1 8B 84 57 5F B0 0D 48 27
 57 0D AD AE 49 93 3A 08 BF CC 66 7B 85 48 AB FD
 0A FB 74 BE 23 96 21 07 85 37 00 28 58 DC 7D A0
 39 5E DC 89 00 5A EA EA 2C 67 F2 EB 40 11 94 BB
 C6 AD B4 D9 C1 69 EF 3A C1 54 3A 85 40 08 40 52
 E5 E6 A4 0D 11 05 8F B7 66 B1 A3 73 99 E9 BF AE
 F8 AF 98 EF 56 95 50 20 EA 39 D0 AE FF 58 B8 59
 FF D4 7D 01 F6 1E 6F 3D 3B 1A 69 FA D5 21 9E 61
 CB 37 40 FC 5C AE BF A9 DF 6E 70 5E 95 78 26 E6
 C5 45 3A A1 BD 29 8F EB 43 58 C5 E4 7F 59 E8 28
 7D 9B 11 83 5A 12 FF 3D 70 07 5E 43 A3 6A 69 92
 52 B8 4E 1D A5 45 9D 83 30 A9 61 9A BA D3 A5 8C
 F9 5B 71 23 00 94 78 DD 4A 8E 42 6F C4 BC D5 B4
 88 C1 FC C0 FF 48 CC 6B C2 DB A7 E9 E6 FD F5 F1
 DE FC 08 8D EC 09 DA 4D 6F 98 B2 C6 54 4E 5E BF
 55 39 B2 FB 29 3D 7B 0F BD 34 A9 0B 33 BD 7A B7
 D0 51 AE 6E 3D 54 E9 A8 59 D8 CB 44 E9 93 2F 5C
 F5 15 93 76 90 77 C2 72 3C 0A FC BF 4C B6 D1 4A
 72 71 9B 10 70 B8 BA C0 2A 33 68 0F 52 3D 3F C6
 08 23 2E EB 10 FE A1 87 2C 41 80 99 60 8C CF 45
 41 33 2C AA 18 9F EE E3 54 30 1F EA 86 F6 12 B8
 96 47 E9 41 7C 9F C7 AE 18 5B D7 6F DC 51 8E 1F
 CF C4 7D 4B C9 9C 0F 4F AB EE 37 50 29 A3 A7 35
 89 ED EF F4 AF D4 D7 2E 17 C1 B3 35 A3 71 31 B6
 C7 11 F4 40 73 C1 66 43 7C FD E2 6D AD 6D 02 12
 03 D8 D6 D1 B3 73 60 40 79 D6 7B 21 BF EF 84 B9
 C3 9E DF 60 19 EB E8 67 72 13 E7 13 48 3C FD 30
 5A 18 4C 87 A5 87 6F 44 95 C8 3A 51 09 58 23 02
 76 29 30 40 16 9C EB 4C B5 A6 D0 07 57 56 35 11
 62 9C 27 44 D6 67 CB 86 D0 F0 42 D9 24 AF 4B B3
 1B 88 35 54 B3 C9 CC CF EC 3B D6 CC 9D 48 BC 38
 37 AB 1B AB 99 E9 B2 79 E7 A8 A1 C6 88 1C 2E 2A
 45 B4 80 EF D6 0C 75 B6 F2 BE 14 B0 EB 0B 14 54
 89 0F 26 F2 79 DF 7F 04 49 34 01 F3 05 2E 6B B3
 87 A2 01 78 AD 3F AA 0D 97 B0 0F EE BF 97 C7 DD
 3F 3B B8 C9 6F 83 2E C6 26 D1 94 8D D1 14 FC B7
 40 1D C2 51 93 BC A1 96 CB 81 DD 95 2B 05 C5 84
 AF CB E5 60 4F DE EF 99 B6 C2 4E 26 FD 27 F2 81
 E7 4B AB FA 8F 96 B1 3B 0C 6A 43 FB 2C BC B5 76
 F2 24 2B 7C A8 CC 99 0A 68 4E 1B 20 F8 C1 EF 66
 F0 96 DC 22 75 21 7B B9 B5 EE 55 71 68 78 7F 3A
 04 D4 1C 58 97 BB C8 9E 65 B8 16 75 83 16 AC A0
 6D EF 0E EF B9 84 E6 FB D6 40 22 21 EB 2F 4B 4F
 80 79 0B 9C 49 1C AC 96 0B AE 1F 72 F0 49 E2 2F
 65 BF CC 9C 21 8F 24 7D 87 B6 05 93 B6 FB 81 E3
 17 78 4F C4 E8 BD 93 92 B1 E9 B7 FE 08 96 56 08
 CC D6 79 07 73 81 F3 5B 8C 90 7F 42 FC AA 45 84
 F6 2F 20 C6 9B BF 5F 43 D1 DB C1 45 81 32 71 6E
 98 99 80 82 64 AE 06 C7 C9 0B BB 0F 9F 1E 52 8A
 4E F2 EF 1D 4E FE 50 85 66 83 FD 74 69 29 9F A3
 DC 9F F5 03 04 33 AD CF 59 9B A2 04 A3 DA 53 F2
 3D B7 20 B3 B8 1B 2B AD 83 5A 1F 7E 99 0F 31 90
 38 E7 B9 82 35 C1 BA E9 E7 FF F4 0E A6 25 CD B8
 84 C0 23 1A 44 88 2C FC 33 00 D2 46 A1 FB 81 EE
 AA 93 D2 C3 D1 23 71 CD 8B 51 4C BE 10 5E 42 34
 AF 24 5A 8A 3A 1C C8 42 27 A7 5D 86 A1 0E 80 DE
 ED 0F 14 9E 38 8B F0 D6 93 D4 21 FA 4C 62 D7 0D
 38 A2 D4 BC 59 49 62 BD D9 91 F4 CB 42 D5 9A 04
 DC 35 00 74 73 F8 15 34 1A C9 06 F3 53 FD EA 91
 3E A3 CC 40 26 72 5A 30 FD 55 5C C9 5A 02 CE 0D
 B3 9E 1B 1E 99 9C 6F DE B9 77 80 A0 E0 B0 D7 F7
 A1 9C E7 28 EC F9 CA DD 5B D2 82 28 B3 C0 CD 3C
 02 87 60 A5 93 C0 4C 8C 04 F5 A1 33 2E 09 1A E9
 65 BE A7 84 88 9A 45 80 41 29 8E C3 FB 90 D0 41
 D9 CA FC E6 74 11 53 1C 34 6F 8F BA 78 CE D6 E0
 91 6B FD 1D 76 DC 1A 87 3E 3C 40 96 94 90 13 32
 9C 1A 3B 45 B3 05 0F 9B E0 48 B0 AE C0 91 F0 6C
 6F 43 66 2A DD 37 B5 F0 AB 18 8C 1A AD 18 2E 97
 31 51 FB 4B B6 3D 98 DC E0 F4 4D 71 84 72 B9 2B
 3F 8A B0 AF 21 A3 CA 54 FD 50 6E AC AB 11 2C E0
 3F CB 31 0C AD 17 4F F6 90 AD B7 3F 05 23 82 66
 EA 09 65 39 0E 32 3C AE E4 E0 91 1A F1 ED 1B A7
 A2 A8 83 7A 42 0E 1E 49 53 C2 83 2D D6 CF DB 02
 56 7F F2 E6 0D D5 34 CB 12 DD 90 16 61 54 5D 0F
 8C 4C 8C 2F 28 76 11 F4 43 AB 42 F5 1F 2B 24 46
 5C A9 50 1A 27 FC 0A DC 5D 6F 5B CF 3B 95 24 4F
 99 02 E6 56 E6 97 67 92 99 A6 A0 D0 02 6A 32 6F
 C0 48 C9 9A 8E 1E 87 89 7A A0 68 9B CF 0B 02 21
 8C EA 7C 57 80 CB 41 07 92 12 58 1D 46 B3 6E 0E
 D5 85 CA 6D 21 AD AF 86 2B A9 9C B4 75 46 86 CD
 F6 F0 95 68 E3 3A 21 9E 99 CA 69 A2 B6 2B A5 3F
 31 87 5E F9 D7 B7 9F 38 20 FD 12 6B 60 D6 2D B5
 4B AF 9B C6 63 7F 8C 48 BD EC 08 D3 10 EE 60 DA
 E8 72 09 16 92 FD 54 1D 95 66 5D 85 4A BE 0F 17
 7C B6 D9 82 43 C4 1E 6F 60 0B 35 16 61 45 C9 F9
 13 05 C2 6E ED 6C D6 5E 28 11 1A 56 AF E7 D1 86
 55 51 34 44 D4 93 8A 5F B1 AF B3 04 65 03 F4 32
 01 AE 4D 69 DD 2B 1A 96 FE B5 B8 31 34 3D 6A 29
 B3 25 75 90 D0 B3 DF 7F 8F 52 F3 BA 73 8B 95 F9
 17 F1 DF DB 54 4A 1C 49 D1 64 38 2A 95 80 79 88
 1D 2D FB 1C 9E F8 0F D1 C2 0F 04 CA 82 4E 95 4C
 11 E0 81 2A DC 89 62 E5 5E 2B 01 D0 91 2A A4 9B
 15 72 10 DC 33 84 BB D9 5B 7C E8 54 05 5D B0 88
 5E F4 23 74 78 92 62 5D CA 8B C3 2B 81 A3 66 77
 1A 24 FB 3C 58 6D 7E FC 14 3F D3 97 B6 1B BD 7E
 77 98 D6 63 EA 19 91 19 3F 4D 06 1F 56 7F BE 08
 F1 77 3E E3 1B 34 DF D4 53 CB 56 F1 B5 26 BE 1F
 C7 A4 1C 24 17 B5 2D 95 13 6C 91 5E 63 FD FF 5D
 6A 72 29 3F 90 72 38 0B 42 11 18 D9 80 31 60 EE
 07 8B 90 B7 9D 81 20 9B 63 CA CA 0D F0 9C 51 A9
 76 12 2A 4D 32 FA CD AA 0E 95 EE 17 BF BF 1D 31
 E5 5E F1 8E C6 21 9B 1F 00 F9 88 93 9D 1D F5 AC
 ED 59 10 C7 1F EF FE 64 EC DA F7 6A 1C 18 75 0D
 7C 07 06 26 62 5D 56 BB 30 7C 4F E2 74 AE 34 CC
 78 2D F7 B2 9E 33 8A 0F 30 D1 AF 4E D2 C6 71 D1
 01 71 60 4B A8 54 71 C8 69 56 93 0D EE 8C B3 46
 E9 8D 80 72 B4 6E 80 A9 3B 92 E2 AC A9 DD DA 74
 F1 1E 34 88 27 5F 3A 79 68 13 58 9D 0C 17 94 0C
 6F 4D 94 52 7E 4F 9A 8B B5 41 BF 58 04 C5 7E E6
 4E 8D 10 2D BA D1 32 A0 C2 8C 92 B8 3A 80 F3 C1
 E9 79 31 15 AE F7 55 F6 B6 3A 2B C5 79 55 81 22
 9F A1 8C 97 C1 FB 11 73 86 BB 16 5B 99 A9 E2 27
 B1 83 85 6C 77 C9 CA 4F 44 D6 9C F6 2F 81 EC 29
 17 54 F7 25 76 00 A9 A7 F8 91 97 15 8F 98 5B B7
 38 35 C4 66 D0 DA 90 6A 03 3B ED 9C C9 88 DA 03
 DD 4F 2B 35 34 B5 D1 22 35 3E BD 59 ED 5A 9A 39
 A1 49 01 71 3B 9B BF 58 66 8F FB 8A 20 41 24 D9
 A3 88 94 7C 13 0B F3 B6 ED BA BF EE 0B 70 D7 E5
 1C 2F E2 17 7D 2E 23 7D 29 57 65 05 47 C8 0A B8
 86 80 5B 49 41 23 7D 5F 89 68 9D 4A E7 E8 A6 58
 76 42 53 75 3C FA 9F DE 82 87 2B 60 52 56 87 6E
 38 FA 33 CB E5 5C 39 77 BE CD 67 A5 1C 0E 75 8C
 28 71 A0 7B 3B 12 AB CA BD D8 A6 FA DE 99 6A CB
 C7 75 02 97 32 27 5D CC B5 50 8D 72 25 1F 85 91
 F4 15 7E 96 6F 12 4F 51 20 96 D1 DB F4 8C 91 B0
 F0 C0 94 D5 13 63 E6 C6 9D FD 38 60 A6 5A D3 F0
 26 97 72 9E DE 56 F6 02 D5 55 0C A4 84 60 87 D8
 B0 C6 BF 38 C7 EA 97 C3 00 7A 00 18 C5 92 7F AD
 B5 B3 06 2F C4 EE 40 61 23 D9 71 91 71 8C AC 58
 26 0A BB 63 7F E9 E9 F0 6C 31 1C 78 BE 3F E5 D7
 1A 1D 08 68 98 11 21 28 93 03 33 63 3D 77 70 B0
 E3 47 72 11 83 6D DA 48 1B 0C BC 79 74 9C 18 57
 68 AC E6 BC A5 8B 80 8F D2 A2 17 65 AB FB 5D F0
 0A 90 17 D8 AA F9 50 55 21 2F 3D 40 87 42 10 DF
 15 4A 8D 1A C2 19 9B F2 3D 1E 23 0D 6D 42 47 A1
 A1 FC 30 6E F7 F1 1D 50 98 5D F6 7B FB 35 6A 12
 8F 80 42 91 77 6C 70 B4 9E 86 98 9A F9 31 5C 38
 0C 8A 84 6E 4A D8 2F 02 F9 9E F4 40 BF 0E B3 F3
 12 4A 33 74 A2 4A 5F 8A F4 0C 92 26 5A 28 D8 BF
 58 A0 9F 8C BC 89 52 59 88 6C F8 6E BE AD 66 9D
 54 2C 16 0F 0C CD B5 40 5B BE A6 38 4E AF 7C 95
 82 E6 81 55 29 41 44 70 34 EA 97 66 A9 0B 2A 51
 7B CE 5B 50 E4 54 4A F2 40 56 CF 96 8F 95 80 31
 F0 82 04 80 71 3F 72 07 B1 10 39 2A 84 72 F8 58
 07 46 F0 AA 5C 9B CE 20 BF B1 B2 D9 20 00 27 34
 80 7E 15 82 8E 51 E9 51 E1 03 4B 86 B6 6A 03 A1
 61 E8 0F 10 C3 5D 38 70 54 9A 4D DB E7 EB 33 F6
 72 53 7B 78 2B 57 37 3D D1 AE C5 1D 4E B7 82 0A
 E4 2E AD 32 FE 33 4D 0B 40 46 62 6F 47 E0 53 E9
 80 84 E7 A9 CD E5 79 24 5D D4 52 6D B7 18 E9 14
 E1 D2 98 0B E1 FF CC 33 CF 69 CB 92 D9 50 EC B2
 5D 67 50 16 01 A2 44 3C 1C 93 14 64 37 12 A7 C3
 46 F9 91 60 95 03 07 E4 DE 51 0E A2 47 15 53 88
 B8 D0 11 0C 40 DB E0 58 C3 26 9A 5A D4 EA 35 5B
 71 D1 38 71 B1 F0 95 05 2B 79 42 FC 45 33 8A AC
 08 C1 DF 79 ED B0 D9 0A 79 3A A6 7B A9 16 05 73
 C1 58 8A 94 F3 FB 65 BC 92 2F 41 44 85 68 B3 42
 A8 59 3D AC 96 57 98 EE 5D D6 7D 18 06 93 7C B8
 3C A4 2C D0 8E 68 C8 DE 0D 56 8B 96 63 CC 78 AA
 35 51 21 29 5C B2 B1 3F 6D D2 7B C8 9C A5 1B AD
 7B F5 A8 DD 4A 0C E9 55 17 F2 F5 84 3D 8B A9 85
 56 5D 5B B3 4C D7 99 97 58 6C 61 16 2B A4 4A 03
 58 54 0C 4E 1F 50 71 00 A9 E7 1F DF B3 A0 7B D1
 0C 63 2F 8E 9C 34 A0 D3 72 DC 37 63 07 CD 2B 12
 20 54 1D 54 20 35 68 91 37 54 6C E9 E7 FC 1B 7E
 2B 31 02 80 B0 E5 30 36 24 45 FC AF 6A FA 71 4C
 70 C8 EA CB B3 36 AD FB E0 7D 55 1D 05 51 D1 6C
 8B F4 5C B4 60 C3 77 73 EF F6 0C 41 5C CD A2 F3
 B9 9A CD 40 23 A8 5A 02 F5 CE C5 BE DB 74 A8 7A
 D4 AC 42 73 B9 F1 E9 3A 98 EC DF E7 6E 72 A8 1D
 24 A1 CB 97 AD 4E 55 E4 57 AB 69 47 B2 3E 49 B2
 97 8F AF 54 BC 1F 24 39 F3 C2 25 EB 0E 1A CB 79
 54 63 32 59 72 94 1E CF 13 1B 6E 73 88 4F 37 A9
 73 B9 22 CD ED 11 0F D2 E1 6F B2 0A A9 27 52 B0
 AB 5C 6D C7 FC A7 A3 45 FF A9 A2 14 E8 2B 31 A2
 8B 3D 23 AD 46 BA 55 12 13 47 1D F8 2C DA EA DB
 34 5F 05 F9 05 FE DF 10 99 C0 6A 55 34 85 EC AF
 A9 96 9F 62 B1 6B 0B 74 F4 DC 26 FB C8 1B E8 43
 98 6F C5 8E B7 E8 25 CA EB 1D 67 17 4D 77 34 91
 21 D9 B9 2F 82 8A 44 FF 47 E8 BE 05 F8 1F 27 DF
 D7 25 93 AB 73 79 19 8A 05 F1 6D F1 81 8F 24 53
 7C 1A 98 8A AD DB 3D 5D 8A 22 3F 33 4C F8 BC 38
 EE 3C 11 CB 7A B7 EC 4C 84 D4 A1 B2 33 3B C2 BB
 52 E4 A9 13 D3 D2 8D 5B CB B6 D4 AE ED FD E6 74
 76 6F 68 46 25 97 9D E9 A1 86 66 3D F5 32 69 33
 A1 9F 67 D3 8E 6B B4 16 E5 99 77 C1 E1 D8 C6 D4
 B8 E8 B1 6D 10 BB F0 11 F8 1F B8 94 71 2E 0C 05
 11 F1 82 A0 8C FB 90 79 13 D1 16 5C 85 F9 AC C9
 33 59 46 F0 22 47 CB 0F FA 0A AF E1 86 D7 8B EC
 B8 24 F2 40 24 0C A2 9D B6 EF 65 EE 9C FE F5 9F
 1E 81 86 35 DA 5B 7E B3 77 EB 9E D5 D1 51 B3 69
 C0 3C AD 35 75 D2 0B D2 C5 20 EF 85 59 98 D8 E1
 A9 BB DC 77 6C AF CC D3 C1 B5 E7 34 96 FD 48 0A
 CE 2D CB F9 15 52 06 9A 5C 2B 21 69 D8 33 E5 EE
 5D DF 6C 36 18 65 3D 16 E0 0F D8 C8 69 B5 C2 25
 FD DA FE 7A A4 E5 86 28 25 CB CB 10 CC FB B9 F2
 1A D6 75 5A 95 3D 10 16 63 C7 B7 29 A7 3A 3B 85
 50 A5 16 5C 45 4F 07 32 BB 70 2F D7 9C 9C B1 20
 95 A4 B8 F4 EA 53 CB 0F 40 FA CB 8A AF 67 F8 44
 F8 3B CC 4D 7E D7 85 BD 0A 8F 12 96 54 20 7B 7B
 C7 7F EA 62 C1 22 DE C5 38 A1 AF DF 9A B9 FF 4E
 56 6E BB 53 C4 45 9E B9 44 D1 55 72 87 C6 1C 76
 89 3A 5A 74 1D 0D 65 61 34 2C BD 1E 43 11 78 51
 C6 32 B1 2D 9F 38 05 40 90 AF FF D9 66 0D E6 66
 17 95 C4 4C 8D 43 51 26 74 33 0B B5 18 D3 3F 33
 94 30 54 EC 9B 3B 53 8B 1F 4D D8 08 17 21 97 DF
 78 67 23 FA 7C 96 E1 D8 9F 0F 80 FA D5 64 EA 3E
 F0 C1 81 7D CA 06 49 23 D5 4D F4 C5 51 66 D4 74
 5B B6 6A CA 54 8F 9D 73 4C E5 8F 28 6B 51 0A 20
 53 DA C4 B5 E3 B1 B9 DE AA 9F DD 3E 3D 40 04 E9
 6F 8B 89 47 6F 77 36 27 F6 95 B3 5C 27 25 BA 7E
 42 8B 2A EC 37 F7 FD 34 B3 14 E8 64 C0 1F 23 1C
 81 A7 CE DA E7 CA 3F D8 6A 89 90 61 E2 C7 37 97
 B6 7E 3B C3 CC D8 8D 02 B5 E0 7F 79 D0 FB 9E BD
 81 C1 22 24 4F 23 52 95 21 E9 CC 6A 82 B7 E0 91
 E2 73 AD C0 3B F7 64 68 21 EC 2B B2 B6 72 EF 6E
 2A 81 F8 B0 60 64 BA 83 E3 21 F6 C3 99 4A 94 CE
 BA 9F 88 5F 84 38 F1 B9 74 09 2F 70 4B E8 04 E8
 41 18 E5 4D A7 F3 18 4E 1E 26 F0 FB B5 42 B4 84
 09 8E 09 D8 01 F7 5B 7D E7 43 73 0C 26 38 EC 42
 DE 07 70 E8 D3 C9 00 8E B1 BD 47 38 00 24 B8 0D
 41 02 95 43 73 00 4D 83 5B 42 49 DF 2A D2 3D EF
 54 D2 F8 97 9C 94 D9 A4 F6 11 7B 52 FB EB 35 2B
 29 2B 68 97 51 F5 6B D4 78 77 B3 D9 99 6C 1F AF
 BF AD 11 C0 8D 05 E3 25 19 BD DD ED 72 90 EF CA
 8A 94 BF C4 DF 8E DB D3 1E 65 47 D0 BC 91 A8 BB
 DE FE 17 53 CC D1 A5 AA 32 C7 97 3F A3 E2 15 38
 09 18 E3 5B 0F 66 2D D9 4D B4 A5 6C 9E 37 9C 50
 A2 64 D2 D2 77 E3 9A 3E 53 B4 C1 BF 47 79 EA 7A
 4C 5F 69 A9 D8 87 5E EE F2 A2 D6 26 0F 9B 8D DC
 49 C8 8A C5 CF 1C 4B E8 3B DF C1 A1 37 FD 33 A6
 1E 27 6A E3 77 82 92 05 A4 08 02 BF F0 AF A7 7C
 0A 8B CC E4 EF C8 CF 4C 47 C2 5A 00 84 66 8B 7C
 5B C4 CD 0F F9 9D 00 74 23 EE 88 05 7D 6C 3C 67
 B9 18 38 E4 69 14 D2 1C 58 13 EA B4 0F F1 79 85
 96 F1 D9 44 3A C0 FB 20 31 27 5B 0F AC C5 E1 19
 DF E2 4E 0E 7D 38 7D 9A E8 2F 2F 98 9C 4B 60 2B
 BB 78 93 D7 E5 36 D0 C7 4A 14 0A 8E 6E C8 E4 1E
 F1 C6 3C 57 4E 96 4F 78 BC 52 CC BB 0F D2 43 10
 21 50 91 C0 AE 56 F3 47 0D 81 B8 8D 41 11 6D 2C
 19 7F 39 F8 5E 2B 7B AA 30 3A 5B B8 A3 51 0E 72
 42 07 76 09 40 95 96 74 09 1F 15 CE 10 F6 1F 25
 5F 76 F7 AB A2 30 96 B8 13 E7 2C F4 C9 31 CD AC
 4F 0E 0D 10 09 22 72 9F 50 11 22 5F A3 6C 9D CC
 6E BD 7E A6 35 71 C4 7B 88 AF BC 51 59 42 6E 37
 25 3B 3B D8 4D F9 A1 91 5C 47 C3 00 9D 09 3A 79
 B8 82 77 4D 06 A3 3F DD A8 6E 6C 29 EC 7E 99 99
 63 F7 F3 17 76 EA D9 F8 7F C2 05 5E 32 8A A6 C0
 E6 C0 82 0D 58 77 C7 DA 98 1F 0A 3B DC FB 85 17
 64 03 1F E7 78 BE 3D EA 63 3F 9F 3E 73 22 45 C2
 C0 2C 99 10 0B 21 1C E5 DA 10 EB 32 F5 83 DA 3C
 23 58 C2 3C B3 41 74 C1 28 25 54 2C D6 49 05 54
 ED 58 BB 18 2E 8D FC 20 CA 5E 91 FE 43 74 7A 24
 E2 CC 71 1B 1B D2 51 B5 C0 38 BC CC 13 D9 7C 92
 B3 3A FA 85 84 35 76 14 DF D6 6E 42 0A 2C F6 A0
 DB 5A A8 7F BD CA 0E D8 47 32 FD 4B 40 33 9D BE
 47 5F 88 42 26 E9 CB B4 A2 12 59 E0 9E D8 60 B7
 DC 9F B0 C7 5A CE 9D E5 26 9C 66 60 80 EA 7E 95
 5F CC 8C CF 06 97 09 F4 C1 F2 F2 88 C3 94 0E 47
 F1 D9 27 B6 A5 DA 52 63 CE AE 5D BB EB 40 00 F9
 BB 26 08 C0 A0 F5 18 13 94 EF BE 5B 74 DC 93 97
 F8 98 35 E1 5E 85 EC 61 EC 8B E1 34 1B 49 EE B8
 F7 63 96 AD CB 8D 9B 16 5D 83 17 32 36 CF C2 DA
 A8 A1 50 73 6D B1 9B 26 0E CD AE D0 31 BA 05 34
 F0 1A 61 11 88 93 D1 B4 36 8C 40 DC 60 03 AC 8E
 07 9F 6B 53 9B E1 AF ED 9F 26 ED 60 5F D9 52 32
 EC E0 D6 C0 C4 5F EA FD C4 D7 E2 F3 86 23 E8 01
 B5 1D 77 16 8E 88 C9 77 0F AA BE 0F 88 53 6A 8B
 3B 3F CC 37 57 07 F1 85 13 0B CE BB 09 41 1A DE
 BA 05 A7 66 64 62 CD 1F E2 E3 5F 0B 4A DC BD 43
 84 E0 4F 29 86 00 12 28 A8 A0 26 BF 8C 58 1C 86
 81 8A 47 8C 40 92 39 7B B7 DD AA D2 45 DB 0C 50
 B7 28 58 3A D1 46 93 9E 93 53 F4 1D DC 3C B5 83
 FA E5 C7 06 0B 34 26 3D 3A B5 BB 0D 9B 67 FF EF
 F0 B5 7B CC E5 43 BE 70 CF BB 57 73 A6 F7 80 5B
 AF 3D 0D 72 98 1A A0 EE BF FC 99 17 6F E2 2D FF
 E4 3A D8 D7 1A 2F 2D 18 4D DE E3 FC 39 28 B7 37
 E9 44 38 0F 68 FB A1 76 DA 15 BB CE 63 F5 E8 BB
 62 6A 32 7B 6A FE 0D EC BB 90 D8 C4 AE E9 F6 A3
 58 70 A2 30 18 B6 D8 38 43 08 97 5F 9F 1F F3 3A
 DB FC 8E 2A CB 43 13 33 78 61 72 6E 3D 7B F1 B0
 78 78 A2 E3 EB 70 E6 AC F9 24 4A A7 D6 CF 61 8D
 79 BF BB F9 49 70 AB E2 7D BE 0C 13 74 8C C9 F4
 1D 26 8D 59 E7 48 9E 17 78 16 29 4E 1F 8A 78 9A
 B7 46 BC 72 26 60 01 E8 DC 4E E6 3B 6B DF 4D 8F
 25 1F 15 5A 11 8A C8 B4 39 9A 37 28 A8 11 06 E2
 19 44 75 F0 A2 67 1C DA DC 58 BF 18 8C AA 1A B9
 C5 62 69 54 33 9E 23 8A 82 AB 28 19 1F BC 34 9C
 A2 7B 87 30 35 CB 48 A2 57 E8 23 09 2B 57 C6 06
 C9 9B 4F 1C 82 E5 CC 9F 6E D4 E0 F0 DA E2 0C 19
 90 F0 43 FB 08 11 54 FD 8B 73 98 CE D8 27 82 DE
 69 0B B8 A6 61 63 CF 39 9E 23 D8 5B 36 CD 39 F6
 1D 23 78 88 9B 6A 36 EF 8E AD 6C AB 49 A8 4E 45
 4B 22 17 9F 76 E9 A6 90 F0 A1 7B A1 16 99 C7 51
 B8 49 7F E6 DF 59 E3 64 8D B8 37 E4 54 91 30 8D
 FD 22 76 32 00 71 59 E7 32 A0 62 09 52 EF 3A 0F
 CD E6 3D 84 8C E9 21 38 BD D8 6C 19 4B AD B8 89
 0C B2 CB 5B 1C 3E A8 F1 76 08 F3 73 13 BC C9 9C
 76 20 9F 50 6F 14 A7 9C 41 FE 18 02 A0 FB DB B0
 EA 48 47 11 4D 92 13 80 E2 2A 57 B5 62 FA A0 75
 D5 E8 80 4E BA F0 A9 91 FD 39 BE D2 0A EC 67 09
 6D 3B E5 74 C8 42 9E F1 54 72 7D 23 A2 91 4E 85
 1B 15 88 62 EB 77 65 BA 8D EE 10 E3 1A 39 57 D8
 3D 86 03 CF 23 3A 16 25 EC C4 57 58 C8 65 E3 72
 55 C7 68 13 77 4E C1 C0 AF 58 8E D0 2C B1 52 05
 5E 46 A1 14 7D 6C B4 B8 07 A1 78 4C 83 72 04 E7
 7A 35 B2 83 F9 5A EC 28 38 A0 20 B9 36 57 5E 1E
 D0 98 05 AF A9 2E AD 36 0F 8E 5E 76 52 F4 0C 5E
 84 45 84 40 C0 3C EB 33 64 B1 18 0A 87 9B 43 BA
 96 C3 54 22 BA F8 D7 76 0E BC 24 37 0C B2 52 39
 B1 A5 B3 E5 D5 32 9D 90 6B 95 36 DA F8 63 9D 1E
 3B F7 C2 C5 0A 5A 3A E2 8B 1F 54 B4 29 56 76 3E
 23 19 72 81 CA AC E6 EE AD 41 F2 ED E6 2B 46 E7
 9A 9C F4 A8 BD F0 4E 9B 29 EA 09 14 CE 8F 05 05
 E5 51 BD A3 85 CC 6E 41 A4 4F D9 F7 72 F0 EF 90
 72 4B 23 B1 CD 12 57 72 42 8C 6F 44 7C 78 B3 B9
 44 84 23 56 BF B6 0C 1A CD 7F AA A1 EE 26 A8 E1
 C6 E8 78 23 E8 F2 2E 76 2E C2 E8 3B 14 3A 0D 5B
 F1 34 AC 00 03 27 71 DA 6A 2A C3 51 DF F5 AE B4
 47 EF 2B A6 E0 3E 29 36 4C D2 E0 6E 27 64 56 9F
 A2 8F C2 2D 9E F7 EE BC CF 40 E2 A2 69 6C 45 39
 56 C5 25 F3 2A 84 92 D8 1D 91 F7 AA 5E 6D 17 FF
 48 39 8B 73 F0 2D 8F 97 38 94 91 4F BB 95 7F 5F
 41 05 EC DF 16 36 BA 21 B9 02 AD 41 26 D7 F6 57
 40 2D 76 B9 CF 55 59 A9 C9 A0 B1 BE 42 F3 50 FA
 4E B1 60 39 54 60 25 14 7B 8F 9D 35 BA 30 AD 5F
 D2 70 E4 47 26 69 35 7E 1E 67 66 DA 40 E2 24 CD
 31 67 59 AD 5C 41 5B B7 F7 81 C7 5D 1C 5B 52 41
 4D F3 DC 01 F9 41 8A DC 9C 7B 3A F2 EC 4F A3 5F
 E9 B9 C6 E1 C7 8A D6 B6 51 B0 5F C7 CA BB 61 88
 64 F0 FC 3F AD EA 0E AB DF 14 C0 FF 78 37 41 B7
 C6 44 6F 9F 47 E7 39 4E E0 ED 8A 7E F1 A7 F5 F3
 43 BA 4A 94 28 9E 48 3E 04 23 0E 14 25 DB A0 BF
 35 70 6B C1 47 52 1F 0D 1B C4 9D A4 A1 FD E1 50
 EE F3 EC 04 F2 9C 0B E6 F2 68 7C F5 A5 F6 0C 92
 16 6C 8F 8A 69 E7 60 50 90 31 0C A7 28 BE EA 69
 20 79 26 45 E7 58 44 A6 2F 92 EF CF DA 73 06 12
 B3 AE 59 0F FB 12 B0 6A 29 52 25 8E 11 CC 14 B2
 B8 2A FD DD D2 6F 0D D0 D7 07 58 9E 04 D3 1F 4D
 55 0B 70 66 5D A4 8C D2 2E 60 55 8F 42 7A 6B 67
 8B F3 59 D2 A0 BC 3B 51 3A F8 0E 5D 06 FA E3 51
 A4 A3 1A F8 56 BA E3 F0 79 E1 10 13 20 E4 AF 9F
 53 DA 96 F5 AE AF DB 52 26 C5 59 CD FC 13 81 87
 A2 18 89 1A 9C 4C D8 63 29 E5 A2 D4 D7 45 88 35
 0E 7C 28 EF D3 3E D2 D0 94 37 2A CD 2F E8 17 A5
 A3 43 5B 3F F6 E8 85 32 B4 54 F6 D1 18 8C 60 7B
 72 48 08 C9 26 B7 9D 4B B8 F2 50 4F A9 A7 5E C7
 E1 34 A3 B2 07 D9 63 73 1F F5 9F A1 54 B4 4F 51
 BB 01 BE C7 ED CF 5B 38 BD 7D 86 C1 5D C9 2F 6B
 1B 8A 91 F1 3A A5 6E 29 8C 1D A6 05 9E FC C9 C6
 E7 0A D0 89 6B A1 FB 2C 13 2F EE 0B 49 C1 98 23
 C5 B7 85 08 88 7E 44 AB DD B1 54 AC DC 19 3E DD
 B0 8B 15 19 AD FF FE CC 9E 4A 97 EA CA 13 39 7E
 1A 1C 37 FC 7E BE 94 68 08 0B 9C 74 C4 8C 21 73
 E3 08 60 2F 28 7B DF C2 74 4C F4 35 6B CC 43 8A
 2D BB 8D 4E 1B 15 D7 37 33 5F CC A8 D8 02 B9 CC
 8E 14 A2 22 76 F4 DD 38 52 40 33 45 34 47 4E 04
 34 EA F5 75 00 A1 C6 58 6F CB 30 CA C6 BA CA B8
 C5 17 AC A6 56 DA AF 37 46 25 A4 7F 4C 26 E8 97
 15 C6 0F 5D A9 0B 92 2A 7D 4C 49 D7 E0 9D 4F 95
 B9 E8 3E 80 78 D2 FF C6 FB 73 F1 AF AE B1 7B D0
 8E 1E 5C 88 BC D0 B1 A5 00 93 72 AA 07 CD 9F BD
 EC 04 9E 2F 9F 76 FF E0 B2 43 FA DE BC 9A 7A 0E
 F3 21 96 A2 8C FB 9E AD 38 BE 4A 4E 11 E7 8B A2
 A5 99 26 7E 30 27 A4 DF 8D 3B E6 9F 80 D9 0B E4
 66 56 00 26 57 F7 C2 B0 B1 34 AA BB 9A 7A 0D 7D
 D2 DC A8 35 D6 B2 B6 2C E7 5C 70 3C 7E 55 5F 6B
 0F 7F B4 19 40 F7 BC C2 BD 30 D2 35 85 01 E1 2D
 15 A4 B9 48 37 81 8B 58 F1 03 77 82 60 08 D1 22
 07 AF 7F 3A 1C DA 10 ED 3F 35 C3 E7 75 05 A6 A8
 C3 1E FB B2 9F 9E 81 67 1A CC 39 01 C0 22 EF 9F
 57 9D 77 31 D5 A8 52 9E A2 C0 8E BD 29 59 F8 94
 90 BF C9 4F 12 CC 0F F9 37 6D F6 BB A2 BD 6A B9
 A4 F4 91 0D E5 4A EF FD E5 AC 9D 5E 00 67 18 1F
 92 9E 87 4B 74 18 52 40 D5 C9 B2 F6 D4 4A 0A 51
 FA 05 9A 14 80 E4 BF 17 46 1F 2A 97 A8 2F 31 AB
 4A B0 D3 DA 14 B5 69 9E FE 29 7B 36 DF 16 D1 14
 F8 55 94 00 F0 8D B7 44 51 47 38 90 67 67 DE E7
 B8 F6 C5 04 0A 84 80 34 E2 67 BD 60 4B F3 50 39
 4A EA C5 C6 CF 8D 85 77 D6 0E E5 42 61 13 D0 7E
 84 54 28 2F 9F 76 C5 EF EA CA C9 5C 2E F8 3C D0
 29 46 25 3F E1 BC 2F 58 21 47 C0 36 D6 28 53 9A
 15 A2 AF 83 60 B1 A3 B1 C8 51 54 C8 ED F5 98 B9
 D6 BB FA 42 38 59 3E 46 1D 1E A3 F4 09 C9 A4 BD
 54 02 B2 30 65 E9 B5 2E 85 33 1C 1E 1B D9 A8 88
 B6 D1 FB F3 68 64 23 CA A6 C4 1C 73 E3 BE BE BE
 4D 49 C4 65 03 60 0C BE 94 FD 45 B7 10 D3 4E 87
 7C 30 C0 64 6D 5D CD B3 7E EB 58 A7 15 E8 96 6F
 1C 6F 7D F5 6A E9 8B BB ED A6 CF 0C 20 CA 4C 10
 0B D8 C4 15 70 EC FE 38 59 54 8C EA C3 1E AF 89
 E5 B2 AA F6 15 CB 8E 00 05 14 4C B1 19 7E CC 24
 F6 53 1C 31 1E B0 3B 72 7D FE 08 BF DC 65 D6 A0
 86 8A 36 8A 2F 89 CE 86 89 BE 34 BC 31 A2 82 DE
 8F E5 0F 75 69 04 16 11 11 64 58 51 74 E8 70 7B
 57 29 54 87 37 CD 41 F4 B1 90 A4 6C BE 7A 0F C5
 68 8D 61 0D 7F AC 0F 3C 4D A6 77 85 78 57 24 6B
 26 FE 39 AF 24 00 B4 10 4E 0B 99 B3 F1 CD 2F 3E
 77 98 F1 42 74 3E 78 12 48 9C 52 64 D6 F0 8D 81
 EF 28 4D 96 AC 85 DE FC 16 6D 45 46 0F 25 70 30
 7B EB F0 90 D3 1F 92 2A 10 5D 93 85 76 E1 FE 0B
 8F C8 89 16 22 1A E0 FD 8D 6D 9D 3A CE F6 70 FE
 B0 8B F4 8F 1F 4F F6 F0 46 F9 6C 37 98 30 58 01
 55 26 A6 74 30 B2 E7 E0 85 72 69 D7 D4 FC 11 A9
 71 79 09 ED 45 FF 1D 2C 8B 44 C0 5E 7F 83 84 21
 8B 58 C4 4B A5 65 89 F9 E8 DE 2A 63 6F E6 3C 1E
 95 36 C5 ED B9 43 BF 7C 1D 0E 7B 55 72 C1 36 A9
 9D F9 50 DD E0 2F 1B FC 2B 60 67 32 59 9E 6C C2
 7E 71 00 80 DA 90 3D 28 7A A9 7F DD 40 43 28 78
 0B 09 E3 FA 43 40 75 67 3A 90 F4 2E 81 3E 0D A0
 A2 0C 87 DC 37 EF 8D 5B 1F 88 28 EE 50 5E CC E1
 FC D1 FF 97 C0 9B 8C C9 C3 97 11 21 7C 6C 7B 2D
 9F 3E 60 0B 4C 17 84 6A 53 78 71 41 0A D8 C6 22
 CE 4D 3A C0 16 3B 55 3A F0 44 6B A4 AC 47 D6 8E
 70 41 2A 5B 8B 87 64 1E 9D CB 9F 3A F7 CE 5E D3
 0A 35 B8 BE EA 48 3C 2D E5 A8 35 8B AB 32 FB A3
 48 43 A9 64 3F 05 AE A6 24 36 15 93 67 37 2B B0
 3C 19 0B DF E3 0D 78 39 64 B9 C4 F8 8C 33 51 60
 32 25 FB B3 F0 41 7E C1 4F BE F9 34 E3 08 7C AD
 57 86 CD 6B 45 58 9B 6E B8 74 69 E2 9F 23 47 D6
 A2 96 22 BE 15 33 DD 02 7C 93 DC 60 FD 04 FF 6E
 ED 51 C0 9D 6D 8E FA B0 B6 75 75 92 6E CB E5 F0
 2E 6E 74 23 9F FF 31 A9 2C 6B B5 F0 27 25 AC 15
 16 4B 3E F6 BB 0D 36 B4 54 99 2E FC 61 A9 78 41
 A8 DF D2 4D 3C 5F 47 B2 E8 35 E4 E6 88 AB A6 E8
 4D 7C FB 7A 5F 59 C2 5B 4A C5 E0 1D F4 DC 78 E2
 54 06 C1 62 F5 F0 E0 42 6E 6D 43 3C BF 21 78 4A
 B1 91 09 BF FE 1D 28 F0 74 2A 62 F9 72 79 0A 39
 A8 CA C0 E3 FD F3 94 BA C4 DD 96 7C 43 41 37 D8
 F9 F1 DC 84 A3 79 76 BA 11 C0 A8 31 8A 03 5D C3
 03 8A 1B D5 E8 CA 01 E3 7E 92 12 61 19 46 20 BF
 7B 77 89 30 93 6D 1A BA 28 4C B0 1B AE 2B C4 33
 92 DA 78 FA D4 02 EF 4A A4 E2 D6 07 C7 E8 6C D5
 56 F8 3B 56 DF 52 0C 55 9E 8A B3 7D 42 66 E5 7E
 63 F4 55 A8 96 58 CC 69 10 D6 8A 9C D9 3C D9 67
 77 63 43 A5 05 64 AB C1 B0 B4 B1 5D 42 DB 40 26
 56 1A 69 15 C8 D4 A3 69 80 38 C9 E8 79 85 45 19
 79 35 54 B9 46 98 E2 83 A1 92 75 1F 3D E7 3A 18
 8B F3 E2 75 BB 69 03 E8 69 6F 9B 7C 76 CD 6D 95
 40 9C 31 C2 84 AB 9B 4A BE 14 66 21 DF 95 91 84
 D9 85 39 0D 08 A7 8F DA 40 7B E6 B8 65 1B 86 04
 5F EF 96 20 09 A0 62 6A F8 AF 68 19 6D 47 B9 8B
 13 27 DF D8 73 20 27 C0 0E C6 F2 B0 C4 30 77 5F
 58 70 F3 E5 D9 96 90 DD DB 14 C1 11 F0 9F 59 CB
 7D 6F 91 EB C4 80 59 AA AA 7C 50 D4 1C 9F 74 FE
 44 F4 9E 34 99 8B 7F E8 26 A0 CA 80 18 CC 52 A1
 18 A8 1C A6 94 BC 3D C8 24 58 5C 75 AD CE 6D EB
 C9 66 ED AA 9E FD F8 4D 9A 76 3D 1F 71 26 22 DE
 F8 44 91 23 2E 5F FB FE 76 2F 71 75 52 76 0A A0
 AF AD 11 8E 30 6E FD 2F FC 66 2B 57 12 F5 CD D2
 44 81 F6 6C 70 4A 50 14 57 87 E7 26 31 1F 54 03
 1E 54 E9 8B 3F 4F 8C 58 D5 68 AE 62 35 64 80 53
 2D 00 74 68 21 43 28 FE EF DB 4E 33 2D F8 F9 F6
 FB 6C DC CB CC 53 F4 93 C8 48 24 AC EE 52 44 99
 C2 11 B2 38 0F 41 E0 08 3E 1F 79 25 15 4B 46 4F
 22 79 35 53 B1 98 F6 AA D4 1F 72 93 89 02 17 6E
 FD C0 0B FA 8C DA 59 2A F8 64 C7 C5 0B 9B B9 45
 2F 86 F0 D8 D8 E3 95 51 3F 1E A7 1C 25 6A 0A 14
 AB B6 12 DF B2 1F 41 5F 5A CC 38 BC F8 E6 9F FD
 9F B5 37 D7 A5 0A E8 9E 4B E9 87 CF 8F CF 15 BE
 A9 29 E9 C4 79 13 9E DA 04 A4 EA DB 68 BD 23 A2
 8A EA CB EC 52 BD F1 6B 87 0B 6E 98 00 2C 88 3D
 11 7D EE 95 25 44 46 64 45 51 C7 9D 84 AD D8 39
 B3 69 65 BE 81 76 F5 90 E8 53 D2 BA 73 5A DE 30
 25 4F 20 A4 7C 7B 36 74 EE 54 A1 CF FC BE 87 04
 69 77 CC FF 7E 3A 0D 7F FC 61 12 BA 3B 6A BE AD
 7F 4B B0 54 68 AD 5D 30 12 16 74 9A 27 3A 3E C0
 D6 86 B5 52 A5 E4 56 E1 DA 1F BE D4 0F AF DB 82
 76 F7 7C 41 CF 16 0C AD DD C5 0B 9F 9C 70 ED F5
 E8 FE CC 0A EA E2 55 5D 31 40 5E 3D 68 9A 11 6B
 FA 93 C3 1D 5D 77 98 AE 8A D7 63 78 BF 55 2F 41
 92 89 8A 6B 0D 91 3E AD 75 1F DC 30 D5 CC D9 FE
 97 DB 71 40 86 4C AD 26 98 88 74 EB 9F A4 5B 45
 91 82 27 4C 50 04 EE A6 48 07 06 57 F7 B8 FF FD
 A6 62 A6 B4 F3 9E D1 3A 7B 09 D7 CE 9A 02 3B A7
 AE DF 55 D7 A4 93 99 A4 77 8A E5 81 3A 9E 25 6E
 69 4C 08 E5 48 94 D2 0D B9 EA DE C4 13 2B E3 6D
 2B FE 11 51 5F 00 75 F8 A0 B8 F4 62 02 4E 30 D2
 A3 77 49 5C D1 FA D4 D8 56 17 45 DC 6A 9C 7E B9
 D8 5F F2 7B 98 BC ED F6 FD E8 9D 40 45 80 96 B0
 CE C0 74 01 10 E5 A3 80 03 3C A0 30 B7 FB DD D5
 D4 F4 46 C4 30 E6 EE 0D DF DD 55 8D 8E E8 75 20
 73 1F 4D BB 5B 5D E8 D1 2F E9 DC 48 4C EC 2B 2D
 A6 C2 4C E1 5B 77 83 59 3B 9D F9 59 F2 F7 7C 66
 C6 0F 5A 16 90 B5 76 C0 32 EB 4D 99 8D 3A E3 E5
 DE E4 4E 12 4B 89 42 9C 46 CB DB 30 A7 5B 7C 1A
 C6 D4 0C 50 02 83 39 EB 3D 0F 88 4C 22 3E 59 60
 A0 B9 08 CA 07 36 1D A4 8D 86 ED F9 21 05 DD 43
 9F 97 06 63 0D A2 95 72 02 8C 62 4E 7D DB C9 45
 C0 99 37 AB 8D 89 74 DE 47 35 C2 9B 24 53 69 2C
 07 09 91 A7 B9 6C FC 0A 1F AB AB 90 78 4F 65 12
 18 B2 40 4C 63 52 53 37 5D A0 3A 94 4F F0 AF 8E
 13 75 0B F1 10 32 38 F5 05 B7 92 FE 29 D9 5C 77
 84 49 0E 0C F6 86 FD 30 C8 74 50 02 DA EA 2F 1F
 81 0B 77 13 E7 7B EA B3 AA 94 40 3A DD E3 15 73
 1B E6 19 8E AA 64 30 8C 78 FE B5 36 AC 51 68 E3
 7B 1C 58 E8 6E 4E 71 E2 75 6B 66 65 E0 E9 F5 58
 D2 B6 90 6C 8A AD 4B 21 6C 56 8A D3 59 AF 2F FA
 CA 91 99 16 1E A1 28 3A BE 5D 8F 64 23 CA 44 6B
 3C 1B 2A F1 67 E2 9F B5 F5 6E 5E 13 B4 AF 9C 99
 D3 32 72 4E 43 DD BE 75 BC 6D FB 34 C1 FE F4 CC
 07 85 40 F0 C3 B9 FE 3C C4 1A 82 AF AA BE 95 61
 59 93 2A CC E8 22 C5 3B 4B A0 D3 89 34 C8 F9 39
 4C 85 7C C0 84 CA 87 83 CC 06 39 E9 06 69 E3 09
 9F 3C 60 DB 62 98 3E C1 5C 24 43 2E D9 89 6B 5C
 2E 41 29 1B 8B 1F E5 F6 F0 5F E9 38 73 A4 54 6F
 8B DC 05 DE 4C 16 B1 3B A1 11 E2 94 AE 6D D1 31
 AE 92 40 61 A0 A4 86 48 F4 F0 4F 70 AC 08 46 BC
 77 EE 44 5E 4E B2 23 05 08 BF 00 AE 21 4C 28 1C
 F7 7E 4D ED 6B C0 95 7A 26 1F 2A BE 2B C4 D1 9A
 69 C0 1F C9 FA 35 FD C7 78 A8 CC DE CA 2A 3E 10
 27 BF DA BE 37 EB CA 03 B3 CE D2 19 0D 6D 9A E8
 78 35 2D 48 F7 B7 B8 CB 4F DA 76 66 4E 02 D0 9D
 90 CA AA 06 D4 81 B9 13 4B E8 B9 68 C8 62 95 F4
 45 A7 67 99 4E 08 32 53 E5 F8 7D 52 D2 B3 65 ED
 44 C9 26 4B 62 92 36 8D 8C 84 38 AD A1 1E 27 04
 B6 9C E1 11 1A 08 6F F1 57 7A 33 AB 77 E0 CD 48
 2A F0 A6 E7 00 F4 C8 67 4B C6 13 09 7E 71 02 31
 B8 0A CC 6F E4 44 75 49 0F F3 96 C8 71 94 AF FD
 24 15 BD 8C 62 4F 05 C2 7D 05 A3 CF A1 27 62 22
 96 A6 75 18 86 E4 C1 8B 2B CC C9 53 EC 9B FD E9
 8C 10 CA 52 D1 F4 B6 44 67 1F 13 E0 AD B4 3A 45
 90 BE 8B 2A 1A C5 B5 E3 A1 34 C2 E8 57 05 42 2C
 62 DC 1A CD 51 90 01 44 F2 E8 F7 14 BD 4B 59 66
 2E 06 F2 99 11 66 B1 74 7C 8D 68 BA CA 28 2A 43
 11 37 66 50 B7 ED 1D E7 B8 05 55 47 B5 7F 21 98
 61 60 76 24 9C AD D7 C3 2A 41 C6 6D 88 34 AC 80
 ED CF 01 21 FD 29 BA 96 F8 71 9C 87 AF 36 9D 1D
 97 F8 C8 C9 EF C7 18 EB 52 D5 3A 53 7A 11 91 E2
 6A 18 02 EE 57 DD FA 61 DD 35 A5 04 69 78 18 2E
 20 90 EF ED 6E B1 5F CF 74 C1 FE 8D 76 64 B7 2D
 C4 20 67 9B B3 57 6D 88 74 6D 59 E4 73 1A 83 40
 4D 87 ED 46 51 78 AA FE 67 30 FF 70 57 A6 B9 E1
 AA 0E 22 DE D0 86 BB 6B 02 4B 2C A4 49 69 C3 30
 AB 7B 55 91 8D 57 DC 84 A1 B4 8E B3 71 62 E8 DA
 E0 91 40 83 23 8A 06 13 52 4A 74 CD 65 F3 81 7E
 76 15 92 27 BA CE C3 DB D0 19 11 1B E0 EE 18 21
 4F 43 62 F7 4B DD 88 E0 2A 2D 47 01 DE BB E4 67
 3A BB 94 2C 28 10 C5 1A 6B 9A C2 FB EF E8 C5 D7
 37 0C 13 98 13 1D 92 49 F6 C7 65 A5 C4 25 64 EF
 88 1E 71 0F 7C 50 C3 38 48 AF 9F 47 54 06 9D DA
 17 BE 3C 9E 44 E7 4A DA 0A 51 4D 8F E7 8B 74 70
 66 F5 5F D5 F6 D3 A3 8B FD 95 6F CA 60 BD 3B CE
 F4 E2 59 84 B3 8E 16 20 77 A9 1D 5A 70 63 FD AF
 78 0E 87 CE AB 26 40 1E E3 95 97 F9 E2 4C 18 63
 4E ED A9 44 B4 EC 30 1F 3D 17 75 15 78 76 75 93
 98 42 E7 AB 8D 80 53 8E 94 75 35 D7 FB AD 4C E0
 D4 63 AA DE 9F 9A F1 D7 7D E0 72 D9 1F B5 16 39
 C5 89 69 98 EF 9F 82 4B 36 09 F0 C8 CA FE 64 66
 0C DE EE 3F 72 CE 15 92 CB A0 7A 1C 4B A6 74 FA
 29 92 11 50 1A 57 9C FB 95 AD 01 99 0F 94 B2 C5
 4F A8 7D 36 DA 2F 77 2B A8 7D ED 5A 8D 66 1D BF
 6F 00 A8 F9 CB C0 2D 0A 5F B9 24 32 30 D9 8E 43
 48 0A 12 E6 55 5B C5 90 E0 B7 7B 45 E5 D0 48 08
 3F D2 CD 91 61 F9 98 5A B9 AE E0 27 2E B9 66 70
 0F 90 0C 65 0A 3B F1 C6 FC 38 88 FF 5C 9E C8 61
 F5 8B A9 11 35 05 D2 37 32 6B 47 34 A6 F8 5D 68
 C0 91 64 80 26 9D 82 55 1C A2 B1 86 EE 8C F1 D5
 BB C9 66 DE 8F 3D AE 11 1D EC 49 94 BF C6 84 86
 E7 61 1D 32 B4 5E EA 51 1A CA 65 52 6E A3 59 19
 33 14 EA 59 A8 6A 27 18 C4 62 58 43 74 39 FA E5
 05 0E FD D0 30 49 88 ED 1E 08 B9 65 34 52 CE 0C
 FB 9C A1 53 1C 3F EB 17 B0 48 89 A9 E1 C9 7E 2D
 65 1F 8E 83 E9 81 9F 06 85 8F 0D 37 23 05 E6 D9
 90 BF 8E 3B C3 1E 9E FB ED D7 AA 1B 91 A9 85 15
 8F 17 62 D0 23 EB 7F E0 2B 65 E5 DA E1 CB 38 B1
 FE 45 E4 24 39 D4 CC 58 14 DA 8C 7F 38 9D 72 52
 5D B7 ED D6 DE C9 6C 07 8F 8B AC 82 96 51 31 D7
 3D 00 B4 84 59 E1 65 B5 99 50 31 F1 50 4E CC 05
 89 84 DE A5 46 1D 22 E4 8C E3 7F 4B D9 B1 08 6E
 73 AD 87 EE 03 0E AC C1 7B 50 5E 67 54 BA BF 9C
 8D B5 02 FB E3 62 B2 71 FB 33 34 D0 F3 3E C3 5B
 3D 80 40 51 44 87 16 B2 30 DD A1 A7 4D 65 F1 40
 C6 27 33 47 92 0A A0 DB 01 1E D6 EE 64 27 E6 6E
 3E 65 3A 64 F2 99 94 9A 4A 59 77 C0 7F 6D EE 68
 79 9C 12 44 9F 8A E1 85 0B 74 59 0B D1 7B C9 9E
 77 2D 04 EB 0D C6 C7 36 2E FF 08 CF 6A FF 92 C8
 9F 54 7D 42 41 65 84 87 26 38 86 60 16 B4 19 21
 9F 8D 22 36 72 F3 4B 9D 94 EF 0A 96 4D B7 6C 02
 73 8B 2E B1 A4 08 4A A7 A6 FF F1 FD 23 55 72 BB
 F2 B0 B0 07 56 58 DE 7B 01 C8 BF 75 37 75 A4 A8
 71 77 76 2F 5A 8D CC 0B F8 A1 F9 EA 9E EE 42 4B
 BD 49 72 5B CC 69 51 B6 85 E7 06 CF 83 D7 85 09
 3D 2B 60 28 D0 6C 4C 0D 64 75 5C 1E 33 A1 69 37
 38 AF ED 30 1B A9 ED F7 68 E1 43 7E 42 F9 80 F6
 26 26 7A D8 F3 A4 AD 36 3F 10 FB 27 15 2D 61 B5
 49 A9 89 38 43 1B A1 28 2C 23 EF C5 A3 10 47 FF
 4E 3F C4 70 57 6A 6A 32 3B 26 6F CE 31 52 14 64
 32 72 67 C2 39 74 AB 47 80 7A A8 93 DC 40 17 AB
 30 17 81 39 3B 03 29 30 5B 1C 67 62 39 1E 35 F6
 74 CC AD 03 5E 2F 0A 65 EB 7B CE EA 01 72 4A 7E
 A1 26 CF F0 03 3F 43 1A 19 5E 5D 84 A6 A1 06 E3
 B2 B7 93 C5 0D BD 62 5F 5F E0 F4 53 98 E7 C1 B3
 7A 0A E3 C6 26 DE AE 45 D4 AA 23 98 9E FA 29 00
 91 FE 33 5C B1 14 C8 13 CD 60 01 9C DB F9 BB 18
 C6 8D B9 E2 98 57 0F 89 97 0B 56 7A 67 27 A7 16
 9C F3 05 1B A1 C1 5F A3 A3 63 FD 47 87 09 2D 14
 02 D1 35 25 F4 8E A8 3D D2 B6 3F 18 B4 D8 0D 97
 A2 A1 EE 50 05 E2 65 30 D7 80 D2 58 D8 1F 62 E1
 A6 14 61 2D F3 23 83 6F C2 31 1E 41 79 0F 27 D3
 8C 6D 98 F0 2D A8 66 CA EE FD E9 0F CA 98 57 40
 97 48 F7 67 3F A8 94 47 72 1C 29 DA E7 80 40 B1
 FC 2E 01 06 36 25 78 91 C2 04 6F DA D7 82 C1 7C
 45 BD 36 6C 49 BE 7D 1E D5 F6 CF F7 02 D5 43 AF
 8D DF 11 2E BF 72 F4 3C A4 B8 9D EF 5F 44 DE 45
 57 37 30 16 7C EF D6 71 B5 18 58 07 D3 FD 98 90
 6E 44 04 DA D1 A7 45 3C 01 66 87 12 5B BA 77 39
 1E 21 8B 62 88 B9 BC A6 D1 C4 39 AE 20 5A DD 28
 C7 0D 94 A3 DE D3 4A 61 C5 36 4C 0F B3 A5 71 5C
 77 1F 09 DB 7B 86 02 AE 73 F5 DC A7 78 71 4B 67
 82 F6 F4 55 B1 D1 9B C8 B1 F1 5F 03 19 40 C8 5F
 40 7D 7D 19 BF 35 DC 01 92 25 5D 4A 65 33 04 4C
 8E F2 52 EF A3 81 D9 E4 6C 64 96 DD D2 21 DC C3
 14 19 20 19 53 A7 16 8A 5A 5A 7A 5A 88 A0 1F 7D
 AD EF 9A 4E E5 8E A7 E2 3C 7B 3C B2 0D BD 5B AC
 AD 5F A0 76 0C 53 4D 84 CD 13 BE 9B 0D C4 CF F0
 55 21 D0 5D 40 ED 2E 69 65 17 30 F1 65 B4 E1 A2
 95 9D CC 5C 1F 79 B5 35 4D DD CB 80 CE 1E 77 54
 A1 8A 5F 0E DC 67 FB D9 E6 4B 98 5D 64 D5 AA 19
 55 A6 05 29 2C 3F 24 ED A0 E5 C9 B2 53 CC 48 87
 F4 20 01 86 59 10 62 B2 B7 89 A7 60 A4 EE 47 91
 AF 0C 64 8C 42 8B 3B CF 6F D8 80 3F 0F B1 20 CA
 BC AC 94 93 3C 81 C8 0F 97 C4 BB D8 6D B0 E3 28
 AE 03 34 E0 A8 E3 A0 F2 E1 A2 D6 83 03 95 00 14
 10 02 D7 F9 F0 C9 1A D3 82 6E 4A 1B 85 84 47 31
 45 AC 6B 95 50 AB 72 67 CD 66 59 83 E9 38 B1 E0
 38 91 0E A7 52 8B 2E BA A6 9E 69 5B 98 1B BF 22
 B5 70 A2 AF A2 73 89 86 D1 01 8C 59 5C 8D 05 D8
 5E F1 DE BB 5E F9 BD 3B 47 92 32 B5 78 1B 94 FD
 3D FF 3A 77 20 00 F7 77 53 32 F0 0E 41 53 14 EF
 C2 72 47 62 91 F8 5D C0 7C 4B EC 02 71 63 14 ED
 BF F9 7E 1E E6 B6 29 19 EA 20 2E 99 06 0C C3 87
 21 61 66 03 04 45 BC 53 DF 01 09 50 F1 05 FE 73
 6D 1C 06 C0 82 B2 8F 7A C9 91 4D 12 68 6E 5C 63
 D8 9F EC CB 52 90 AB 09 6F 87 F2 94 19 EE CC B1
 3D BA 4A E1 5B CB F3 FF AC D8 3B DB D6 E4 60 07
 A9 72 0A 8E 39 7D 3B 8C 1C D4 C1 18 A3 54 40 CF
 F8 B6 CC EB 96 09 00 BA D4 66 79 F5 08 42 A1 D5
 9F E5 05 9A C0 35 8D 48 D0 86 8C 3C 5D 14 DF 8E
 4D D0 B2 D7 0D B2 60 69 AF 74 C7 4C 84 98 E0 09
 D4 AC 37 5C 09 F6 36 37 A8 E4 90 2A 66 00 CE AE
 F3 63 42 5C 5C 1F 8C A0 64 10 F3 71 CB 95 9B 28
 48 D0 E3 CD D1 8A 65 AA 30 A5 4A E8 F2 26 39 0D
 FA 4B E3 87 7E 14 C8 5B 87 55 D0 03 92 77 20 B8
 81 EF 4E 76 26 57 2B F9 7C DD D9 64 90 F3 AA E8
 49 69 F2 78 7F A4 E6 27 C0 3E 80 97 C2 0E 8C F1
 FA 25 9F A5 32 2A 36 32 43 55 E9 A5 F1 42 E6 61
 B5 3F 15 2A DE 51 D0 C5 CD 3C 02 AD E6 5A 36 4C
 1B 4E 88 96 24 8B 09 78 37 F1 A8 76 B8 96 F0 CF
 3C 10 3F 36 D4 3F 5D 3E D2 39 00 5C DF 32 49 95
 82 46 3E 17 0C 61 39 3C 53 76 6C 62 51 D8 A4 C5
 F5 B6 17 6C 77 EA E9 8F 8E 3D AE 2F 87 C1 D7 B5
 34 0B 35 65 98 33 F7 1B 50 4C D9 23 45 4F 73 70
 C4 FF 8F 7B DA 65 83 2E D4 E1 03 50 37 C9 3C D5
 0C 68 87 1E D3 DE 9C 0A 1B DF 9E B1 4B 31 74 9B
 50 31 7E 75 3C 63 5F AA 75 14 FF 19 69 23 CA 18
 8B B8 1E 7B B4 40 A1 ED 5A CA D8 13 CE 42 81 C8
 28 1A 4E 89 35 F9 B4 29 76 FC 7A 33 8E E9 1F 6D
 D8 BC E3 6D 41 26 76 9A 7A 24 4F 88 AA 89 C3 86
 01 53 8D 81 B1 26 D7 5A C1 56 38 92 FD F0 B0 63
 81 5D CB C9 66 8A 58 5D 42 20 0E 45 2C 05 E4 CC
 7F F3 90 07 EE E1 4D FF 5A B3 E3 43 07 6E E1 01
 F8 27 5E D6 AA 63 27 B2 C3 20 4C 38 08 17 24 6A
 09 A9 4A 8B CB B7 03 80 3B 63 D7 37 74 E4 4A 2C
 6D E5 DD B8 9C 01 C9 F0 CA D1 EE 94 1F B3 F5 43
 3B 8F B9 53 97 3A 6D FC EF F8 85 52 02 E4 B6 65
 90 15 75 9A 20 97 94 7E 51 14 B7 02 B0 ED F5 AB
 24 50 6A F6 7D E3 84 8A 5E 55 DF AC 36 4E 28 4E
 EA CB 10 1E 04 17 DB 7C 76 B2 B4 21 E3 54 0A 6E
 A8 04 80 AD 28 2D 04 D4 23 50 9F 8E 37 FC 8F 09
 7B D7 D3 F3 57 19 31 49 3A 1F 31 D8 38 0C 5C A1
 E4 2E 67 E9 04 7B 31 E1 AD AD BA C5 C3 62 58 E3
 B6 8E 3E A0 E0 B7 4A 62 7E 37 38 C0 A0 BF 81 06
 19 BA 0B 4F F0 7E 61 4F 1A 10 AA 16 AC 6F F1 C4
 A4 9E B0 55 5D 98 FC D7 21 A0 79 B5 A6 42 18 D6
 B4 61 32 E8 BD 37 A8 45 BE 7D 2B AE 0D FF F4 D9
 9F FF 43 8C 75 04 61 02 80 52 84 77 CB 1A C4 F4
 76 9F 5F 37 85 C8 F0 3B CA E6 FF 41 62 7A 93 D7
 6B 4C 31 76 81 FD AC 9D D9 CE 92 C8 B9 F7 52 EF
 08 AC 11 1B 19 52 B8 A8 17 55 A5 FD DD E7 C2 5A
 5F 95 33 2E 2C 9D D6 1D A6 92 8B F6 3C E5 52 BA
 D9 33 90 25 B6 11 BB BB A8 E6 81 63 AC 77 69 95
 42 70 63 58 A0 F1 94 C4 E8 3F E4 E2 7C EB AC 1A
 0C F6 B7 ED D0 E3 F6 9D 4E 1B 63 5D 02 2D 20 AC
 E0 BB 5B 6F AF 13 77 ED F7 FF 93 35 47 D1 76 CA
 89 12 1C EF 0E 8D DA 74 E0 14 1F 84 60 25 F3 CE
 1B 7C AF C2 F4 8B 0D 75 9F C0 AA 44 57 F8 2C E8
 19 AA 83 47 45 61 00 85 0A 88 D1 91 10 44 87 EF
 89 4E 63 0F D2 5C 16 29 21 4C 6C 2B F9 19 CE 10
 FA 03 8A 03 D4 0E 05 41 1C 74 26 4B 20 08 92 B4
 F7 BB D4 6D C6 C2 95 F8 89 DA E7 AA 55 34 4D C5
 8B EF AF 63 34 67 E9 8B D1 D6 6C B5 5E 58 5B 1C
 FA 91 97 74 72 66 51 EF 18 24 DA 60 E3 71 A0 6C
 2C B3 38 01 2B B7 FB A1 4B 82 97 80 2B 06 DA 06
 DA A4 B2 35 57 1B 00 A6 82 A1 EC 78 54 EA 3D 6F
 62 58 C4 66 1F E7 45 AA CD FE 56 75 27 1B 00 A2
 36 9F 11 D5 CC 70 EC CF 4E 9C BA 97 38 29 81 5F
 05 71 EA B7 8B 45 A0 FF FF 3E 94 85 E7 FF BE FD
 2E 92 76 43 25 A9 A3 D8 22 B4 77 58 A1 74 74 F0
 7C 35 6C C3 45 12 25 AB 57 E9 0B 97 0C 62 91 2E
 B4 7B 5E 13 A2 AB F9 D9 54 4E 15 73 45 0D AC 47
 50 9A 8F 62 CD CF 87 F3 60 E2 61 75 17 A5 39 DC
 08 D9 9C 56 DC 7C 8D 27 04 4F 73 39 BB 4A E9 42
 5A DE 1E B1 90 21 5A 61 76 E6 F4 33 42 6C 1B A5
 74 57 E8 D6 C8 BF 74 A3 3C A2 67 8D 47 77 43 C5
 AB A3 02 EA EF AC 0D 8D 13 5E ED 65 D3 3D 28 F7
 C5 E7 AD 84 B2 C6 14 FD D7 B4 A8 9F 8E AE A9 BE
 86 0F 90 B7 00 60 25 D5 CF BB EA 6A C4 87 15 CF
 B4 C5 29 51 25 94 9B FA 98 E6 E0 83 F0 42 42 4B
 B4 78 C7 B7 D8 FE 88 A5 77 F2 22 8E D0 D7 5E 5D
 F3 AC 34 59 60 A1 23 D7 F8 04 51 30 0D 0E EF E9
 6F B1 77 B7 E8 29 ED C2 49 48 0D 82 C1 15 95 0B
 A9 04 0B F8 68 23 24 9B BD EB 4B A1 A5 E9 E6 A4
 B7 2E 7F 59 DF E9 D1 BF D4 0C 2C 5D A6 19 F7 0E
 C1 90 09 83 06 A3 83 52 A3 D5 EF 76 AD 67 93 EC
 EF E1 9A EF 69 D8 75 F1 B4 89 E0 29 CC FE 0E 05
 69 CF 25 1F 6A 99 B1 BC DC 51 C0 69 47 BA B8 93
 45 F4 B9 F8 C2 F9 4A 78 F8 00 E3 16 15 79 9F 53
 57 71 E3 11 CC 93 7F 7B E2 40 36 BF 81 DD 3E 9C
 59 85 93 90 F2 ED 68 54 E1 64 EC 61 7D E9 CF 02
 79 B9 A2 BD DB 5B 29 39 E7 B5 6A 6B EA 17 92 32
 A1 DC 4B C3 21 22 12 05 91 33 62 9B 7D FF 50 34
 77 0A 09 E5 A1 E6 22 C1 97 FE 68 1F 1D 73 AD B8
 42 4E 6A EA 2F E2 BE 7B EB CA 97 6F A7 C7 3B 43
 EB 1A 81 A8 BD 02 42 10 9D E9 18 23 B1 E6 D0 D5
 3E 5A 95 EA DC 38 BF C6 F8 9E CA 63 5E E8 CD A7
 A4 7E 27 E3 3D D9 09 D5 CD 4B DF 94 18 85 59 0D
 75 C1 A3 8C 41 AB 7C 2A 21 04 CE 3A 2C 58 84 07
 9D 10 BB F8 F2 51 DC 44 A2 E1 D0 49 14 AF 56 B2
 D6 85 3E 9A 93 6B CB 05 B4 50 31 DD A5 D8 47 FC
 2B 11 20 3A B4 D0 BF 40 99 3D E3 7F E7 E7 EA AE
 3E D8 D4 AD 3D F5 A4 60 EE B4 C3 EA 91 93 D5 07
 85 67 1D 9E 6A 02 FA E1 C3 26 F8 7F 86 94 EA 33
 2E 45 7A 66 41 B8 88 84 6D EF 06 3E 35 90 F3 2E
 71 A1 BA 73 E1 E9 77 02 42 09 A7 63 D3 69 A5 5E
 8C 0A 39 74 26 0A 94 05 58 B6 D0 6D 7C 13 F7 7D
 4C 02 40 49 B3 BB E6 3A 29 38 97 07 C4 B1 57 F0
 49 F7 DD 3A BD 38 E8 AB 6A 98 49 74 22 83 5D 97
 3B F7 41 3C 13 B4 09 BB 9D 59 36 A7 B0 EC B0 A7
 40 83 60 CE 6C 4B F5 E2 CE CB EA D1 DF 08 E6 B4
 96 14 E4 4E E3 BA 10 D9 90 5E 5E D2 68 13 96 59
 31 04 E6 27 FD 42 8E 2C FA 03 1C FE 16 E7 04 6D
 47 F8 CA 25 68 C0 3F E0 90 AB B9 61 AA A3 0E 03
 82 64 8C 6C 49 73 68 35 70 33 65 70 56 C7 91 18
 0D 1B 88 1F 2D A4 CF 4D 96 A7 FF 43 79 C6 75 B3
 EA 42 8D 1D 93 E7 4D 39 B3 D2 C1 34 D4 10 6D 9F
 A6 30 01 DD CF 4C 62 0D EC 99 37 2C 79 9B A1 69
 03 9C C2 3B 83 93 03 83 B7 5F 35 5F 8C AE 61 0F
 99 AF 94 5A 75 B4 D6 B3 DD 7E 46 93 D2 62 E6 33
 C0 E7 55 73 28 4B 56 85 56 A7 1F D8 B2 21 03 F7
 4A CF AC 99 73 FD 27 BB 33 E1 99 5B 86 42 D9 4E
 C9 E2 72 78 25 CA 82 D3 00 9E D7 E3 C1 0A 48 38
 81 EE 51 E4 7A B2 52 05 D9 42 3B 0C D3 00 67 6C
 A2 3E C1 6E 55 3F 21 79 DD 70 7E EE 8D 32 22 EC
 55 42 80 33 65 D1 61 C3 E3 A4 80 F3 A7 99 4A 66
 23 F0 A4 9E FF 8E 32 B9 37 93 2F DA A9 A8 5A 67
 B0 E6 99 E6 64 D9 36 C7 F9 EF 34 12 87 8B DF 21
 F2 95 7E 82 31 98 CF 87 C0 4A C6 D9 AD 7A 3E 53
 E1 73 0F B9 45 53 FB 35 CD B9 09 F7 06 C1 C6 98
 E3 29 DD 1A 01 CE 37 51 15 AC 85 08 51 CC CA 03
 83 A7 11 FF DA 45 25 1B 81 EB 94 12 79 43 9B CA
 C3 9B 26 DF 4D 12 F4 23 E3 95 A7 C5 B5 15 49 96
 F8 CF D7 83 A2 52 9D 12 B5 60 9B 73 DB D4 CE E9
 CF D3 CE E4 8F D3 4D BB A5 DC 97 F4 2E 3D 0E 26
 3E 86 CD A9 C7 19 66 81 9D 87 E4 66 56 0A 75 D5
 F8 D7 3A 95 65 EF ED C3 6F 6B 65 7C 79 0B 48 51
 B2 ED AE 8B 7C EA 65 1B 6A 85 5F 6D 2A 9A 67 2C
 BB 1D 0D AF E5 91 E8 52 25 A0 4E 1F F1 50 99 F7
 C5 FE 5F F5 18 2F 3C F3 D4 7A 36 62 74 3D 31 D2
 29 97 53 22 CA 90 0B D3 D7 C3 CD 17 9C 4B 91 5F
 5F 19 1F 7E EE EF C2 6C AE 42 A5 D1 15 48 CA 46
 02 C2 27 21 8E E3 4A 3D F1 D2 F2 43 BE 12 02 42
 AF 5F AA D5 FC FF 2F B0 5F D3 F7 89 07 E6 39 A2
 0D 55 9E 01 1F 45 72 22 F8 32 CB 4C FC 1F D8 7A
 23 05 45 96 B6 D8 0B A6 FE 03 01 8D 70 6F 79 44
 5E D5 E5 46 1C AD 0F 7E 7A 41 02 65 E3 C1 21 B4
 64 A7 D0 C0 CD 08 36 49 7B 11 A5 E1 60 F0 ED 5C
 DF 36 7D 7C 1B 13 DC 45 4E 81 62 4B CF A4 33 1E
 D5 C2 D1 41 71 20 20 08 33 CC 17 66 86 E1 32 5C
 57 F6 DF 1E 8F 8B 6A D6 6D 46 59 AB F0 8C FD 15
 90 5A 54 B8 D2 F5 2A 6D 5F BC C4 D7 97 F9 3E 82
 62 61 0F 7A 90 49 6A 27 76 39 4B 23 75 E2 37 72
 3D 7F AE DC 9A FF 03 34 F1 48 66 B9 A2 C9 F0 17
 2F 4C C7 22 BC 66 21 E8 8E 2B 58 C0 61 E1 BA 96
 47 DD C9 33 C1 96 B0 2C 9C 0E 25 AF 66 E8 D0 1C
 CD 33 CD 2E 6B BF 63 1C 86 38 AE 23 CB E8 8D 26
 88 E0 97 E9 8A 16 2C 91 92 9B E1 AE 5C DA 88 7D
 91 49 E6 8C 9C 89 01 DE 07 50 6F 1E 0B D2 1F 2E
 54 73 45 C8 39 EA C9 13 66 EE A8 01 76 92 B7 A6
 27 76 35 4B 70 73 A1 71 09 91 B6 89 85 ED 33 36
 44 ED 86 8F 9C 0B 43 46 45 CC 03 AF F9 F5 8E BC
 44 E7 94 4F F6 33 A3 41 0E 3E 6C 7E 3F B2 19 3B
 B9 36 0B 34 DE 11 F7 43 45 CA 16 54 3B 16 35 ED
 46 A4 6C 77 9B E1 13 61 59 42 50 9D DF 66 30 C6
 83 03 4B 34 A4 18 2A 4E 96 2B D3 DA 7A 56 6A F1
 93 11 40 16 89 99 1B 90 8E 68 72 B2 E7 8F CF 8C
 A9 52 9D 92 18 29 CC B5 E6 5D BC AE 71 AF 04 9C
 49 E9 A6 74 84 16 96 A1 6B 60 F5 49 9C 85 EF 14
 7A 7D B4 C1 A8 68 58 23 5B 33 57 9C 1A A1 D5 10
 FF C9 70 C9 AC 29 5E 24 63 03 89 C6 10 69 35 83
 29 BD AD 11 A1 22 DD 76 21 21 D4 5B B7 71 FD 96
 80 64 D0 F7 FA 4B D0 20 41 98 1C 2C A7 FB 03 E8
 8C 23 63 24 EF F2 FE 68 1B DE 28 19 C6 F5 8A 6D
 9A DA E5 24 4E 7F 9F BB 3F 21 A1 1A C4 CB 01 B3
 C7 CE 0B 8E AA 39 8B 5A A1 8C 1A 06 98 8C 3D 0A
 B5 17 25 A2 97 8D 1B E6 6C B5 2A A1 D3 3D 47 56
 DD 34 99 5D 47 A8 FD 03 CB 88 84 55 89 1C B6 33
 ED 91 BA 5D 5B 31 5D 04 4E A3 55 46 F1 36 10 A3
 11 80 ED 57 0F 10 7D 10 51 82 B2 26 D8 D9 7E 20
 7E 5B 29 DF E6 BD 9B 17 D2 49 9F BB 08 04 36 F7
 DB DF D0 EE 1F B4 F5 0F 52 1A B5 17 A7 EA 7A B1
 47 02 42 22 66 23 EF 1E 09 B2 28 FC 0F 74 72 F9
 FA 31 75 52 E0 79 F4 0E BC 8C A1 93 54 33 77 1E
 A7 CF 8A C9 B6 12 58 1E 81 37 D1 2E 70 70 CC 81
 8D 65 EF E7 F1 A6 2E D9 53 56 17 8F 2A A8 BF 87
 32 09 3E A3 2E EC E3 CE 49 AD 67 F1 E9 02 7C 84
 CF F0 EE 87 C2 B2 3A 74 42 1F E2 5C 25 96 63 1E
 DC 67 85 21 B6 AE 67 ED 80 1A 8A 31 93 B3 20 69
 1D 6F 32 7C E7 04 BB DA FB 2D 59 DF EB B9 CD 76
 D3 52 FF 04 06 FF C7 73 A1 7C 94 F8 33 DA 90 56
 C3 E1 CF CF 86 4A C4 C3 94 22 49 2C 1C 27 FF 45
 1B E7 01 A7 AB 35 6C 5B 4B 84 78 66 A2 3A 9A 08
 E9 71 29 D8 07 1E 37 A2 06 BB 07 E2 27 75 E4 20
 2B E6 A4 4A 9D 51 79 18 4C FE D6 50 73 B2 55 A8
 A2 AB C4 71 02 BA 80 11 40 D7 C8 CA 6C 42 E9 5C
 16 CF BF C2 3F 92 E1 50 5A E7 51 3B 8B C6 F0 CC
 14 9C 45 CB 78 F5 B7 66 A5 DC 68 D9 45 B5 DA 33
 2C CD 99 CC D2 7F D7 C7 BF F3 E7 D9 0E 18 C5 14
 FD 07 1B B5 0B 5F 22 13 7A 8A 5C 9A 52 7D 18 70
 97 00 26 D8 2A C4 EF C0 AB FE 69 ED FC 14 D9 98
 AD 93 50 FB B4 9E B5 5F E7 B3 A1 67 8C A7 9A 19
 C9 78 A6 88 31 13 40 08 2F 5B 3E A1 94 76 BF AE
 13 44 B4 6E F7 7F 08 40 B3 51 92 7A 94 2D 5D 71
 FD D1 42 29 BB 10 FF A1 52 76 73 F2 E7 65 E3 F8
 59 E5 C9 FA C8 4D 95 19 CE BE 96 B8 F7 BA 46 E7
 39 0B 57 A4 8A 44 30 B4 FA 5B 4C E1 2B CB 26 89
 78 FA 0F 89 A9 71 53 5B 88 CB DC 2C 06 19 A2 93
 84 B8 22 D9 A4 BC CB DF 7D 3C 8F A6 82 FF FC 14
 00 3C DD 0C 34 B3 A2 B0 AC 2A 3A 2A 57 AA C8 A2
 DD 67 29 76 BA 23 7C F2 90 4A 0C 1E A6 AC D7 18
 85 16 F8 A0 B9 29 82 4C 08 6B 10 8C 29 58 F3 83
 3A 7F 6F A0 9C 6A E7 E2 5D 94 86 45 5A 93 C7 53
 5B A3 E1 68 22 9D 64 06 4B E4 95 07 A4 39 96 C5
 EB DA E1 13 BA FD 78 C9 C5 4C 5F AF F2 2F AE 09
 47 D1 BB 44 3D C2 86 89 62 B0 C4 03 E3 36 28 5E
 4F 42 CF CB F2 2B 3E 91 EF 96 D1 6B 18 0C CE D3
 6C 2C 8D 77 23 88 80 A9 9A 99 A2 DD 0D 77 E2 9D
 0D 7F CB 2C 41 CB 7E 20 A5 67 CB 16 B9 F9 8E EE
 2E 4B 21 F0 26 BA 28 CA 9F BF 55 F9 D3 B4 E3 91
 64 A1 2E 1C 85 5D EE 38 42 F8 F6 3D 49 E3 47 1D
 43 05 9B 7F 95 1C 8B 37 C4 EA 68 5A AE 5F 69 2E
 98 2A 39 E3 46 25 39 09 CF D7 DB 46 73 A9 0F A1
 AA 05 C3 AE FD 73 8C EB 14 9C 28 F1 07 21 C1 C0
 9F 9D 4F 82 84 98 A5 8A FD 1C 91 D3 5F A0 40 2E
 43 06 C1 EC E5 EA C5 61 4D E7 C3 7C 8D 1D 1A EB
 47 12 CD BE 95 CB 62 60 E2 69 A0 A9 3D 62 61 B2
 DC 6D F2 41 18 2F A7 65 7F 7F 91 0F 5A 75 C7 88
 94 F9 A5 7B 2A 87 42 04 21 2F 48 AC C8 E7 90 2C
 67 9C F8 C2 AE AC 23 7F 19 46 93 95 B9 67 38 18
 CD AD 30 6B 92 9B A3 E8 A2 CE 21 F7 82 30 9E C2
 0E 8A F1 A9 F3 8F 6B FA 0F DC F0 96 C7 0F 8D 1E
 44 E3 FA 7E 79 8A 87 67 94 70 82 60 96 95 8E C8
 E0 02 BE A3 A3 E0 4C CF 82 E5 55 07 5D 8E 25 37
 E5 DA 18 0F F3 95 83 DB 24 B3 1A 0D E6 52 99 9C
 82 D4 71 7E 9D 6E C0 D7 08 F6 6A 01 8D 44 0D A1
 C8 BD 19 94 88 C6 72 65 82 BF 02 CB 6B 78 C5 06
 02 8F 99 BE 69 62 82 B5 09 5C 39 93 65 81 C3 B6
 84 5B 43 68 20 19 7D DF 76 1D CB 5F 8A 01 5E 61
 7C FF 10 1E 64 A0 10 FC 26 AD 6C EE 61 82 93 E4
 F4 4A 53 8A EA BC 6B AA 4E BC 61 87 19 33 38 3A
 42 34 05 74 87 96 07 5B 6E 09 EA 71 7F C1 01 22
 C2 89 1E FA BB 59 D8 54 61 AF CC CF 39 F6 15 84
 05 27 B2 F8 CC D0 59 0B 22 DE CD 1C 8C E3 1B 03
 84 4E 7F 40 85 6F 85 DF B6 5A D5 25 71 2C 3C 9D
 67 80 3A 47 A7 84 C7 90 02 BB 9B 5C 67 D1 B5 30
 B6 C5 6E F0 B3 81 38 52 23 7C 11 09 7F 26 8C 01
 B6 BA 62 54 36 7C 54 F8 9E AC D0 5D F1 65 2E 36
 B5 48 56 38 7A ED AA A9 49 CB E8 F8 BE E3 7D 65
 B6 F0 23 C5 0F A7 62 81 20 D8 96 05 E6 43 DF 4A
 5B 23 41 F8 4F 26 F6 14 72 67 00 67 9E D0 38 81
 8A B0 44 E4 56 F4 98 7D 47 28 C4 A6 18 FC 4B 81
 08 73 BC 0A 0D 29 E7 2A B5 21 43 FF 7C 49 D9 E1
 EA 24 0C 69 71 A2 46 E7 BD 81 57 76 D4 FC 88 DF
 EC 00 9C 32 78 E4 67 5B 71 D7 9B 9B 18 31 6C 83
 27 9A 9D 05 E0 6A 44 09 0B 80 7E 9D 60 59 94 CE
 D7 31 85 9C 21 93 14 6F 50 9E 01 85 5F 5A F0 A3
 B3 76 DF 63 4A D6 B8 BE 49 27 0A 8F 1F D8 DB 0C
 5F 06 15 74 0E 5C F0 1E 6B FB 28 A6 59 5C 83 2D
 BC CE D7 29 AA 6B A4 E8 6B FA C6 EC 40 F1 EC 44
 23 5A E7 B1 A8 7E 1D 0A 56 B0 51 E3 A7 C9 69 3C
 3C B2 7F 7F EA CC 03 F6 E8 7D 99 BA 97 54 29 BB
 B3 EC 53 47 DE DD 2C 8B 57 36 F4 98 65 32 91 4A
 D6 FB 40 4C 5A 56 B0 44 30 22 F8 6D E9 0E D9 44
 02 3F 48 2E 86 85 CA F9 6C 1E A7 83 83 0B 19 3E
 33 8E 55 13 A5 49 36 04 CA E0 EA A3 6B DB DC 58
 97 4F A2 DE 61 D0 5B E9 97 85 43 FF B1 EA 5B DF
 5F 00 81 1A 19 A3 F8 AF 3C E2 D2 83 B7 30 CC A6
 F3 95 B2 6B 75 57 83 CA 71 96 CF 0D E8 35 CA 0A
 2F 78 C6 BE 86 D9 02 55 28 64 59 24 01 AA D7 40
 82 FE F1 25 01 C1 C3 3B B0 26 B4 9E DB 2B EC 55
 BE 3A A3 73 DA 4B DF AF F5 D7 84 08 BC 2B AA 9A
 ED 41 34 36 5B 8C CE 06 1F 2D E9 74 CD 38 4D 16
 FA 04 EC 5B D0 FF B1 DD DC 4B 3B 5D 0F 22 65 54
 DF 02 43 FE C3 64 F1 CD FC F1 2C D8 D6 EB B5 40
 EC EB 4E F4 E9 FE CF 8E 2F F5 82 35 53 22 D8 38
 8B 86 FA 5C 54 8E 27 82 D5 BF 41 50 DF D2 FF 2E
 23 92 24 A5 F7 59 20 2C CC 7E 93 78 22 91 64 B4
 F9 73 0B 6C 6D D0 9C 00 92 75 CA 09 10 76 93 AF
 C1 26 89 BE 2C 26 CD 68 4E 2E D1 A4 8A C7 EF 15
 F9 F0 B2 20 D5 E4 1B 37 6E 6A 26 74 8D 8D EF 92
 3E 40 E6 28 D5 41 DD 32 31 FD 49 5F D0 F5 40 02
 31 3F 10 A3 5E 87 3D F9 27 D6 6A 2F BD F2 D2 09
 6D 31 D5 FA E0 73 BC 07 FE 8C BF 53 1E D4 2B 15
 7F 33 8F 0D 0C B3 63 32 15 E4 08 C1 16 C2 1E CE
 B2 7C 80 68 5A 98 13 A7 A6 86 D1 6B 47 CC AB A1
 A6 D7 4D 42 BC 4F 02 A7 DE E6 F9 B4 4A D6 24 F8
 C5 51 05 04 3F A1 59 45 21 62 80 F7 8F 0A E2 0F
 94 7D BF 29 AA B1 9F E3 03 1D 07 F9 96 9C 03 C8
 11 85 13 1D 20 58 18 CB 8C 4C 6A 55 0F 2C 8D 92
 34 09 17 54 56 4E 69 F4 2D 17 B7 25 D2 17 3A 54
 0A B4 B7 8C 6D D9 44 1C 46 0A F6 DF CD 8D 50 65
 EC A0 EA 80 92 9D 25 AD 01 9B 7D 51 DC 96 B1 BD
 00 63 10 15 80 72 F3 02 A3 7A EE 68 A3 C4 07 0A
 4A FC 26 AD 4E DD 2F FF CF 02 D2 CC 27 5A CD 3D
 22 03 81 0F 62 3B 9E C3 BA 1C A6 97 64 6A 4F 89
 B7 96 BC E7 85 B2 A2 06 DB EC 7A 23 5D 72 4E 63
 3F 8A 1B 21 C8 39 81 DD 5E EF 40 0B 2D 38 74 76
 05 3B 2A F1 08 33 3D 1F 92 C2 E1 C8 77 F2 EC 24
 AA 3E D0 A7 BC AD 1C 5E 91 02 AE 86 99 2F 43 AE
 F4 61 48 26 00 3C F4 E7 AD 1F F3 09 B2 8C 23 BA
 6D 50 A4 C0 A7 6F E6 01 C5 60 FE 47 7F 4C D6 18
 CB 75 AE 60 C7 CA 42 75 D7 58 40 24 E0 FE 3F 1B
 F3 94 8C 46 EF 1F E2 53 E8 A2 6A 58 B0 39 EC 2C
 64 3F A5 24 84 03 AA A1 88 E5 FC 5E 82 AF DF 05
 C1 39 6F 98 DD C9 62 E9 C1 54 5C 20 7A 85 73 B5
 7B 72 89 6B 75 5A 6F 12 BF 07 2B 6B E5 BF 36 7B
 65 75 C4 21 87 95 45 58 C4 C1 14 92 87 0A 86 B6
 E5 68 74 43 58 BD 61 FE 04 DC 51 0A B9 FE 29 FE
 0F C5 51 EA C6 1D C9 B7 D1 01 51 B2 DB 15 CC A0
 18 8F 13 B6 1D 75 4D 6E 88 FA 0C F4 98 7B F5 88
 96 A9 CD A3 BE 40 16 EA 3C 9C E8 3F AC BA A3 D2
 FB 5C 35 1E 0B 53 F7 8C 6A 63 F5 4D D1 EE 5E FE
 68 D5 1D 1B 54 27 5E 4F 35 BF EB AF D4 E5 90 12
 00 F2 1E FE 77 5A 92 06 3D 02 58 80 B4 71 FE 22
 94 89 C5 13 4A 03 CD C5 7A A0 FA 92 47 76 1F 5E
 F9 0D FC FB 54 B1 C4 64 01 B7 F6 3D 44 90 29 CB
 2A B6 3F 3C C6 EF 2B 44 5E F7 98 CC 32 53 69 7E
 AE 44 FE A1 21 F7 9D 2B F2 1A 61 CF 58 74 0E 3B
 98 12 EC 81 0B 60 BD 53 48 D2 44 83 43 D1 AF 00
 CD 06 DF 6F 14 0E 75 AA 35 A6 A7 05 B6 CA 50 5F
 BC 2E 5D F9 6F 43 88 C9 2E C3 7D 74 E9 76 5A 36
 03 57 F8 BC 4E B7 EC E1 21 FD 42 6E 68 60 81 FF
 19 D0 86 68 DC 3E 7E FE FB FC 09 82 99 9B 52 A0
 12 70 7F 0D 71 1C F5 74 7C FF 8A 53 FD 06 D2 28
 A5 7A C1 EE 53 2B B4 25 5B 83 0A 76 13 9F AA C8
 77 5C 6F 9F 40 A9 FC 06 B1 BF 41 DC 96 52 D5 92
 A0 AA 79 71 27 B7 33 2E FB EF 48 B2 3A 25 DC 3B
 44 5C 6D B7 97 4F 46 4B BC 02 0F 43 CF 51 16 12
 82 92 59 5A E6 DB 03 A0 68 11 83 A4 6C 0B 2F AC
 AE 56 7A 1E 3E 35 C5 81 40 73 C4 B2 A5 17 6F 66
 8F 43 44 C4 78 98 29 D3 B5 A6 7B 7C 9D 35 F7 84
 F2 D1 C1 7C F1 33 AC A6 3E 46 6B 35 B9 D7 C1 F3
 1F 7B 82 1C 30 81 E1 53 71 C3 84 31 D0 D0 07 57
 FA 53 85 9F 97 97 DB 1F 75 27 AA 08 92 3A F7 B3
 BD BE 06 9B B2 9E A6 98 FA C7 AC 74 15 97 E5 0D
 FD 95 97 E5 D4 30 A1 24 D2 06 D6 03 45 BC 51 76
 5E EE A4 32 E0 A4 95 9E DB 51 2E C8 2F 48 24 56
 6F 2C 45 C5 21 FF 1A 23 38 B1 67 A3 90 4A 16 2A
 51 43 D2 CE 5F 4B D1 2A 95 5D C6 11 B0 46 1F 63
 3F ED E7 FD E3 55 33 AD 62 E3 E6 A1 80 E6 C4 3F
 C4 1E 7F B0 4D 08 75 F5 85 94 E7 7B DC 85 EB 0B
 C6 2C 3E C2 A9 05 34 24 BA 6F 07 47 A0 46 84 24
 F2 7B 9B AE FC 76 8D 9F 73 54 97 0F 59 81 C2 6B
 EA CF 47 42 9B 9C C1 9B B3 E2 55 62 A5 DA EC 08
 73 A0 B1 DD 60 4A 86 6B 76 95 31 05 DF D2 E3 F4
 6F C9 0F 9A 08 EF 4F 03 D6 58 B9 F5 69 57 78 6E
 20 1A 72 A9 C6 98 C3 13 E5 90 F0 2B 33 A1 B1 32
 76 A0 C4 09 12 53 41 70 C1 7F 82 CC A2 4E FF 42
 A2 3B F3 55 14 45 F0 74 60 68 30 27 50 7B BA DF
 C6 9A 75 37 C5 1C 8B B6 71 18 91 70 5B 1E E5 FB
 2C 4E 2B AC 69 9D F5 CE FE 24 8E 9F 8A 91 2C E2
 C5 6A CF A7 05 68 F3 9F 75 9A 76 7F 77 DD 68 0F
 71 24 64 D5 73 DC 7E 9E D1 D0 A7 91 51 3A F1 82
 79 1E CD 1C FD 51 AA C0 60 91 5A 46 1F AA 60 83
 71 18 F9 22 B4 2F 98 5C BC DD 9F 7B A0 1D 7E AE
 69 85 0D 4F D5 F3 2F 10 49 A7 2E B8 55 6B 8B 51
 09 5B 90 3B F6 00 67 78 5F B9 B4 C2 C0 08 C0 DF
 BA D6 46 84 95 8D 9E 80 BD 54 39 7D 0F D2 FD C6
 9B F5 80 83 57 A5 6F 2E 7F B1 F1 3E BA 64 70 C7
 E3 85 76 D4 12 E8 12 C9 E1 37 1E CC 95 B5 02 33
 C5 0B 81 92 DE 22 B8 1F 58 3A 2B BA 3B 6C B5 34
 88 39 78 50 3F 04 20 7B 8C 4C 39 3E 33 60 C5 68
 BA 9A C3 DE 6B 80 F0 F0 65 94 E8 86 B9 6C C5 32
 55 7C 88 C3 1F 0A F5 15 5F F7 36 79 D4 4B B1 20
 E2 DC CE 1C 63 C2 3E FA F2 36 B1 41 72 C6 BC 9E
 E6 C6 57 71 7A 11 8E 18 7F 45 A8 82 2D FE B3 E5
 D5 50 43 DF FB EC 71 25 34 4A 63 F1 04 EA F9 79
 DF 0F 73 FB E8 46 1E DB 0A 5D A3 DA 68 3F 7C 0E
 60 22 B5 03 71 1C 24 C1 11 6D 5C AD CD 62 42 C3
 5C 1C 2F F1 8A 95 E0 65 0F 5E 9F 00 AB E0 83 04
 54 C9 A1 6F 34 3F E3 61 98 10 C7 13 40 B7 8A BF
 C9 30 2E BC 5E 1F DA 96 7D CE 8C EB 78 54 3D 1E
 38 DE 3D 57 44 83 23 08 62 AD F0 68 C8 8D 9B 75
 69 A7 80 0C E1 73 3D D5 37 B2 A6 1C 54 FD DC 7C
 F9 27 AF A9 65 1C B7 BB FB 68 B3 A3 DA F5 24 E4
 E0 0D A9 C1 1A B6 A1 BF 29 C6 E9 14 F5 34 B3 62
 D6 DC E8 4F C9 03 F1 01 69 06 3F 40 B9 01 5C E8
 FD 4A 50 BD 06 B9 7E FB 75 D8 07 94 F5 78 29 B9
 60 F0 28 92 99 90 A5 61 B1 E1 C3 1B 41 24 5F E9
 D8 FF 6E 73 11 C2 37 C4 03 2C D1 C6 2D 10 CA 76
 04 BE 47 CC 75 D5 0E 65 C6 14 87 56 DA A6 54 41
 EC E0 75 96 74 E7 3C A3 0E 92 6B 2C 88 80 85 02
 89 A3 50 49 A5 2D D1 71 73 80 D4 01 64 1C 6C ED
 C1 98 99 C3 D9 1D CB D9 F9 73 8F F9 9E 55 8B F6
 80 3C 0F FA E2 8B DC 0C B9 B2 79 D3 93 43 6A 74
 E2 0E E0 3F 82 50 D3 83 2D BD 06 17 FE 79 15 6E
 AA F0 45 41 93 3F FC E8 A6 41 D6 7B 2D DD D7 D2
 24 4B CA AF 3A 99 36 35 DA 85 73 EF D9 2A 32 8D
 E2 CF 15 E1 FB 47 51 2D 7B FF 58 67 78 7E C8 60
 1F FC 4E C4 61 63 D8 AD 1D 64 68 7B 2F 3E EF 17
 C1 BA 71 55 11 07 DF 4C 8B 28 48 8F F1 DC D9 59
 99 29 8F 14 E8 40 7C A6 65 74 CD FF 3C 5D 41 9C
 99 AD 87 07 88 90 B7 FC 1E 48 F6 CF 24 25 0D A8
 FD 16 77 95 E2 D6 F6 3D 08 BF 26 0C 9D 87 29 E0
 38 82 FB 93 DB 89 9B 7F 4D B5 9F BB 13 B6 34 F7
 5A 96 5E 40 8A 3D A0 66 70 B5 4A 69 81 F8 2F 6E
 1E E0 00 E9 1F FC 19 AB 59 27 98 22 C6 B5 B2 CD
 34 8D A6 72 59 CA B2 EA 51 69 E5 84 90 88 BB C7
 49 22 EF 4B 50 10 66 EE 86 06 05 82 96 58 AD 31
 AD F0 DC DD 10 17 82 D1 77 EF 9A E1 5E 18 21 37
 A4 1C 85 50 39 13 DE AE E3 B1 14 78 C2 20 35 F2
 9C AE F7 10 17 D7 FD 4C 07 0B 75 9C 47 1A 7C 1B
 C4 EB 02 0B F0 E9 02 59 53 AB F5 C0 6E 7D 8D 62
 F1 1E CA 66 0E BB 5A 5F 02 BB B4 1A 58 84 4E 25
 4A 50 D6 B8 99 1D 84 5F 47 59 85 D0 B4 2B 55 EF
 C4 7E FC F9 CC 69 A4 D8 DE 1E 4B 0B 22 9E 2E AA
 47 6D 4A 26 D1 D0 26 40 27 EE DC 5C 02 EA D6 8E
 15 AE 55 C6 CB 5B 05 C2 AF B3 C5 90 9A 90 F1 D5
 A4 36 45 58 82 6A FC 89 46 CC 4F 67 AA 8E 63 F8
 2D 32 23 B4 83 D5 C1 A9 57 A0 23 CB FD 05 8D F8
 A4 B1 FC EA FA BE A5 DC 7D 8F DE 4B DD B7 80 0A
 15 38 BB 58 56 F0 19 A2 CA E3 69 05 52 2F F6 AF
 FC 89 3E D4 16 5B 85 0A E7 05 D4 05 93 7E 30 65
 66 44 44 60 83 A6 88 E3 99 57 D7 B7 46 D5 23 AC
 7E B9 E3 62 3B C3 EE BE 24 32 71 71 48 18 4D 55
 0E 16 70 5D E5 D5 59 7C 80 2E 38 45 9B 73 80 61
 D8 D1 7B 9A 2A E1 72 4D 61 F8 DF 38 45 F3 1B E0
 90 F4 FA 5C 65 35 01 D6 49 A8 26 BA 99 08 39 08
 1B 84 D8 6C 8E 60 22 E3 E6 AD E5 D1 EA D2 43 8C
 BB 0D 15 BC C4 D9 93 62 71 18 12 49 8F 8A 9D 65
 17 C3 FE 07 F1 F0 CE 42 14 21 FD EF 24 1E 4D 10
 F4 4A 57 98 76 DB 05 C0 79 06 70 65 B0 12 B5 B4
 13 F1 4D 71 1F 22 4B FF 62 A3 15 D1 D4 66 51 EA
 06 A7 F9 CC D2 54 3C C8 48 30 00 70 3E 8A C0 91
 66 99 69 8D C8 59 D3 99 A8 D5 CB F1 76 F6 F3 74
 01 91 10 DD 82 FD B6 0A 6E D6 DD C7 F6 BA B0 80
 88 55 8D 64 E4 9D 22 85 62 4B BE 4F 92 E9 77 36
 2C 3E 19 72 78 BB 86 53 2A 3D 80 0C 82 C2 85 A1
 AB BA BD 0F 9D 7C E2 95 E9 64 02 5C EE E5 0B E9
 B3 76 77 E7 7E B0 82 40 DB BD B4 FA 6A 9A 5E 9F
 AC 4E F6 C4 B8 D3 1E 26 3D A5 E7 2B F8 AC C2 72
 10 3B 94 9C BE 83 51 BD 92 89 4A 7B 60 1E AE 99
 30 BE C1 63 C2 CB C3 D5 B9 58 AE 95 8B 33 C0 5C
 96 C6 6A 5C 94 ED 1C 0A 95 7C 06 6F 56 1E 99 C5
 4A 39 12 E0 BA C6 61 B2 6D D2 4C 1F F9 3D 66 14
 73 3A 8B DF 1D DC 8F 23 4D D3 86 B3 98 4E 83 07
 45 6E DF 23 AA 63 2E D6 63 D3 BF C1 83 48 8D DB
 21 5F 88 8D 19 EF 8B B2 B3 4E D1 0E E7 0F D3 49
 7E 77 D1 12 86 0A 46 FD AE EE D7 52 20 80 9C 32
 D7 81 18 DE E8 83 0F 59 94 D2 70 A4 0D 34 25 C1
 FE E3 A3 60 FF A1 18 F4 4D EC FE E5 28 0F 7A F6
 29 A8 AC 19 A5 05 2E 17 C1 48 07 3E 5F 9D FC 3D
 EC 36 EA 24 09 EF B4 57 7E 9F 67 25 37 04 8B 1A
 07 A0 B3 67 27 61 4A E0 20 15 61 33 8A C1 46 52
 5D D7 3D D4 78 2F 7D 87 2A 36 5C A1 B9 F5 61 E0
 13 C3 94 FF 07 54 FD 22 F6 48 05 F1 E3 14 4C 1E
 6F E7 83 A1 2B C9 59 50 52 EA AD FA 6D 9E E1 D0
 06 6F B7 57 14 98 C2 9A 69 59 37 BA 3C 88 13 92
 23 77 84 48 AF 38 82 93 B6 B4 3D 60 FE DB DA 4F
 0D 58 F3 E8 D3 71 ED D9 B3 65 5B 82 93 9C FE 11
 29 9B 70 6E B8 14 09 73 3B B4 0B BA B7 F8 5D CB
 0D 66 4A 59 07 92 04 27 15 8C F6 DB 7C 99 F9 8A
 2B F9 56 85 DE 87 47 12 74 EE FD B9 C3 EB 23 F5
 3B 6C 89 72 95 C0 E6 7F C1 39 15 C0 8E BF EB 35
 FD CA A1 C9 74 4D 1B B0 75 67 0F 72 07 A0 AC A6
 A0 3E 27 E2 D1 CB ED AE C8 37 CD 32 87 AE 11 CB
 A8 1C 07 0F FA 3B 88 77 E1 03 D6 52 97 D6 1B DE
 17 F8 66 D3 92 4E 3B 73 4E 8E AB 07 3F 21 22 A7
 26 F9 8F 3C 0F 05 1E 8C 62 AA 7E F5 37 DF 0A A9
 BC E9 9B 9B FC C4 22 C8 28 50 DC A0 37 12 9D 86
 CD C4 DF 76 43 BC 2F 5C C0 D0 2D 2E D6 CF 71 41
 D0 B1 39 FF 9A 5E CB 27 7F E7 24 CA 54 04 BA 42
 AF 89 FA D9 56 14 98 E2 CC F9 58 4C A9 64 C8 71
 F5 61 A5 0E FF EB 09 F5 EF 61 38 3A 12 01 8E 5F
 74 A3 47 28 43 88 22 8B ED B8 6F 4E 06 1C 88 17
 29 71 B2 E9 A4 97 FB A7 24 42 D2 BC 35 FC 1F DD
 59 BE 67 D1 D6 D0 04 55 2D 3F 61 31 AD 3E 41 50
 EE A5 C8 C2 FB 4E B5 23 A9 C3 FF A5 D3 1B F6 A0
 07 85 01 65 8E A9 B0 14 E7 67 5D 87 13 52 2B D5
 A5 B0 7A 9D 6E C3 A5 8C BF AE E6 90 F5 CA 7B 51
 D8 65 97 DC EA A8 E2 09 02 C9 1A 1E B4 CB 1C 21
 08 2F 49 A1 76 0B 93 A9 A9 C1 A6 69 3B 7C 89 7E
 F7 1B 8F CB 6B A1 46 BA E0 14 8E 8C 2C 3E B3 76
 4F 77 C1 44 C6 35 B6 86 24 68 DE 7E 99 40 14 D3
 BC C2 52 99 18 37 F3 35 66 52 20 DB 39 8B 4B 47
 4F 36 36 2E 2C C5 23 D3 07 F9 4F 2C 08 0B 40 36
 91 41 CB E8 60 FB 60 3A 49 BB 2F D9 33 5B 95 D6
 AC 4C C7 AA AA 9E 4E F1 14 9D F3 20 E5 07 4F 2B
 41 77 9B 7E A4 42 9D 91 86 E6 18 22 15 2A 30 EB
 BB 38 28 38 F4 12 0E BA A4 5A 3E 01 42 43 71 6C
 7C 36 9A C5 08 6B 6B 26 9A C9 BD B8 CC 2C 06 BD
 A9 2F E0 DB 36 1D F0 EC 7C 1A 88 3B D2 F3 BA 13
 5C 75 3F E2 FF 0C A0 55 57 B3 B1 9E E9 D3 E9 6A
 AA F1 7C AA 24 39 67 1C 99 34 FD 6B 49 C5 4A BE
 B1 03 A5 32 09 FD 5A 83 86 DF DA E2 F6 21 91 C4
 32 B1 FB BC 08 4E 01 CE 50 22 C9 1D 64 AF 36 12
 AC 1C 42 C3 B5 DB D1 01 62 08 84 AE 61 4D 6C CD
 33 24 8E 67 BD 49 C1 22 1B FC 41 0F 71 3E DE 7E
 C4 A2 E7 73 54 A2 87 FF CC 16 33 47 68 5E 75 EC
 13 97 B1 38 C0 35 4B 61 30 A4 1C E3 7E 18 69 79
 98 7B 86 94 F9 BB 4A 71 DA 58 E4 80 32 98 19 4D
 75 98 94 0E 66 77 7A 10 61 9B 22 D9 7D A8 EE E4
 EB 42 60 DF 63 26 A1 19 E4 47 07 3F CB 2F 15 80
 75 FA 22 F5 CE 7E 62 C8 AD 84 EE 90 E7 1D 82 0A
 9C B4 0A 1C D2 84 5B 0C 06 59 B8 FA D1 63 E8 9D
 5E 0F 26 C2 3F 6E F9 DE 0B 02 FD 5F CD 3E 1B 17
 32 39 A3 3B 70 95 44 80 18 E5 CA 66 79 18 0F D3
 7F D0 DF A6 77 A5 A7 1A 39 ED 87 FD 62 53 3E 35
 33 6A 69 53 08 CC 64 3D 6E 3C C8 13 FF 17 7F 67
 0A B9 9F E4 12 03 81 5B 9E 27 A0 A9 69 51 84 4E
 48 E9 DE 02 26 2E 8C 63 80 1C 61 E5 B3 44 AD C9
 62 69 38 4B 0D BC 5C 89 CC 21 C1 2F 6A C8 C5 B5
 7C C6 1B 7A 37 A3 06 F3 B0 61 BD 87 C7 45 FB 7F
 C2 4F 8E E1 BF EF A6 F5 42 F9 ED 8E 27 2D B0 B4
 60 0B 6B 03 57 7B B7 D6 AC 9A 61 F0 2E DC C9 49
 7F 49 10 00 5A 06 DB F6 F3 5A 47 DA 94 E0 29 18
 11 44 EC 61 DE C2 3C 18 74 C1 3C 61 84 AB 02 98
 D0 49 1A D5 E9 AE 4E C9 E4 21 71 FE D4 5B 4D 70
 E4 79 53 C6 DF D4 BD 71 CD D6 0C 62 5E 7A 53 DB
 88 A3 31 8C 5D A3 FF 22 CB 0A 57 B4 D5 26 33 10
 14 83 E8 F0 9E 4C 4F EB CB 1D 94 F9 13 DE 00 4F
 2B F4 08 BC DE C9 2E 3C 97 C2 AF 87 79 BC 3D F1
 30 E5 E8 59 2A E8 3D 34 88 B8 50 5C 2E 86 9A B5
 8E D4 E0 F5 ED C4 85 A1 D5 98 DE 67 BC 20 58 43
 3A 23 51 5F CA A3 6A 4C 58 6F DF ED 74 F5 16 F5
 E0 A8 35 A0 D9 76 63 81 7A 3F 05 9B 43 FD 9A F3
 21 6E AE 82 00 47 F4 55 38 99 56 CE 19 C7 32 E9
 A1 80 24 11 84 77 97 F5 64 C5 EC 0A C3 47 F2 F2
 0D F7 2E DE E1 59 9C 8F 10 A3 5A 16 5E 38 9B 5C
 38 32 48 B5 1A 9C B5 16 FC 7F 34 2F C2 0B 9D 21
 27 7C 78 B7 73 4D 0F 85 C9 F5 5D 3F 7F 75 88 C6
 29 F6 D5 84 B0 D8 2E 13 0B 18 10 ED AE B7 9F 4D
 39 26 C6 48 10 2C 86 C9 EC BD B0 D0 59 F1 60 1A
 B2 6F 21 26 9A F5 24 C2 75 A7 F8 28 89 41 59 B9
 C5 65 45 8E 82 B4 03 85 49 F9 69 25 86 C6 49 CB
 6A 33 B9 D5 A5 89 17 93 D7 61 7B 11 E9 53 6E BC
 71 94 30 D5 94 FC 31 53 8B 25 6B E4 12 3C 7E 82
 00 93 A3 1E 1D D6 3A D7 53 22 04 84 D5 BE 56 36
 1D E3 3C 25 0A DC A0 7C 1F 1C C5 87 FF E2 AE CA
 53 93 D1 8C 5C 9F AF 16 33 1A D4 E6 A5 AB 96 86
 F6 24 C9 E7 72 CE 8D 13 E1 91 0D FE 0B F5 31 53
 48 0C 7B 06 2E D0 10 35 D9 2A 17 93 50 E4 C6 C4
 69 94 28 63 92 A1 6B 7F 3A CD 13 1A 4C 61 2A 7D
 8B FE EB D5 0F 57 9F C1 53 29 C7 35 1E 26 B7 83
 13 1A 12 F2 0E B9 CF C0 8C 96 C7 4F A9 82 E8 2B
 B4 4F 8A 31 0E F6 BF EA AD 4E FD 07 F5 69 BE C9
 00 89 A5 04 F8 90 93 A5 E8 7A 34 4B B9 53 46 FB
 39 48 A5 59 37 BC E5 1C 06 87 EA AD 84 A2 EB 6C
 4A A3 DF 4C A7 F6 AB 70 FC E1 8F 9B 20 11 A7 37
 FF 6B E8 BA 85 58 60 AB 3F 30 0A AC 37 EF AD 6B
 21 8C B8 AA 21 90 5C FD A6 64 1A 45 22 78 C9 E0
 D0 22 AB F9 CB 85 01 22 97 14 E7 75 0D 16 50 23
 83 A1 FA 1D C8 D8 E3 37 C1 8C 36 16 9C DE 38 A6
 1C 76 C1 83 CA 37 5F C1 1C 9B 96 AC CA ED 64 72
 0A B1 4F DF 25 D6 27 E7 8E C6 14 B1 EF 0B 2B 63
 28 E0 65 C7 7E F5 4A C7 7B E4 EF C8 9A FF AA F0
 B9 8E 27 22 58 EA C8 82 BF 42 5A 14 15 C8 7F 13
 E3 06 43 96 45 32 97 10 F3 66 65 E5 C9 41 43 A7
 A9 C8 9A 0B 58 87 53 97 E3 DB 1E A0 6D 31 AB 47
 4F 0C 69 12 23 EC D2 EA 06 EB 5C A9 16 B9 46 74
 54 1D 43 BB 5A CB F6 21 73 F2 57 70 64 67 82 5A
 1E 2D 33 7C 52 71 D9 B4 32 E7 B5 08 F2 40 DA 06
 8D 29 A5 7C 3A 4B EE 72 DA 31 F3 EC 4E 52 F1 AA
 B7 4E 29 E7 7A 38 59 96 D9 FA 2D 96 70 E9 C9 8C
 36 D7 6A 9C 62 04 AF CB AE 69 FD 31 4B 29 A6 69
 8B E4 02 56 A9 0F C6 4F 3A 88 1F 5B A0 C6 CA EC
 AA 2B 6D EA 55 DA 92 C5 B9 C8 84 D6 ED AD 97 B1
 DB 08 F0 E7 AC 5C DB 1E 99 15 7E 39 45 CC 30 8E
 74 D0 14 E1 64 16 F7 A8 73 13 C0 F0 1E 81 66 85
 4E 62 7A 32 5A 0B D5 EC 76 C9 30 DB 09 56 66 7A
 E9 7D 25 99 EA F8 1A 3E 05 91 2D F5 5B 2B 84 FC
 29 89 38 E0 74 AF 83 04 00 0D 7E 01 A0 8B CE 67
 D7 94 6F 8C C7 B9 6E B0 12 31 99 72 C6 4C 99 81
 B1 E8 BE 11 D7 F7 93 9B 3F 9C 22 A5 5B 99 4A 45
 D2 56 E7 B2 68 7C 83 F2 34 F4 B6 0F 90 A2 2D 50
 26 6F 39 25 AC 82 FB 0E A5 BF 35 1A 6D 4F ED 9B
 C6 D4 EB EE CE 87 E2 55 E0 81 E7 1E 4E A8 52 C2
 AA 09 A9 2D 63 71 40 D0 A9 88 EE D5 FB 32 DE 47
 73 F8 21 18 12 A9 B0 A1 6B A9 09 FD 8F 9E 40 08
 BB 96 3E 65 F1 32 D3 8E 3B 2F 6B 70 D8 A2 8C AF
 E2 B1 5C 68 B7 F4 DB 3E 0B 00 C1 37 00 F8 3C 94
 34 AE C6 C6 61 CB E4 80 3D 95 9C F9 49 B1 09 99
 54 6B 01 42 6A DF 74 44 59 BB 31 89 51 70 11 BB
 49 6C 50 4D A8 0E 49 4E CE 65 BF 80 B4 CC 93 2C
 EC 05 51 C9 8D C1 08 C4 19 BE 4A 28 15 B4 42 D3
 6D F8 54 C2 B5 A6 0A E8 30 24 0E D0 C0 02 08 83
 D8 EB 6A C6 12 C3 92 5D C9 6A 0D 8C AA BF 6C 70
 79 6E 7F 35 09 58 98 BF EE C7 60 A1 13 40 3A D2
 DE 24 00 07 45 3A 02 FF A0 C1 B1 57 F1 29 E3 88
 F1 DB 0A 14 61 5B 39 64 EE EF 6E AC 4D CC 3E 58
 85 0D 98 D3 2A 53 78 F8 65 B3 20 FE 15 8F 8F A9
 08 15 B2 72 E8 4E 2E C6 02 A4 89 4D 7D 86 8C 86
 14 6B AF FB 5A 02 E2 BA 22 71 C3 CF 34 15 76 64
 25 57 6F 95 17 9F 0C 50 D5 C0 28 FF 6C 17 4C 8F
 11 02 83 66 4C 2D 06 9D 7B C3 62 E6 2E 34 00 C5
 63 1C 0A BB F4 22 EC FC 84 22 72 98 83 A6 E5 B3
 76 0E F9 3D DC A3 94 E7 95 B9 A6 8D 78 5B E7 72
 00 8D B1 D6 17 65 FA EF 59 A8 E8 95 49 E7 9A D4
 BA AB 9D C0 7E 42 B5 E1 A3 07 33 8D 3E C0 FE 85
 48 00 F4 60 5D DE FC F4 1C 47 0B 3E 13 2B 4C 29
 04 5A 1F AC AF 47 11 A8 CE D3 BB 3C 92 B4 CE 14
 08 53 04 7A 4E 79 7F 33 A8 65 8A ED 7B 2D 37 AF
 B7 6A 6D 10 97 7F 55 8E 84 36 9E 45 26 C2 82 52
 8D 51 AF 4E 59 15 FC 3F 8E D0 AB AB 2B 91 D7 A6
 F0 A1 6E 71 7F D7 8D EA 56 77 99 9B 40 EA 7C 50
 CA A8 EF 20 A0 3B 46 62 DA 6E C8 45 BC 37 B6 6F
 E5 B1 E1 82 DB 76 58 29 33 57 87 9A 43 67 57 9E
 64 F0 24 3F D5 98 A4 63 68 B8 98 AA 72 BA C2 20
 E5 01 E2 99 85 E5 06 A9 53 CC 96 72 C7 7E 12 CC
 C4 11 F5 33 C9 8E 10 AE 2D 13 7A 85 3B 6A 97 4D
 08 6C 0F CD 7C 2B 75 EA 75 23 7E FD 02 DA B9 D1
 53 E3 A8 95 48 2B C8 E9 02 E5 5E 26 46 B9 F9 7D
 5B 38 1F EE EA 5B E5 D9 48 A5 71 9E 43 BF F2 4B
 58 4E 94 04 B4 5B BC 2C 31 2F 46 58 D7 F5 DA 2A
 9F CE 24 D7 33 4F BC 48 49 BB 60 04 44 83 3F C4
 74 11 AE D4 30 FB 71 6F CD C9 E1 59 B5 AC 33 FD
 39 78 E1 58 29 92 92 71 7D 06 31 54 1A 6F A8 E4
 F2 A6 C0 0A 61 80 FC B8 52 5F 03 15 5E AA 84 0D
 D1 59 E5 DE 07 2B 01 21 C0 3B 77 AC AE DA F8 12
 7D D8 D2 79 A5 6D 3F F3 60 0A E0 8F A3 92 46 CE
 7F DE 39 4D 2C D5 29 2F 31 23 07 F8 4E C8 1C F5
 5E 13 6E 50 BD FF 72 63 DF 4F F9 88 13 70 A4 0B
 C0 31 10 C2 3A EB 53 18 76 FF 8D 29 80 4B 38 35
 76 A3 4A CA 22 6C 8D B0 52 8C F6 43 00 94 B6 48
 BF 31 7B F4 E6 20 C4 D2 CC 99 0F C4 93 0C 23 EB
 C5 73 BF 26 34 51 FA A4 30 42 E7 BA C4 DC 66 00
 78 40 17 1E 86 65 3F E3 92 6E C6 11 B5 98 C1 BA
 36 A8 2C A4 75 D1 65 50 55 47 AE 7F 94 0E D2 D0
 82 AA 51 A1 0E C3 4D FF 58 CA 2D 7F 63 14 1D 0C
 90 5D ED 25 5C 54 C1 32 26 60 A3 1D 11 21 23 7C
 97 BF 5A 56 68 02 8F 40 F2 FC 40 46 FF E0 E9 3E
 D6 DC D5 A3 7F 62 47 CB 0D 3C 64 8E 7B CD D1 E8
 AB 59 9D 82 AB 37 28 A8 89 97 EA 65 C4 50 58 C2
 BB 0B C4 55 52 C8 2D 94 67 6A A5 03 A2 86 C8 75
 F1 32 B3 25 18 94 56 44 07 C9 05 6B C1 0F AE 6D
 71 84 3D 11 F1 FD 64 1D 2D C8 A9 B9 83 BE 9A 24
 0C 8B 64 23 62 EF E5 E1 BE EB 99 D6 44 8B D2 92
 49 58 34 37 E6 2E 5B 40 F1 69 95 17 4A F2 60 CB
 4C 0A 17 88 BD 3D C1 57 D7 1B 51 E4 68 86 14 7E
 3C AE 88 F3 BA F2 B5 61 02 D5 E7 6E B4 64 B1 AA
 D6 11 E8 B1 D1 2D 7D FD 3A DB 5C 1E 2A 7D 17 1C
 C9 B2 B1 73 41 A4 3E F9 95 7A 9F A1 EA F7 FE D3
 9E D4 F1 2F 05 26 1B FA 35 CF 63 8A 0B 1C 7F 40
 43 6F 35 22 A6 74 92 E1 BE F5 E8 85 B9 CE 38 2F
 40 EA 6A 7C A8 79 CF B4 87 C4 43 0B A9 7B 9E 00
 83 DF 19 EC 1F 5E 78 04 1C B5 C9 56 7D 93 2C D0
 B5 2B F0 AD B3 4F C9 38 0D 41 94 C0 E9 46 70 C9
 DE C3 25 42 77 5A 53 3F 3C F5 F8 50 0B B8 72 5A
 4C DC FE 6B 0D 6A 09 99 4B 95 FF 45 BB 99 EE A1
 EB 7D CB A5 EC 74 E0 A5 31 A9 2C 07 72 10 77 1B
 D3 7D 3C B2 F3 51 68 AD 1B 4D 35 B3 20 92 84 E2
 13 B3 D4 A6 B9 A0 EC 68 5C 41 1E F2 38 7A 7C CA
 02 0D 87 81 17 54 AF 5C C3 39 DF 76 03 4F A1 5E
 88 97 0A E3 66 0D F2 F3 7A 69 1F 87 76 7B E2 8C
 78 D9 57 64 89 28 EA 72 44 F4 B8 D6 9F 9F 4A C7
 E0 B4 B7 D0 51 3B B7 C7 B7 65 C3 24 AE 70 DD 63
 F9 CD 15 5F 7B 87 59 A2 9D A6 88 BF B1 2F AA D9
 B1 3B 46 C5 51 15 00 BD AA BD B8 AF C7 85 ED B4
 7D 78 55 3D CC 94 6F 1E 15 3A C3 1E E2 E5 E5 31
 16 45 13 13 71 B9 81 DE 19 E6 C6 C7 D1 18 D0 F1
 BB 53 85 35 4A A4 FC EE 21 14 39 0F C1 FF 88 E7
 E9 BF 1B E5 C7 25 5A 56 B1 88 2B 59 CD 42 1D E1
 ED 35 F9 61 50 CF A6 43 B4 0F E4 88 65 73 2E BB
 46 CE 71 01 D3 72 18 9B 54 00 91 E5 7B 15 E0 23
 D1 39 18 25 DC 44 E2 C5 19 19 54 E5 E6 E5 0A D1
 8A F5 72 78 B4 CD 7F D1 08 27 F4 8E 5E C3 F7 89
 D3 5E 38 DB 40 33 8E 06 15 EA 63 3B 65 15 66 17
 68 53 43 42 CB 7A 28 2E 75 14 5E EA 31 2C BE BA
 5B C4 F3 93 24 12 92 F9 F3 10 71 BC B2 A5 95 71
 4B F7 20 1A F2 45 0B 77 F8 E6 01 6F 8F 29 A6 17
 80 41 53 D1 F5 A6 6D 90 B8 E4 79 60 64 33 43 B6
 E9 E5 65 1E 6A 1A C1 08 37 1B 79 34 56 F2 5F 6D
 9F 8C A4 7B D8 43 C4 4A A6 08 13 36 94 4E F6 65
 C2 16 16 93 EE E1 BA 1A 96 97 2D A5 55 55 23 86
 B8 6F 1B 28 2C DB F9 11 D3 A1 34 6D A7 AA 6A 53
 85 48 F8 5F 91 BA 4B 58 90 75 CB 5B 42 39 94 46
 40 4F 7E 06 46 86 79 AE 33 43 DD 5B C7 3C 36 ED
 0B 74 50 BC FF 5B AC 6E 3C B4 53 51 E4 0B 9D 48
 ED 8D 0D 82 F5 6D 11 A5 71 BF 35 57 27 BC 3A A3
 E1 AE 53 B1 CA 8A F2 B9 4B DA B0 C0 88 D3 E7 AB
 57 04 ED 94 B6 3E CA 66 57 D7 EE 75 08 EC 90 18
 CC 62 C2 58 AD 85 03 02 23 21 50 FF FD 6F 15 C4
 0F 5B 02 D0 53 39 4C EF C2 F6 0B 2B 3A 32 76 64
 9B CD F8 D1 62 61 2B D9 1A 41 1C 98 3E 8E 72 7C
 68 96 50 A3 3A 82 71 48 DC 1D 00 10 BD F1 0C 18
 7C 15 68 A6 38 48 12 44 8F E4 D9 14 2E 05 70 DE
 17 F2 24 69 A3 06 28 6F 52 E7 B4 CC 30 24 41 C7
 6F F0 BF EF 44 FD 5B 2A B8 3D 43 90 49 63 F0 5A
 FA AC C6 93 2C BF 80 7F 3D 8C 8D 9E 64 0B 58 DE
 9F B2 BD A8 FE BE 21 27 CF 4E B6 BD 36 59 27 A1
 0E AF B2 3D 42 BF DE 74 A2 94 A9 50 FE 83 7B E2
 31 94 AF 73 36 AB EA 58 F3 04 0F 1C A8 3B 7E 46
 E1 C0 74 12 07 DA E6 F1 5E F3 9B D0 26 A9 04 A8
 EA D1 61 2B A1 D0 77 EA FA F3 6B DE B4 12 18 94
 0A 1E 56 63 BD E5 09 53 03 3B 71 00 7C 79 84 57
 9E 08 65 36 12 7A B0 7E 02 F7 1C 40 CB 97 76 08
 B7 73 94 C6 00 B7 B1 59 93 C3 37 75 E7 2F 75 91
 74 BC 28 8A 57 3F 48 C0 54 B5 5F B5 3F DD 6B 2A
 C3 F6 24 47 9A 0F 6E 25 37 D1 25 EB 3C 93 05 96
 B2 54 4A 0B DF 42 CF B6 1C 37 82 45 DD 77 1B E5
 57 82 76 6B 50 BD D2 AF 31 83 D6 72 30 A5 2A A7
 6F 5C DB BC 82 9D 24 AD 33 93 A9 D9 3F 38 54 74
 EE B4 A9 9B 66 3F D4 99 26 7B FF 71 3C F9 44 68
 39 6A 07 3B B8 72 7A 16 18 2C 2E 9C 98 3F 41 7D
 85 D0 45 94 93 5C 02 48 0C 18 90 7C CE C7 67 6B
 73 C7 CE C4 60 B8 B6 7F 11 7F 68 94 33 21 FE 34
 17 0E 10 79 E8 1E 65 7E C6 1D 18 BB A9 EF 98 7F
 D6 23 C7 5B AF C0 05 0E D7 BC 5E D3 EB 0B CD D4
 5C B1 46 1D 17 3F 38 E8 B9 71 3F 4D 0F 9F 4D 4F
 99 62 36 C7 1F 6C 37 C8 9B 09 8E 92 AB BE 08 52
 42 FC EE 8F F3 12 4D 8F A5 41 79 BA 9D C2 D9 8E
 63 84 4B D6 01 84 23 17 F1 A4 87 AE CF 89 07 C7
 4E ED 6C 76 6C 5E 10 AB A0 A3 73 32 CC 0F 95 66
 B2 39 26 63 E3 27 9B 00 19 1F D5 08 D0 C6 F4 84
 DB 13 80 26 8B A7 D8 B1 BF F2 2A 34 8B AB 00 11
 54 3C A0 35 18 21 49 06 75 BC 7D 4D 1A 7F FB 04
 5E D4 18 E4 02 D2 0A 2E 5F 59 E1 B5 95 A3 AE 8C
 02 B0 E3 52 B8 45 58 3C 93 45 B5 BB B4 2E 38 CD
 7F CD 81 A7 72 52 AA CE 94 68 EA C6 F0 9E CA 5E
 85 83 5B B7 46 22 CC 98 EB 84 67 EC FA 36 4D 04
 77 D7 B5 8C 8D A2 7D F6 D8 F6 D7 1E D4 C1 C3 4F
 3B 35 69 14 3D B2 38 CA 12 09 B9 9A 0E A2 62 C8
 FB 0A 40 FD BB C0 BB 8F AD D7 36 B8 B1 A0 94 28
 7F 34 E7 40 D1 E2 5E C0 AD 9F 5A E2 E5 D3 80 CB
 C5 3B 7A 9C FC 29 A8 55 A4 AE D8 E6 49 5B BB 90
 0B 0F 7D BC 47 C9 84 64 61 C9 07 9D D3 04 78 00
 58 70 51 A9 4E 36 91 94 84 5E 46 0F 8F 7F B8 5A
 F7 4F BA 18 40 DC 79 8E DB 9A D6 81 AD 11 E0 6F
 71 43 D3 DC C4 01 26 D9 CC 46 6E 42 CA 6D 69 B7
 9B 66 04 5B 39 C5 01 20 C8 A6 8B 2C 71 84 5E AD
 49 5C B2 6C 35 D7 59 B0 66 87 D6 37 59 83 2A 78
 39 25 61 4D 7B 88 CC 4B EC 96 8F 37 E0 63 BF 86
 64 DE 2F 70 93 FA 4C E9 CA 72 30 47 24 B9 86 5A
 C8 42 3C 7D CC C5 94 EE 4F 79 20 A0 8A BD 7D 77
 A8 BC F7 AD 4D 13 0D 02 DB E0 9D 8F EC 65 DD 5E
 1B 3C 40 A3 EB A3 A9 EF 58 1F 8E 20 E7 ED C3 D0
 09 07 39 90 33 79 92 FB 37 72 F7 EF 8B F0 65 9F
 51 A8 A2 D8 81 98 7B EE 68 67 CA 77 AA 99 69 5D
 D3 0E A4 50 FE 7A 6C F4 A5 0C 50 BF 3A 67 73 DC
 2C 61 F5 82 59 10 71 F3 78 8C 43 E5 69 42 CD CB
 39 B5 C2 49 58 8A AF E9 E5 E6 65 13 B1 09 55 32
 67 70 04 9F 1A 2A FD 48 83 0A EA 76 AB EA E1 5C
 1A 9C 13 AC C1 FD 02 9F B4 1A EC C3 3F 92 81 9E
 1C 67 EB 41 36 2D 44 A9 7A B9 25 08 86 AC 41 ED
 46 F0 E8 F3 3A E7 D4 82 21 C4 BB 1E 5D 90 1F F8
 22 60 17 CE AA 35 EF 2D 16 F0 0B 04 5D AB 68 A9
 F1 00 82 11 49 56 77 A2 D1 82 FD 8E 6B EE 83 19
 16 C6 0D 57 EA A3 10 88 D0 FA A0 6F E3 D3 69 79
 FA 72 E4 00 C7 EB 1F A2 DB B9 46 6A BB 41 40 5E
 C6 55 97 52 3F 5C 5F BB DE C5 57 14 38 6E 37 B6
 77 06 90 7E E0 3D B7 19 A4 15 8A 2D 51 29 87 FF
 9E 78 F9 44 7C 45 D2 DE 2A C8 94 2C C6 24 75 E2
 85 B0 A4 09 B6 89 1F FC 4C 0D 57 4C 22 E4 CC E4
 34 F9 A4 06 D4 62 51 1E 24 FE 00 74 59 B2 D3 93
 C6 A3 BC A5 77 45 B0 A1 32 71 68 91 87 C3 95 18
 15 74 37 4E A0 06 4B C9 AE AC FB 4D 5B 07 21 5A
 D1 9C E1 16 B4 6D E9 F4 E9 B4 75 F8 0A C7 82 28
 20 CE 18 E6 72 29 A6 97 8E F1 2D C0 C3 F1 9D 36
 A3 CE 84 F3 4E 96 29 E8 9C BD 95 08 C2 D6 2E 40
 03 4E DA A5 3A 53 A6 33 EE D3 74 19 4C 2E 1B C5
 9F 51 44 07 BF C0 A6 C9 0D 6A 7B D1 51 4F 25 74
 10 26 01 1D FF BA AB 19 11 9A FC 6D 6B E9 17 6F
 EE 88 A7 3E BE 38 D5 17 3C 77 2D 9D E2 D2 C6 8D
 AA 67 F4 2F 1D 90 5F 12 26 5B DE 5A 5B 1E 96 B2
 EE 40 1D 93 20 50 3F F4 C6 23 E7 92 BF 30 03 14
 01 7D 7D 92 CF F9 02 D8 64 A3 A6 B4 90 D1 C7 DC
 8F 89 E8 4F D4 19 7D A6 05 8A A0 89 E7 89 95 95
 9F 39 54 79 1D 54 0A CB 2A C1 5A 1E F4 F9 FC FA
 3E 91 2D FD 4D 09 7F 09 27 47 5B 75 88 9C E3 ED
 19 23 39 1A C3 38 9A A8 91 4C 6C 84 C1 94 1E 54
 E5 0F 1C 54 AD 75 5D 48 00 CB 72 77 93 85 97 E9
 70 BC 7A C2 34 84 81 01 C4 5D 89 8E AD 81 EA 73
 4F 7E 60 F0 29 6E 9F 4A 7D FD BC 6B E8 64 97 C8
 D3 2D B4 2D 84 95 7E 57 A1 7E B1 92 09 17 55 69
 5F EF 95 1A 94 77 7A E5 06 7A 9C 42 4F 42 BA E1
 CA 83 5F 8B 0E D0 1A 0D 3B FE 11 0F 5B 31 A8 33
 C7 92 74 B8 E4 98 79 D0 AE 13 23 08 7D 55 21 75
 69 99 67 C4 E9 DD AF 0B 70 96 82 11 CE 0B 06 9C
 1F AD 71 ED 69 2D BE BC 5E 1D 9E CC DC 18 65 D8
 97 E4 C6 17 A0 04 89 B1 8B E8 4E 2D 62 3A C9 83
 A9 AF 6A 25 1D 95 1D 4C E7 A1 69 86 77 17 D2 DB
 97 AB CD 85 D8 70 09 37 CE E5 E3 47 F5 A0 1F F2
 0A A8 3F 3D 67 4C 36 E7 2C 72 21 33 40 98 ED 41
 C6 4A CC 45 7F 84 6B F4 FB 92 C3 4E 38 F6 97 48
 89 64 61 65 E0 40 25 BA 86 03 EA B8 5C DD B3 8B
 96 4F A4 30 20 9D 8F E5 44 95 DF 92 86 84 38 B4
 88 A3 C6 39 A9 CD F4 E2 B6 58 2D 4F 7E 16 B2 E4
 3C C6 96 E2 23 88 81 8D 0A E8 8C DD 51 4B 89 BD
 DC 59 D7 C5 A6 E7 3B C2 0B EC 7D 65 80 63 B0 22
 09 61 8B 7E 66 EA 39 F4 C8 4C 4A 10 F0 16 F0 35
 9B 53 EA 4D 69 77 16 BF D9 4B FF 0B 01 01 23 B3
 E7 BB C7 73 01 55 74 87 DE 01 93 2C A9 EE 9C D2
 F4 36 24 EA 25 DF 73 F0 FD D7 BC 7C 79 B5 96 76
 A6 62 64 70 33 E8 CD D6 D3 38 D5 5E EB 41 F7 3D
 EE A0 72 11 37 94 14 7B 2E CE 7E B4 34 7F 24 8C
 1B ED 02 22 96 2C D3 78 3E 80 71 D2 4F 25 B0 64
 6B 23 46 80 D0 C5 AE 66 4D 3C 41 29 3F FF ED 23
 54 E5 54 65 6B 29 19 F8 F1 72 80 80 A8 F0 C2 8A
 76 D3 92 13 8A 56 C2 B4 FB 42 42 3F 05 37 25 FB
 F9 2F 71 F5 E9 20 73 DD 0D 56 B5 43 40 23 B6 42
 F9 86 BF E1 E1 C9 9E 7B FB C2 0E 4F 6E 3D FA C3
 DC 6E 50 26 DB 1C 5B 3B 75 99 EB 1E A2 3C 45 87
 9A 53 05 A1 22 31 A8 B3 F0 36 6C A0 C4 7F 26 98
 35 D7 B5 0E 4D 95 63 BD FB A2 5B 05 85 50 E8 25
 D3 3F 0B 44 23 96 04 51 8C 99 09 5F 9B B9 93 CA
 75 4B 55 DB 03 51 28 82 47 D9 61 77 0D F2 4F 0B
 CB 10 F9 0E 5E 15 EB B2 42 F4 FD 92 41 97 C4 92
 20 5D 89 9B 16 75 7B 91 71 11 A3 44 80 F9 BA AB
 5A E1 0E FC 0E AC 3A C9 5B 5F 66 27 97 60 39 F2
 0F 4A 45 D2 C8 29 30 A3 5B A7 77 C5 29 AD CE 44
 5C E5 CD D3 CD 33 8C 34 CA B5 73 6E 54 4C EF 0E
 36 BC 80 11 1F 1F 58 10 56 2A A4 90 59 DD 4A 19
 18 51 9A FB 49 4F C3 A7 F9 CE 98 FF D3 DA 6E BE
 3F 34 49 55 A5 B1 62 34 F7 E5 18 CB AD 90 C3 33
 D7 BB ED 63 11 97 B1 F7 69 EF EE F1 1D 1F 85 B8
 82 9A C0 63 C6 4D AB 76 56 0E E2 F6 78 C4 31 42
 B8 FD 11 AA 18 AD 0D CF 33 B7 C9 D1 1B 4E 7C D1
 90 3F CF C9 29 C7 FF E6 13 5C EE 96 19 40 E5 40
 EF BF 5C F1 F1 08 35 67 F8 F9 B1 05 9C BB E2 00
 A7 35 52 44 B2 AB 20 2F 44 EC E4 A0 3E 61 F4 7A
 48 7F B3 D5 1B 27 CF 98 67 04 2D DC 71 DB 73 B0
 67 F9 10 EA 9E 3C 6C A0 D3 F6 39 84 B6 E7 A1 82
 86 D7 C8 FC A2 16 41 18 79 96 AC 71 65 83 57 25
 F7 D4 FA AF 64 F9 A5 F3 C2 6C B6 E0 4A FB EF 93
 A8 1D A8 20 A6 28 32 D9 34 07 58 1E EC DB 2C 80
 7C 20 22 92 29 FF 46 29 31 0B DC 9B E2 C9 B8 B0
 C2 38 86 4B 9A 5D 41 85 E5 3E 1D E1 C1 0B 4B 23
 A5 CB DF EA 98 A5 CC A4 A4 9D 9C 32 6A 2E 3E DA
 65 D2 20 89 15 B8 1B 3A 8E 8F 15 6F 72 3C 55 0B
 51 BE F8 87 49 11 16 F3 7A 9A 3B 87 DA 66 9D F3
 55 88 9A 87 A3 BD 3D 87 1E 8E 95 38 65 4C 94 5E
 90 EC 11 54 8C 3E 8F 47 EE 7B 46 F9 7C E0 0F 56
 A5 05 CC 53 D3 77 0A C7 FF 43 C0 C4 48 D6 E0 21
 B1 59 45 F4 8B 89 A8 F9 18 06 28 42 70 65 7A 5F
 CA C4 52 E1 CD F2 CF 4C 8C AE F0 C4 18 F8 A4 8C
 15 E5 FA F6 50 FC 36 38 C2 FA F5 FD E4 40 DF 39
 77 5B CF 0C 6E 94 D1 68 AE EE 9D 3F C0 02 31 3E
 2F F8 AF CA 30 00 EA 76 03 C9 C3 F8 6C FF C3 F7
 C0 1A A2 12 E8 A9 E5 62 7B 4E 1A 9D A2 10 AE 69
 DA A4 BA DC 9A D2 2F 56 31 EA 76 E1 B6 79 F2 6C
 63 E9 ED F3 18 BB 27 80 F6 11 E2 44 6F C7 00 8E
 9D E9 46 59 9D EC 13 61 34 56 AD 1F F6 7E 9F 1C
 22 2C 4E 5B BE C6 3C E5 CF 6B DF 8C 08 CE C1 1F
 DA E0 89 E1 19 6A 2B D0 02 60 64 D5 5B 58 BA 56
 68 72 D8 5A AE F6 FC DD D6 95 99 B5 8A F3 4B 03
 37 CC C0 5F 59 81 6E 2F EC A6 C8 41 CC BA 5B 87
 D7 92 10 7F 7C FC 64 B7 CD C0 54 B3 12 6D 7D 30
 93 39 A9 A8 EF 3D F8 08 7E 33 F4 FD 2B 98 E3 2F
 F9 86 A1 06 A2 59 52 42 8F 36 D9 73 C3 F4 7C 8F
 F0 C7 56 4E 0B FC 15 EC 65 72 42 EE 50 C8 77 74
 A5 F0 09 E8 63 93 C4 49 3E 58 28 2F 66 57 E7 D1
 B4 DF D9 44 4B DB 3E 18 7A B9 11 B2 D9 04 9C 99
 5C 58 29 D1 6D 56 E3 EA 47 55 5E EE 83 27 7C C8
 CA 7C 1F 7D 8E FF A9 AA 3D B1 CE 50 EA C6 D7 4A
 3E DF 71 34 11 F6 FC 6D 0D EF 42 24 2E 57 E0 0F
 AF E8 76 FF 4B 96 A0 58 25 95 C0 43 F5 93 CC 52
 02 1A 00 78 7B 7B D5 53 69 E8 72 69 13 E5 30 73
 93 18 AE F4 D6 3A F8 C9 81 39 45 10 91 54 B1 87
 1B 38 E6 77 0D 0B 6B FA FE 70 17 6F 90 05 18 8E
 8F A3 79 55 22 5F 98 E5 8F 89 BB 43 02 C6 44 78
 66 B0 EE A3 FC A3 13 9E 6C 08 CD 8B 1A DA 63 C3
 92 62 FA A8 ED 55 B5 61 58 33 A0 4F 8B 46 63 A0
 74 04 CE 68 15 99 8A 14 18 18 B9 4F 0A 81 B8 38
 CA 7F CC C8 6C 3F E0 60 FE 1D D0 41 6E C0 5D 97
 0A 50 8A 21 DF 77 61 89 05 69 8E DD CB 91 F5 35
 53 17 F2 6D 65 41 70 AF FE 77 97 25 88 DD E6 59
 10 D6 D8 6A 05 AC D8 DC 43 10 8D 5C 87 B6 3A 38
 EA E3 A7 20 E9 AE 1F D3 90 B5 47 44 CF 55 EC 36
 5A 0C D8 4E 8E BE 5E CF 35 8B 76 C1 46 42 02 9D
 1D E8 AC 44 28 AA 5C E6 CE CC 2F CE AE EE 57 45
 3C 2A 1D 83 00 74 00 C9 FE 32 93 FF 58 1B AD 5E
 D7 CE D8 B9 45 AB 92 59 F7 8D 5E EF A4 97 8D A4
 C0 43 44 D2 06 F6 1A 0C 6B 70 0A 31 8D F4 06 D6
 EF 5C 8B EC E7 E1 CE BF C5 45 B5 70 B4 54 E4 99
 BE 02 10 CF 59 CF B0 49 20 EC 12 D3 8D C4 BA 8D
 5F 8C 35 1E 43 32 A4 D7 1C 3A A6 95 B8 8C 92 85
 9B 42 EC EB F7 E0 FE 09 0C FD F0 1A C9 53 23 1B
 96 7F 86 BE 16 D2 42 39 4D BF 39 12 9A B1 F8 A2
 20 2A A7 66 85 C5 43 B0 01 12 7A 6E 84 95 51 DE
 DE 57 AF C8 97 C5 14 5F 93 38 8F 79 40 FA 84 18
 F8 89 DB 20 E4 E3 54 07 C6 9E FD 78 AE B8 D5 0E
 00 19 8D 7A 27 51 8D 55 26 01 9D 8B BA 05 82 CF
 D9 7F 43 7A 7A 5F FF B8 80 27 28 0B 55 A1 F8 90
 5F 64 48 43 35 20 A0 B8 56 C9 D2 97 3F 7A DA CF
 F8 06 E7 3F 6B 36 25 94 E5 0D 5A 21 29 37 ED 69
 D1 4C AA 55 63 AA 53 8D ED E5 41 AC 5D 06 7E 44
 F0 BF 09 7B 86 FA 43 3F 87 B8 FB 28 D3 77 13 14
 0F A4 C3 50 2B 16 07 BC B9 EE 5C 23 BE 3E 34 D6
 08 B4 91 10 E4 91 13 D2 A6 13 4B 74 48 F3 20 ED
 8F 2A 82 E1 BF 93 9E CE 06 4B 4D DD 2C 67 20 87
 77 EB 1D A7 60 6A 73 A9 AA 09 4D 78 99 81 9F D9
 5F ED DF 73 FB 5B 0A F1 CC 4D 63 18 E2 8F 23 67
 82 AE D0 26 63 07 CC 37 C4 DD 51 5D E2 82 B2 E2
 5A 66 83 1E 8A FA D4 D7 B8 C5 DE 00 E0 95 67 58
 C9 94 5E 67 87 63 E9 56 18 27 CD 07 F5 D7 D3 72
 0C E4 21 1D 6C 43 12 A3 E8 A6 4F 71 7D 50 0F F8
 EE F0 B7 CD 64 1A 6D B8 96 74 7A EF DC 0D 7D B9
 04 B0 70 4E D2 D9 FD 16 E8 A3 D1 FB 68 23 DD 87
 79 1E 49 A5 E9 DE 61 CA 57 63 00 1F 7D 11 59 7D
 D7 1C 2D 36 7F AB E5 0E 9F 62 80 1E 28 94 96 37
 05 F9 5D 8D 56 FE 14 FB 08 06 46 89 AF 91 9A 32
 D7 0C 1D 99 24 D6 D9 FA 30 FB 22 5D 35 DE DA 28
 E3 0F 7A E3 20 80 E4 AE 4F C3 0E C2 D5 EC 36 0C
 F5 27 4C 38 10 78 3C BD 8D 14 EC 7F 0F 14 F4 A8
 C7 F7 B7 E1 68 D8 8F 9E B0 8D 13 1C 6B BD 72 05
 65 86 B4 74 06 CE DF 4D F9 3F 1B C2 D8 2A D0 F3
 63 AD 69 FB 07 2C 0A 7A 5A 66 7A 41 B9 68 12 FF
 35 2D 18 2F CA BB A6 D3 7C EE B0 62 4C 0B A0 3D
 D7 F3 2E 73 D9 C1 4D 4F 79 15 35 83 0E 90 A1 71
 F6 56 96 DF A2 6F 60 4E 04 F2 36 75 D5 AE C8 AD
 25 FA 8E CB FC B6 FB DF 46 64 7F A2 42 A3 E1 92
 EB 71 1D 64 9A 94 40 1B AD 1B 2E 62 41 EB CC C0
 98 E5 B4 00 8B 2C 7B 0B 70 2B 82 B4 16 E8 8C BE
 E2 F8 F0 16 16 5E 9E D8 7B 7E 08 F5 03 7F 06 21
 3F 65 A0 01 73 A3 B4 4A 25 27 0C FF CB D1 46 95
 09 ED 34 10 A8 D1 04 22 F1 B3 AA 47 FB 48 21 A9
 EA 9B A0 92 CA 29 65 A4 3C 44 4D F8 AB 0A 95 2B
 5A B7 83 0F 03 28 D1 32 E0 35 37 74 79 FC 4C D2
 9A 1C 01 86 8D 44 55 34 36 AC 5B 63 3C 04 77 88
 97 56 5F 93 0A 06 E8 24 50 89 83 07 33 6B EA C7
 32 8D BF 2C 9A C7 ED A4 31 9B FE E1 82 52 B8 9A
 6E BD AD 59 3F CF 5C 48 64 09 62 61 3B B0 2A 85
 28 9F 9B F4 CD 4D FD 63 EF BE 04 75 18 7F FE 67
 CE BB 9E CC DE C4 90 CE F0 50 24 C0 67 A2 11 4D
 18 2E 13 B4 E9 E4 9C 7F 1A 60 D0 33 D8 98 15 F9
 99 1B 29 F2 67 92 29 11 97 2B EE F3 ED D2 D3 42
 A4 0E DE 4C 6E C2 D8 5F 00 92 46 75 AD 05 FB 7D
 19 B1 C2 86 70 21 30 90 32 5D 52 BF 52 A1 98 CF
 D8 13 62 B1 95 B9 BC DD AB 66 6A 55 31 CC 9E 56
 C0 C7 24 61 4F 82 48 1F C6 F1 01 22 81 1F 40 67
 E6 A7 40 6C 12 8C 42 89 48 2A D4 6F 02 83 98 8C
 A0 D5 DC D1 2F E9 06 A4 28 2A DD 1C 68 D3 28 86
 FA 8A DB 02 42 7A 9F D3 87 C0 02 B5 BB 92 8F 15
 EC 39 BF C3 64 87 7A C2 93 D0 18 09 84 8A F4 AC
 BF 71 81 CC C2 DE 2C 94 E8 2E 9F 87 93 61 D2 1F
 84 11 35 A1 87 2A A0 54 93 4F 0E 30 B1 BC E9 80
 A2 4D EE 5C CD 73 98 0D 3D B8 0D 6E EB 98 03 9C
 EA 12 41 C3 93 94 05 D6 BA C8 8E 0A EC 31 E1 8A
 E7 71 09 03 77 09 C1 C9 D8 B1 92 54 43 21 2B 7E
 C7 E1 CF B3 F9 0B E8 07 B9 C4 50 DD 19 E9 2A 2C
 54 DC 85 46 45 41 90 4E 7B 57 C4 4A BF 44 9E FC
 D7 62 08 8E 12 59 0D DD 39 4B 8F 07 EC 76 DC 85
 88 D9 00 58 6A 3B 37 50 F0 E6 63 C3 1B 83 39 A9
 4D 7C BA 14 D3 F3 ED 69 16 CA 77 B4 AC C6 FB 1D
 75 C4 35 D3 C9 87 17 B9 B8 57 1A 63 2A 50 14 61
 F6 2A 89 B8 DC 53 5B 40 CB 04 6D B3 D7 D1 D4 3E
 F5 F2 B6 83 CE D6 D2 E4 20 D7 64 7D EA 62 E5 6E
 85 74 C5 DF CF 4D 70 F4 01 5A 7C CA CC 82 1A 9D
 77 36 15 67 94 58 A3 9F 57 62 12 99 4E F3 AB 87
 B1 D2 B7 CC 53 92 36 98 04 41 3C B3 AC 77 89 F9
 E2 F5 84 EA 5B E7 B5 57 2F 20 40 EE 9A 69 30 5A
 30 41 66 35 47 58 B8 4F 5B DA D2 B6 4C E3 0C F0
 3E D0 94 8A 6C 84 5B 98 FF 1D E0 68 24 13 A0 69
 00 B1 55 CB 84 1E 05 0D B8 12 1C 7F 1F F8 13 87
 77 7F 2E 92 4C 2C 87 1A 93 69 B8 69 48 4F E6 77
 A1 FB 0F 10 03 13 87 56 B3 1D D5 F3 4A 35 AB 72
 3F 00 4E F2 87 8D 95 3E 2B 5D 7D D4 C0 53 E4 4D
 3D 46 B8 5F 44 81 2D 3C B6 F6 B1 22 A4 7D 03 E4
 E6 07 6A C0 1D D3 F2 16 07 F0 93 5A 78 64 11 BC
 20 B3 31 55 C4 44 7C BC 36 38 8F 60 DC AF 79 08
 2A 45 0D DE 13 F7 1B A4 05 A7 13 63 97 1B 4C E8
 80 9E 8C 72 82 21 CC A4 D1 C0 63 FC 98 25 C1 26
 86 BA 34 63 B2 86 2B DE 8F 01 9F 45 39 E1 11 2D
 A7 41 FD 13 F7 F2 25 63 DF 86 4F 1C D2 00 EB 87
 7B A2 E0 74 CB 2A 08 C9 D1 C2 21 4F AE 95 BD 89
 39 92 5F EB EC DE 28 CE B1 52 7F F7 9D 03 9B 37
 AA 36 D1 6A 93 B3 AC 30 3E 5E 1F 89 4F 28 33 02
 1D 6D 13 EC 36 67 0B 82 44 DE 7B A9 84 6B 85 33
 DC 1B 01 42 4C DA E5 D2 92 A2 54 8E 81 3A D1 88
 21 6F 53 9F 5C 25 D4 89 2D 39 00 CD 31 3A 2F F0
 67 F3 0D 94 48 FF 9C 34 A9 29 7E 39 74 DF 81 8E
 0F 9A 67 63 C3 15 4B 24 48 5F 10 FC DC A2 ED BA
 C9 09 28 A2 D0 54 63 A3 10 A4 B5 67 95 B7 A5 1C
 1D 3A 95 D5 2B 15 96 84 67 51 A7 0B 02 B0 DF F5
 2C 03 35 86 E8 37 14 8B 57 04 D3 0E 85 A7 0F E2
 C0 E9 1A 06 8D 52 CA C0 FF 78 B8 35 01 73 86 EA
 E9 83 28 F7 D3 9C 0C 69 00 E1 A1 7D DB 16 36 4E
 8E 0E 9B C7 F1 53 AD E4 E0 05 E2 47 CD 4D 42 18
 D9 69 82 E2 EA C3 CB 50 4D C7 DB E7 B6 45 1F EC
 C4 0F B7 49 E1 08 C9 17 DE 3B 48 97 15 92 49 3E
 98 65 2D CE 10 87 25 2F EE C1 51 2E AD 49 FE CF
 33 1D 52 AB 1A 6C 67 2F 96 59 07 1B F1 CB 51 93
 26 6F CB B5 00 79 A1 9C 98 73 1F CE 13 CA 92 F6
 B0 E5 89 30 A1 7B 1F 44 6B 0B D4 04 F2 36 FE D3
 D3 EC C9 95 01 DF 62 2E 08 F8 8E 04 11 4B 51 7F
 40 9E B6 0B 93 39 60 F4 62 FB 7C 15 BC BF 2F DE
 54 CB CB B5 3A 91 CE 81 0E 34 6F A5 37 B6 DE FC
 2B CF F3 EE DB F0 B6 64 C5 F1 8B E5 54 A6 0D 7C
 A6 29 D2 85 55 CB F4 8A 63 02 DF AB D8 4E A7 AF
 EF 68 D2 F1 09 1F 49 DA F9 88 9C 33 EB 5E 46 A9
 1B 95 AC 9D A3 DE 29 AF FA CE 0F 41 A5 91 81 88
 E1 90 7F 46 6F C7 A9 20 C2 07 C7 94 A2 6A F4 5A
 9F C3 B8 58 E8 D4 17 6E 8B DB 14 FD 7E 76 86 09
 73 4F CB D3 C0 E3 E8 9D F7 92 E5 5A 8D B9 6C 61
 AC F9 9E 25 6C 3C 49 5A 55 A4 9E 70 41 78 9C 0E
 DE 3E 82 69 B3 80 85 22 65 5A 93 C5 9E A0 98 E7
 4F BE E4 28 85 B5 72 AA 9C 69 F9 E3 75 F8 1F 5B
 EC 7F D8 8A 38 F2 51 79 FF 74 F0 A7 60 54 0D 98
 80 CB DC 7E 41 0F 7D D2 41 43 B7 88 57 1E E7 1F
 AB 1D FC C0 83 87 CB 9D 4D 6E 10 47 5B 11 21 24
 FA FC 02 C2 8D A6 6D AD 2C FE F5 E9 CF AE A4 29
 0D 00 21 C0 08 D1 01 3C C7 D5 36 6B 77 3A 2F E6
 41 8E 52 55 C5 DD DB A4 2D B0 A4 7F B6 F8 85 00
 0F 59 49 1D D3 67 E4 B5 89 73 9C EB 85 83 9D 70
 62 9B DE 25 69 1B 79 75 9D F2 F2 B9 52 10 51 7D
 59 50 14 6D E7 78 EA 91 7B 94 BA E0 EA 24 59 53
 38 D6 B4 C7 5F F3 C9 D0 DB 1E D4 DE 64 21 F4 F6
 2B D0 F0 57 E0 CD FB 10 D1 13 60 60 5D 96 34 D1
 31 60 1B 5F 35 40 7D D7 63 4F 36 B2 67 6B 01 2D
 34 03 E8 5A 15 4B 80 E8 48 00 F2 48 D7 21 DF 52
 E3 AD 4D 09 21 83 61 04 44 4A 1B 4E 6D 9D 6C 79
 3C C7 DB F2 C9 A9 F5 12 36 E3 97 86 A2 B0 A7 6D
 9F 3C 8C EC A2 F5 FB A3 A0 B9 93 BF 85 3D 29 1C
 33 7F 28 CA DF 83 01 A7 8E 63 A7 9E 5E 7B 60 3F
 1E 22 85 E4 E6 5E 97 30 46 1A 91 5C AF 7A 7E D6
 4B 40 75 6F 2F 75 15 49 A4 2C 4B EA AF F8 BB E5
 04 CA 46 4B 70 7A 9D B8 7F 2E DD CF 34 46 AA 96
 B7 BB 4E AA CB 9B 31 B0 B2 74 20 CA 77 B4 AC 41
 03 F0 A4 26 D5 E2 2F D5 8E C3 BB 34 55 F8 BC E0
 72 08 B2 74 EA 56 87 A6 9F 6E C5 69 B4 CE BE 9E
 82 73 D9 10 31 5C FC 4D 6D B8 7D E8 EE 88 45 32
 54 E9 3C B1 B0 CA 74 B9 2A B7 97 FC 5D B5 DA C3
 09 C6 E3 3D 52 86 DC 74 5B 1C 79 CF 1D 72 D9 BE
 04 14 61 23 B3 D1 16 07 9D EF 58 6F 20 4C 76 63
 F9 56 22 A9 C6 75 49 C7 E3 28 4B EE 53 EE F7 E3
 31 B1 06 7D 8F F5 28 F7 15 FE 83 C2 F2 B5 36 26
 D9 55 07 EF 1E DE EE E8 50 C8 C7 34 A5 0A E9 10
 85 32 28 28 65 F2 38 EC B2 C0 50 00 97 10 D8 98
 18 4B 22 E6 F1 E2 AD 3B 03 B3 D6 AD 68 BC 68 D4
 33 60 5B 57 F0 89 53 CF 56 E8 BB 4D E6 E5 CA 8E
 84 E1 8B 77 F0 F8 C1 05 A3 A0 C6 9B C3 1B 50 52
 79 4F 57 0A AD 2F AB F3 F3 9B 73 D1 C7 49 75 BB
 88 CD 2D CF 70 56 45 E9 DE 06 3D F6 E8 CA 0E 73
 5C 70 BB C4 7C CA 6E 7F AE CB 00 6A 48 75 9C D8
 FC D3 86 05 37 65 88 8D 88 DB 37 CC 44 2A 37 04
 1F D8 DF AC CC CB F9 72 58 2B 09 D9 40 BE 10 04
 4F 66 4F B2 EB BE 3F 8A 1D 32 35 12 46 B7 6B 64
 64 EB 1D E3 1D B3 19 30 74 4F 70 C6 27 DD 81 2F
 2C 96 F4 7E 52 15 57 A7 5D B9 75 00 0B 59 1B D6
 88 A5 80 93 2E D0 13 DC 37 96 87 97 76 44 36 9E
 64 48 DE A4 0F 2A 80 12 E8 1B CF B8 1C 8B FC 58
 20 36 F5 1E 57 08 D5 29 F1 D9 EB F0 CE 6E F9 49
 12 44 72 F5 85 18 1F 14 19 CB 12 AE 6E BD 09 AA
 9B 20 70 AF 23 B3 09 C2 6D 76 23 B6 2D 2B 53 6B
 3A 23 26 37 45 54 88 45 7E E7 34 30 C8 FD 47 DE
 9B 4F 31 84 3A 71 AB 83 29 4D 35 83 FB 46 FE 93
 7D 37 A8 2A F3 7E EF BC 9D DD 0B 1C B1 8A B6 36
 D2 1D FE 14 F2 37 06 18 EA B0 0C FF 19 78 63 0E
 7E 84 77 68 68 DD FE 78 93 43 AD A4 F7 BE 85 A1
 12 D1 CC BD A4 77 3B CC 48 52 47 D8 20 CC 21 0F
 14 07 69 DF E1 90 68 EF 9A AE D1 C5 34 A1 6F D6
 FB 74 F5 F8 4F B9 59 BE 41 64 98 7C F1 FF 95 60
 4F DC 79 23 8B 31 5E AE E0 2C 7B B0 D5 85 78 F8
 C8 E2 2D 85 2B 75 E1 53 EE C3 14 F6 63 76 60 55
 8B DE 50 08 A2 C8 02 35 25 48 49 4E F0 B4 8C DA
 8D F9 91 E0 9A BD D7 BB 13 10 32 32 54 AB 0A 5F
 A6 52 E4 DE AC C0 EA 24 F6 D6 8C 01 8F E4 A7 CE
 B7 BE 47 DD DB 8F 8A F0 BD 7F 99 31 0C A3 63 4D
 51 87 90 FB DF E7 67 60 E9 2E 94 06 2E 09 0B 8D
 C7 89 39 7C 8D 75 C7 9B 16 EA 3D 29 74 21 69 B1
 B6 89 9E CE 1D 7F 63 BF AC F4 6A 97 2D 51 E9 01
 41 08 BE 57 92 EC B9 24 54 B2 A4 94 09 FE 37 EF
 E0 46 65 2B 61 A7 18 AC 56 3B CF 25 B1 50 7F DC
 5D A4 F7 D7 8A 93 AA 01 FD 71 C5 B3 DF 41 35 24
 0F D9 04 C9 27 8B F9 7E 69 1C 5B E4 FC 2B BC 62
 B9 C3 3A 77 3F 28 FD 79 DF 0F 68 60 9B 26 E2 35
 F4 2F 4C 8B E8 3D E5 C0 11 02 5D 7A 8A BE 2A 2F
 27 9F C4 3E 51 78 4B A1 84 9A 54 5C F1 C5 FF F4
 A9 91 1B F1 94 9E 7D 71 89 C3 FC D0 2F 75 4A B8
 F0 21 EB AD B9 DA 6E EE 8F AC C2 10 46 05 E3 E7
 22 4B 76 4B C8 55 BB FF 63 33 F4 34 2A FD 1A E4
 5A B4 58 EC 6D 46 D6 D3 01 99 22 9B 87 F0 E4 D6
 A5 6A C5 A8 1D 66 A6 8E 21 88 83 62 EC 03 20 5B
 3A 27 41 DE CD 36 61 55 F9 76 49 D2 42 16 6A 8B
 A7 28 EE C8 E9 0B 7E 32 65 20 DE 40 02 86 AE F3
 B6 4A D1 5D A7 F0 61 B8 1D 9D ED 43 57 91 C9 37
 4F D6 DB 06 70 FB 73 89 02 EB 6C A4 6E 36 FC 68
 24 BF E2 AC B6 0E 55 44 CF B6 41 4C DB 77 AC A3
 4E 72 F4 4C 68 20 4B AD 59 2D 48 C1 52 8E A0 BC
 03 D5 C1 5B 6D 0C EC BC 9E 0E 74 DE 0F 27 88 81
 3F 8E 7F 85 E3 42 7A E9 65 4D 72 BB C9 25 59 F9
 72 19 FD D2 BA 57 F2 4D 58 AF 37 59 9D 89 1E AE
 C5 10 05 ED 81 3D 7B E2 8A 3A 19 48 97 0A AB 9A
 D3 56 32 EA DB 41 3C AE 79 1E 44 71 7F 89 4C 4B
 BD 76 16 12 29 D6 40 A0 A2 42 9F ED 96 70 9E 0E
 FE A7 D6 A4 87 93 45 FB 66 C3 E5 92 8C 73 9F 05
 93 59 45 7B 5E 07 7D 36 FF E6 41 CE D8 F9 4D A0
 D1 D2 52 3D 62 BD F7 C1 82 78 59 23 8F 2A 2B F1
 EC 18 0A 3C BB 8C AD 8D 21 2C AA 20 A7 5B 40 58
 70 C4 F1 74 A3 86 DB 30 3C DC B5 4B AC 35 A9 C7
 8D E8 4E 01 3E 69 FC B1 CE D0 4B 93 A8 4A 51 61
 35 DA 74 C1 C1 9C 7B 44 A8 E1 1F 88 AF D0 91 99
 86 5B F8 07 11 C2 AB 45 AB 89 81 C4 B7 EF 2D 28
 68 38 F2 53 53 54 07 03 1F EB F5 67 6A 87 45 B9
 98 28 82 DD 61 96 0A BA 4A CA D0 8B 1E 78 96 7C
 C5 54 A0 1A 91 DE FA 63 C5 0B 94 C4 98 9C C8 67
 2C 64 DB 4F AA AC 57 F7 06 F8 BA B3 21 89 8D E4
 48 FE 5B A7 13 D0 28 A0 CC D8 D9 6A 8E 96 8D 9B
 A8 AA 60 17 41 1B 39 C4 19 AA 8B 44 D3 30 CF 2B
 69 28 57 79 7F 1E 8E 13 BE 2A 19 C4 D5 82 77 66
 63 96 0E E6 26 BD 30 A8 AC 35 0B D0 EE 28 57 F2
 79 3D 30 F8 E1 3A AB C5 EA 12 51 1E 3D E7 76 62
 85 B9 53 FE D3 58 F9 F2 76 36 38 83 65 59 05 6D
 9F AE 17 75 3B 09 5F C9 4F 4B 1D 75 43 63 C7 34
 16 54 7A BE E6 75 61 BB EA 9D 68 6A AF 7D 06 F1
 5B 22 01 CE CE 87 B5 3B 88 20 DB 0B 82 A1 E4 1A
 48 46 23 94 55 65 90 08 8C 41 EE 8E 7E B0 A5 F1
 6A 38 0A F1 3D 2E 6A 8D 04 33 AC 87 65 18 B3 1E
 C8 80 C2 01 D6 70 2D A6 1B 4B E1 87 B9 1F 6D 4B
 FD 8C 89 D6 71 C8 A4 E0 20 A1 D9 80 DA 75 CF 10
 AB 3E 94 C9 4C CF 22 81 A7 A3 62 50 6A F3 02 1E
 07 21 9A 74 27 0F BF 57 8D B9 6D 0F 9E 22 B0 90
 8E 46 F0 19 2B 00 52 2A 28 5B D8 11 9F B5 A3 18
 FA C3 70 37 80 20 1F E6 90 8D 50 AD 22 4F 2C 35
 38 52 A2 41 07 87 8D D0 AB D5 23 17 69 17 5E 65
 11 C7 54 F7 E0 91 C7 F1 0A 05 43 B4 25 98 01 FA
 3A 78 8D B1 D2 C9 9A 68 9C 65 CE B3 7E 1E A4 C7
 CF 7E 90 AD 10 2F 8A 76 C0 B6 CE 26 C0 F6 32 DB
 C1 AF 88 FE 38 45 2C 6F 54 79 F5 CA DD 99 65 AD
 5D EC 5F FD FB 62 C7 A8 7E 91 79 B2 4D 55 68 70
 F2 EA 8E F4 90 20 F0 81 67 33 B0 EE 26 C7 32 54
 F3 05 94 92 13 1C 1B 8A 03 DD 54 F1 C0 48 DE A9
 0F 68 93 25 40 D3 66 1B 5F 6E 64 15 EC DF FA 24
 0A CA 84 61 13 B3 D8 F9 AB 1F BA 0C E4 4C 42 93
 68 04 80 B8 79 AD 82 B5 AF DE FC 0C 42 E1 18 35
 F0 11 50 39 6F 8D 9C A3 71 17 20 3F 7E E5 2F 4D
 16 AF A1 E7 08 4B 8D 11 63 68 CF 63 A0 5F 5D E6
 7E B8 39 4C 46 BE 58 4D 9E 38 80 A9 B6 9D AA FA
 7C ED D8 D9 6E 33 63 CF A3 7A E9 E9 B0 FC 31 40
 5A A1 D6 94 90 A8 C2 3E A7 A1 E0 0F 7A 96 05 5E
 ED 71 43 F5 DC 10 C3 DE 92 05 04 1A 4C 3A 6C 39
 F4 89 AE F0 60 CB AC 28 1B 7F AD CC 28 30 02 18
 BB E6 BB 42 20 7D D9 02 48 66 0A 15 04 AD 7C FD
 00 24 A9 DA B1 71 BA 9B 5F 30 3C DC 0F FA 07 3A
 C2 72 A9 23 3E E3 2A DD 38 B0 60 CF B8 6B 8B A0
 32 43 BE 1B 50 1A 8E 0D 22 5A 0B AD EC BF 79 6B
 0C B2 32 48 F8 E2 87 F3 0D 9B 61 AA 00 82 0B 48
 AD 1D 1F 23 30 A5 2C 4D F4 E0 CA 8B 04 DF 72 F6
 F5 E2 98 6B 1D 3A F3 BA CE EB 95 6A E0 C0 BF C8
 9C E4 AC 0E 1E CF CD A7 5B B8 34 91 99 1E CD E5
 00 BA 4F 1D 37 84 AC 0D 04 FF 72 33 91 B7 3C 4A
 F7 8D 87 16 20 AA 92 8B 37 A0 E7 0C 60 14 C5 0F
 C7 D3 0F F2 EC 77 7D FC D9 EB D0 F4 2D E4 5D 11
 59 C4 CA CE 8D C6 87 3E 86 5D CF 79 5D 92 23 0D
 E5 F2 AB 12 FC FE B3 A3 84 15 AC 50 AF 82 47 F9
 03 84 EE B0 F2 BC 57 6B D9 93 24 9A 4A 64 2B BA
 2A 7E 2A C9 7D 49 D0 56 D2 4C 7E 0C E1 CC BC 02
 75 AE E0 3C 2A A0 57 BC D3 C6 E0 06 B8 FF DB 34
 FB 36 43 F9 19 89 1E 18 71 E9 40 3C D2 E3 34 C4
 F4 40 14 CB A7 28 86 E8 4B A3 2B E5 5F 5B FB 6D
 2C C4 90 08 5B F3 A4 3F DC E8 10 78 38 14 E5 F0
 E0 F3 83 50 9E AC CC E1 4C 37 E9 F4 E8 78 18 06
 BA 93 9E EC D5 F1 EE 79 B2 C9 DF D4 01 22 9A 44
 C4 C2 3B 07 E2 2F 4D 00 8F AA 22 67 B4 90 DD 65
 06 1B 14 A1 8F 58 40 C9 1A 8B 5F C6 9A EA 85 35
 01 7B 19 51 32 2F 71 BF EA 4B 8A FC BC D1 08 02
 0C 04 EA D5 5E 82 65 AC 72 F1 E2 59 B2 C4 C1 14
 DC 7F 1E 5A 93 61 72 4A F9 E4 68 F3 7F 1F 98 74
 73 4B 15 10 AE A8 06 B8 DD 49 82 85 1F 4B 52 7D
 E2 D4 84 DA 60 12 87 87 48 35 7A E5 C5 62 11 3A
 5F 69 07 DA CB 8F 39 32 58 59 EF EC 47 B9 F9 73
 2E C8 C8 82 60 13 8A BD CB 66 45 33 EC 4C E6 7E
 E7 A0 25 B1 FC E5 35 5E 62 6F 8B EB B7 8F E2 86
 69 B5 8B 01 B2 3F 20 71 FA DA 44 60 D7 B2 8D 76
 6F 42 B5 33 16 3D 1E D2 98 07 FD 9E CD 3F 36 84
 49 7D D9 D9 D5 C8 DC A9 18 D5 61 36 A4 17 B3 55
 06 CD FB E8 6B BA E3 95 DC 77 21 D3 00 A1 02 FE
 F5 97 45 23 87 10 9B 71 E4 25 1C D6 1A 29 D3 DD
 D6 80 95 3F 1B F8 83 2B AD FF 95 C8 26 1E 70 83
 DB 54 02 C9 F2 0B A5 3C 56 29 48 DB 4F 60 80 4A
 51 55 BF 16 6D C6 E8 27 84 D1 8F 87 96 FE 67 49
 62 2B FE C8 82 4B 82 44 89 44 48 30 1B 93 8A A8
 BF C5 1E 4F 2B ED E7 4A 9E EF 2D 45 10 A0 91 AE
 C0 EE 07 77 35 73 F3 0A 4E 8D 75 A3 84 5D A6 B6
 32 40 51 DB 2B D6 90 17 EA 30 AE 40 01 70 2B CA
 BB 70 91 6A 0D 28 7D 5D A9 D4 F6 09 E1 A3 38 6A
 CC 67 D0 D0 66 B8 18 B8 90 17 B4 BC 4A 6E 05 49
 51 FE AD B3 9E 09 0E F1 39 D2 12 61 86 87 BC 61
 1A 73 AE BB BC 8D 56 A5 54 41 59 75 C1 B2 7F B4
 0F E2 C2 18 F7 1D 1E 07 9F 49 E9 91 EF 38 89 C6
 CD 84 7B 2C CA 56 73 50 46 42 93 1F 4D 33 15 C7
 D2 A1 64 FF D5 B2 C9 72 32 7B 42 70 D3 C5 E8 84
 1D AB C6 DC AA F4 37 10 0A 99 A1 89 D8 F5 7A 42
 7F 6D 9B E2 3B 56 56 62 F2 97 49 18 0B 78 A6 51
 E3 CC 1D B1 F6 19 AC 55 D4 37 8E E6 D0 F8 19 4B
 B6 D2 E3 0D 55 F9 8F 83 AC C0 07 CA 73 77 58 C6
 9A AB AB 91 49 A0 89 B3 C1 1F 4C F7 C9 09 85 58
 E6 6A 62 76 CE DC 38 DE BC 18 44 0A 11 9B EF BD
 CC C8 C3 A5 B5 92 79 E0 8F 35 C6 94 4A 4E C0 08
 AE E5 5A DF 06 D8 6F 07 2D 86 F6 8D 02 D1 8F DE
 1E 8D 1C 66 36 C2 B0 3F E3 47 F4 0D 26 16 1E CD
 50 6F A2 D7 C6 29 18 D6 25 3B 07 5A BA 12 9F BE
 EC 3C A6 74 84 28 A3 47 28 4D F2 AC 29 94 20 E8
 06 A0 43 E2 42 BB 0A 1F 95 31 02 3C 2A 22 4D 54
 C8 2D EA 4D A8 3A AC 3C E2 C5 AA 3B 74 1E AD 8B
 23 B9 AC 1C 75 25 A8 92 9E F7 D3 87 A4 6C E4 D4
 D6 F5 A2 0B 01 5F B4 A8 3C 5D 2C 0D 5E F6 F9 00
 7F 5E 1E 83 FA A6 83 0B 3F 34 16 51 5A CE 20 E0
 5B 6D E1 EE 06 EC 0A A0 C6 48 CA F5 B0 EB 05 2F
 69 E0 1E 93 28 BD 31 41 B0 95 E4 7A 2E A4 41 B5
 A0 FE C8 73 D3 3B 54 0A F3 50 BE 4F DF BF CB AE
 3E 57 E3 CC 7F CA 0C 72 F1 27 08 96 DE EF 8B E1
 E0 25 B0 AD A1 62 52 C9 9C BC 25 38 67 B6 DE 86
 C5 2F 0F C7 14 05 0F 5D 8F 2C 60 2F 08 3F 1B F0
 40 85 61 28 90 A8 B7 F3 A9 BA C5 3D 6D F4 05 DE
 57 88 A8 F7 C2 B7 EB BA 5C AB 1B A8 8C F7 9F 01
 99 DC 26 79 FF 4A 1A 54 07 EA 6F 3A 24 31 2A 3A
 FD 63 31 CB 4D 86 EB 00 C7 4D 27 D8 85 2F 9F FB
 AF 0B 4C 91 F8 80 C9 99 56 C3 95 57 EA A9 B7 49
 AB 90 8E F6 54 E0 DB E8 45 F1 38 56 E9 A3 0B F7
 A3 21 B6 56 BF 10 07 DB D8 CF 28 6C B9 EE 17 5A
 9F F7 A1 10 FB 27 7E 53 17 A8 9D 2C 2C 7D 16 50
 21 3A EC 71 DA A2 47 04 73 2D 58 89 3C 90 F9 C2
 1C 6C 68 F1 40 70 3C C1 11 60 00 8C 32 97 F9 2A
 CD DE 53 FB E9 96 63 8C A7 CA 06 51 AF AA 2F 29
 D6 58 4F 6F 5B 07 3D AD 03 CB 1F E9 C4 87 76 8D
 E0 3A 10 C4 C9 A4 61 A1 19 60 80 93 FC 15 64 45
 F2 2B 75 8F E8 95 F4 13 99 0F 38 92 BE 63 71 63
 A6 22 6F 5E 8E 3D D4 10 5B F0 0D 00 AD 7D FB 8B
 19 13 52 06 33 01 9A 77 75 44 5A A2 C7 DF 90 AE
 C8 4A 67 BE 30 1F 28 3B 6E 37 8E B6 4A 2F 89 81
 80 9D 1E 00 5B EF B4 07 5D C8 3F 69 83 C8 50 44
 07 9A 0C 88 F6 EC 7A 5A 4E AE 57 23 E4 A8 21 5E
 BD C5 C6 49 4E 9F D1 22 44 40 69 E5 22 49 EF B9
 D6 6D 38 DD 49 D7 D7 6E 17 46 0E 35 0D B8 61 FD
 0F C6 BB F8 C1 E7 54 C4 9E 3B 4F E5 B1 7A E2 51
 25 77 84 E7 0B 93 63 13 59 E8 85 FE 0A 7A 00 68
 F1 24 3F 7B 00 12 41 84 79 6F 51 05 81 CD EA 08
 1D 64 75 DF 12 39 28 FE 17 60 72 01 5C 6C 88 A5
 22 95 80 95 04 22 C7 F0 65 9C 4D E6 9B A4 B4 C0
 D4 2D A3 BB 83 97 33 15 13 53 DD 13 FA 3C FF 54
 32 B6 14 52 D8 CA 9A 01 F9 E1 5F E7 65 C5 70 83
 1A 9A 53 B5 BF D6 6B 1E C8 F6 5F FE D7 02 54 F3
 1B ED A5 32 88 47 3D 93 A0 07 B5 47 D4 02 48 71
 42 FA 91 5C 09 76 8B 49 1B 69 09 F5 24 12 10 53
 62 AE 0C 8A 4B 06 20 B8 F0 3F 74 A8 85 E9 46 2E
 21 5A C1 8F 9A B9 49 5C 07 39 89 A9 59 7F 07 6D
 A9 B3 CA F2 99 B6 C8 CD 49 45 58 11 6E AB 5A 74
 E6 3C 77 8C 76 34 E7 63 BF 14 7F 84 F3 C8 D2 6F
 64 BD 20 08 EF 6A 36 43 56 0A 57 69 68 CB 09 58
 08 2E 16 DA FC 71 28 9C 9D 54 1F 14 F0 56 DB 3E
 E9 B8 E9 7F 95 BE 96 81 B7 7A F8 8F E1 2E EE F4
 0C 11 B8 1B E2 5C B9 D3 B4 4D 40 70 B3 1A 95 C9
 92 7B 5B 02 61 1F F6 90 F6 B2 A9 8E F7 61 9C DE
 BF 0B 63 07 AD C0 D3 C6 17 78 FD FB 02 6F 8C 4C
 F3 CF 53 F6 5A 9D 3E 8D 26 77 00 5C 8A D2 0E 2B
 E0 27 83 4B 96 03 C6 3B 1C 43 D5 3E DC 48 16 25
 6B 9F 66 DC 64 C7 E9 6C 28 76 DB 99 04 C2 A2 0A
 39 F4 AE 99 04 BA 50 DE D0 61 01 81 17 00 84 B7
 CB 60 E9 DD 54 8E 82 4A 25 A4 3E F7 68 88 F0 E6
 A8 D2 3B 4D 55 77 09 17 2D 2A 03 2B CD F7 6E 63
 3F 91 9A 03 6F 8B 21 85 4F 78 E1 21 0A 1C B0 8F
 68 CF 03 5C 08 E9 68 12 08 8F 7D 9D 4D 8D F0 A9
 43 75 06 D4 71 33 59 C7 62 37 CE 3F 93 05 E0 7A
 1E 28 89 45 F6 14 0C 77 99 07 D8 FE 21 F0 3A DE
 FB 61 3A 8D 1F C1 60 BC B5 66 FC 95 67 D3 0A 04
 B7 B3 99 B7 02 9A B7 8E E1 7F E7 81 6A BC 6D 3D
 9B B4 28 55 CE 10 56 FA D9 3A 0D 68 CD 8B 9F 5E
 FE 7B 7C 4E 94 30 7D 85 26 FF 01 AD 77 30 E4 2A
 45 1F 4F DC 74 96 BB 98 CE EB 43 CD 2D C6 DA D9
 B1 D3 06 4A 23 64 F6 52 94 DB BD 34 A0 DB AB E8
 EB F3 9D E7 46 B2 59 26 BC 96 B9 9A E3 71 6D 3C
 7A B4 C6 9C 4C 18 D8 65 DF CC E5 DF 3C D2 46 EA
 D1 06 1D B3 4D 87 2C F3 F1 50 49 CF DA 6C 59 94
 B9 8F F6 86 B3 42 F0 F4 05 FD 24 36 18 80 09 09
 43 1F F7 8F 37 28 B0 50 1B 7C 37 1B 60 12 0A CF
 7D 1E 91 56 D2 3B B1 A3 5F F3 0B ED 2B CB 4C 22
 DE 11 9B FA D6 D7 4F 7E E3 5B 13 2D C3 59 96 63
 4A DA B7 1F AA F0 38 F7 57 01 88 5D EE 66 33 3E
 84 3B 98 B3 4B D3 FA 05 AD 8C 55 77 4E 7A FC DC
 01 68 3D BA 9F 6E 84 E7 BC A6 84 5A 0F 8E 88 B7
 2A 69 EC F5 DA B0 3D 1D 48 4A FC FA 15 2D 75 7D
 68 DD 03 3D 00 10 29 34 A4 2E 41 AF 94 87 0D A1
 E3 6C 5E 97 EF 1A 7A B9 4D 52 38 EE BA 3E 0B 29
 E1 F1 DB 64 9D 87 6C 6D DF 49 A9 20 DE 87 7B 29
 0F 19 05 A0 2E 86 4F 2D BD 82 EB A5 7A F6 60 F7
 0F 0D C9 BE A5 DF 35 FD 5C 1D 5B 69 74 4D 52 77
 37 44 9A 1E 6F B7 36 C8 44 33 42 52 F8 68 F9 8C
 2D 6A 29 FB 4D E7 35 10 58 E4 E4 E5 2B FC B2 0F
 A0 49 E1 E6 D4 66 1A C4 55 70 08 87 E5 16 E6 9E
 7D 6E A4 BA 7A 76 57 FE F5 0A 85 14 CE 64 17 98
 E5 37 0A 63 36 9A EB 1E 60 67 EF AE D6 89 82 08
 C6 2B 89 A6 FE 93 50 1F 64 BE A2 71 A2 62 10 05
 20 B7 56 75 44 1B EA 60 A6 52 00 C3 C0 93 E0 6C
 CB 00 AE 31 59 F7 37 81 A9 0B 15 A0 82 24 E9 9C
 AB 15 EC BE A6 B4 27 9A CF 30 5E 98 0E 99 A6 2D
 7D 64 EF 7A 1F CC 2E 2E 31 31 03 C4 87 AC 8C 83
 2D 46 D5 39 78 FD 5D 58 EE FE EF D1 80 A4 A1 88
 16 D2 10 F2 38 11 35 BD 2B F4 1E 54 17 07 71 32
 21 6F 8C E0 9F 39 8D 1C 07 2C 2C FE 43 19 05 D5
 78 A2 3D F6 77 6C 24 13 8D 13 61 6E B4 FE CA 16
 2B F7 20 19 11 E4 4A DE B0 27 1D F1 65 ED EC B9
 55 DB 56 3C B4 01 51 36 E7 31 E9 BA FE 0A E0 65
 56 36 7E 8F D5 E7 AD EE DE 84 C9 4E B4 B3 95 FB
 20 C3 D5 A3 4E 53 98 AE 47 7A 2E AD 6E 00 52 D3
 6B 5A 71 F7 B8 E5 A1 BE C6 AD 12 07 0E 7A 68 C7
 B8 62 86 D1 43 68 8E 87 D7 1A AB 0B 4B 4A 8D 5D
 50 CD 60 D8 9F EB 82 D4 C8 55 0F F2 FD 0D 99 08
 25 D6 95 61 F7 16 C4 19 21 B7 F6 CD 8E C2 4D 9C
 9E 13 D4 7A FD 41 1C 0E 1E 72 6A 0E 95 1F 2B B8
 F6 33 1C 59 DF D8 C9 06 6A 3D BC 5E A8 67 61 50
 79 6F D0 4C 2E D2 83 F0 46 5C BF 3A A2 D6 38 65
 12 0A 30 F3 91 A8 6D 67 7E 68 72 89 4C 64 F6 81
 F8 88 CB 86 16 72 BD 1E 50 85 88 C6 D4 A6 EA BA
 2B 05 7C 5F C5 49 39 CB 4C 9D F4 49 36 78 6E C8
 47 5B 13 65 86 41 87 F8 4D C9 89 EC 83 F8 16 B0
 FB 20 02 86 2C 42 50 74 9E 4B 53 3C 8C B9 A6 DF
 39 61 AD 1B FF ED 68 7D 35 ED C4 F8 81 72 8A D0
 6F A1 7F F5 C7 BD FF E6 8F 20 18 73 45 69 12 83
 63 28 15 80 31 EC E6 82 67 62 AA 53 63 32 6C 9A
 A1 03 A5 85 6E 13 A1 02 D3 C1 B1 24 F5 40 C7 6D
 A8 E5 03 15 66 68 15 A3 A7 01 6E 57 7F CE 70 92
 41 4F 9D 71 54 8C D5 35 C2 CB 5F D6 4F 37 67 9E
 65 0A 1A 76 7E 13 4A E5 96 E4 E1 A3 6E 87 A6 B5
 10 12 AC B5 15 BF 2B B3 23 48 17 42 52 37 57 B1
 9E B2 6A 44 10 DC 10 81 95 C5 B9 A4 B5 CC 4C B5
 BB B6 79 C0 E9 26 32 F8 61 E6 23 E2 25 FA A5 8F
 65 1B 83 55 04 A8 03 DD C1 25 6B 87 3E 51 79 4D
 EB 8E A2 28 78 C0 D6 07 B8 39 F9 16 49 9F 3C 2F
 4E 0B 64 C8 92 13 65 FC 3B 2C 7F F4 4C 80 44 0F
 06 7B D7 84 B6 6D D4 AB D3 61 C6 5B 02 92 9D 3A
 68 EA AA 3B 92 B6 30 01 37 C0 27 4A 5E 18 E2 13
 01 F4 CD FF 94 19 24 58 77 D0 28 5F DA F2 EA 2A
 A0 7C 50 5D AE 8D FC 26 17 96 C0 E8 62 A9 CD 3B
 4A 6B 3A 7A 21 F1 D5 36 12 02 80 5A 24 AB 08 96
 BF A5 E7 FC 5E 45 12 A4 26 2D 94 92 8A 82 DD 68
 F2 56 4C 3A 5E B6 F4 B2 1C D7 04 8A 66 28 37 CA
 6C 3E C2 4A 93 38 61 F1 31 8B 86 46 DC 78 DD 04
 AD 46 35 BD 6B 12 87 7C 01 00 91 60 A3 3E 94 14
 63 5B A2 AD 99 DB CE 9B 71 C1 F5 40 5F 47 9E 46
 A2 FA E6 EE 02 60 9F 6A 34 0B AE 06 20 8D 47 8F
 33 78 92 F4 96 E7 05 1C E7 39 85 44 DC F5 DD B7
 79 AA C8 0A D7 E5 91 37 6E EE E5 26 79 E1 97 F8
 9E DD 5F 3E 30 75 A8 5D 0D 79 19 33 0D 93 F8 A5
 84 8D 7E B8 D8 87 C0 37 0A 15 45 F5 13 32 8E 17
 F2 2E 40 9D 50 F9 D7 B1 D7 39 96 CE 83 B5 4E 82
 58 6F 5F C9 FD 98 96 3C 06 6A 6E C8 9E EE 81 EA
 DD F8 60 06 4C E6 2C 48 68 8E B8 CC 7D BB CE 77
 33 8E 1E A0 4C 32 24 49 6E D4 68 15 08 83 3E 2C
 01 CD A8 50 42 6A 6A 35 92 ED C4 05 D9 CD FC 88
 5F C1 51 D5 39 08 E1 1B 92 7D 1A 84 60 95 F0 AB
 61 7D D3 6E 37 4A AB CB 2B A6 6D C8 4E 50 9E 06
 B2 30 92 41 62 76 6A 7E D9 42 C3 7A D0 C7 82 CD
 13 80 31 0E 85 E1 71 69 A7 C6 AC FF 91 5F 4B 86
 5A F0 34 08 03 20 35 BB C0 14 84 29 02 5D 28 C0
 C9 46 A2 52 2F BD 8E D3 5F DF 53 A6 77 22 A7 65
 2F A1 2D 95 70 38 A7 37 A4 84 4F AC 04 BA 65 68
 21 21 B4 6B 77 B1 66 95 94 4C 96 AA 5C CA 0E 53
 2E D5 21 4F DD C6 95 92 D7 B9 84 1F D6 0E C4 F9
 56 57 2C 52 73 6C 88 0D 7A 8F DC F2 96 31 8C 8D
 FB 87 C7 C3 28 96 A2 C3 CE 8C 20 46 9D 7B 9B 05
 78 2C 87 09 23 05 95 89 99 7B 81 DE 07 15 34 FE
 23 3E E7 C4 15 68 3F 13 70 93 E5 FA 23 36 71 3A
 2A 2F E7 FA 7F E1 04 24 83 19 03 89 B1 34 BC 82
 72 A7 BF 3D B9 0C 21 77 54 BC 3B 57 E5 15 F5 3C
 45 2F 92 C9 7F BF 4E F3 2A 00 B4 C7 AC 1C B1 40
 DE 59 39 55 41 E6 3B BF 5B A2 F4 6D 85 35 14 82
 F0 EF 45 FF EE BD B9 A0 10 DE 11 9D 9E C9 7D 81
 D2 36 06 D2 A0 C0 41 E3 70 63 E9 39 D9 DB 00 83
 DB 7A 2B 0F 95 95 E8 2C 41 AE 7E 46 30 F7 60 73
 1B 2C A2 AD 17 CD 9A 38 50 EE F6 E0 7A BE BD F0
 D9 34 E2 59 C7 8E F7 AE 42 98 32 0C EE 48 78 DE
 25 8D 5E 94 ED BA BC 24 64 D0 4A 1D 55 97 DD A4
 79 A4 3C 5B DE C4 03 24 AB FB 2A 3B E3 71 74 B5
 F1 44 28 E5 06 C8 B5 18 96 DB 71 74 0A 9C 79 1A
 FC AD 91 F7 05 2E D5 C2 2E E0 75 EB 6A 26 FA 3F
 DD 34 C6 41 C8 BC 1B 35 80 0F 1A F3 38 68 39 0A
 DD F4 18 43 FC EA 6D 49 35 AC EC 5E EB FB CA 6D
 3C 71 59 74 8D 20 B9 BC FB 30 5E 99 2D CD 2F B3
 3A 4D 7D 8F A0 2D C5 FA 49 84 8B F7 1F 74 21 DF
 7F 89 6F FE E2 4F D6 3B ED 83 B8 76 40 5D 4A 15
 C8 C1 63 B3 AD 92 E3 35 0A 58 B9 47 B7 03 C2 63
 27 C6 A8 4C 41 DF 34 69 FF 6F 54 D2 34 EA F1 14
 E0 C4 70 8A 20 21 A6 4C 19 62 B6 04 A1 E5 59 78
 45 92 9E 3E E3 95 D7 D0 44 20 9D 92 5C 80 D0 6F
 85 D7 E4 C5 C3 50 53 E5 F6 DA 79 29 F3 22 1A 85
 3A B7 99 54 31 28 7B E1 64 DE D3 33 05 83 AC 2D
 13 39 3A 50 8A 05 15 A9 EB D2 44 2C 23 44 84 32
 31 F2 9C B0 F2 92 C5 D3 A7 91 98 C3 3C 5E 7E 25
 ED EF 25 F1 6F 64 47 15 D8 71 C8 BF D4 1D 27 90
 AF 05 66 CC 8D A2 AA 02 EB BA 33 44 91 08 06 35
 8E 3B CB EC 57 6D 63 5E C3 7F D7 45 30 D6 D9 BA
 2D D0 ED 66 35 90 24 D4 FF B1 0C E4 2F F4 9C C3
 98 15 E5 55 ED AA AD EB D7 41 8D 07 A5 74 8A 8B
 88 7A 56 BA 60 55 54 5B 36 2D 8E 6F FF 92 3E A8
 66 3D 6F DF 85 9D 17 CD 11 1A F8 0E ED 05 A6 54
 CB 52 40 1F C5 B0 7D AE E9 3D 3C F7 F6 89 97 24
 C0 93 00 74 02 05 D3 0D 64 89 63 3D EE 08 25 D4
 32 53 A2 08 C7 56 35 97 29 90 22 1E 48 52 C4 CA
 78 91 66 14 88 89 02 7C 67 7D 9B AE B4 57 09 67
 10 77 F7 D3 14 05 3A 6A 90 62 1F 44 77 AA F3 2E
 AB C2 53 CD 1A C5 33 DB F6 16 5E F6 BF 5A F2 12
 48 EB 7F 74 9F 8F 32 15 4D A0 43 93 8B A9 F0 62
 CE 1A 65 E6 E2 B6 49 D3 44 4A 18 F7 8A E7 17 EC
 EB 4C 88 A0 28 99 A2 27 7E 11 30 41 4D 35 54 D7
 EC 8A E4 86 BF 79 CC 5E 07 CC E3 D8 BA 30 7A 9D
 44 D4 13 FA EF 99 C7 29 66 23 64 B7 42 0C 7B 46
 B7 98 88 9E 8E EC 3F E7 C6 86 90 00 65 F9 5A 1E
 EC BF 2B 10 00 0D 0A B2 88 07 54 26 28 52 3E 6E
 CF 3B BF 96 CF AD E5 6D 26 1F E1 73 08 44 80 FF
 03 B2 DF 01 59 A2 76 6C 44 17 1A 54 91 4A CD 72
 38 A8 C8 F5 56 C2 D9 15 58 C0 EB 12 38 1F 8B 79
 5F F2 C6 77 B5 20 30 41 BD 0B 13 6A 71 56 22 95
 F9 CB 51 AC E3 D3 E5 61 68 56 6A C5 43 58 C3 66
 9A 5E 53 62 F3 0E E1 46 44 AF 11 9B 05 50 16 B7
 23 39 8E 46 1E 5E D4 FD 69 72 26 2B BD C2 C1 E8
 29 C5 87 98 01 4F E8 79 BB 51 6C 3D 2E 05 C3 9E
 EF CE C2 F3 F8 28 B5 DA 90 71 56 7E B9 D0 A5 B6
 6B 5C BC 77 B1 15 17 02 9B 9B BD 19 A0 AB F3 25
 CB DB C5 FB 57 A3 93 27 03 7D 95 02 DD B0 EF C2
 D2 0E 3D B2 26 E2 51 CD 8D BE 14 51 3D 22 EE F1
 39 8A 63 37 5C 23 6B D3 5E 53 77 21 4D 44 B3 33
 A4 6B 51 14 1F 1F 92 47 F2 F3 02 E0 1D C5 AA 37
 DD 4E 61 ED 1B AC 21 0F 85 A2 26 2F 69 34 6E 2F
 71 60 5D 5D 8A D3 FD 79 AB D0 3C 92 2C 0C 74 D6
 F5 7E 8A 6B 23 E9 87 5D B6 8D 01 5B 66 F6 6E 78
 C3 FD 31 C4 42 13 3E 38 62 8C 78 97 A9 5B CA 52
 8A 50 78 AB E3 0F 86 B5 74 01 87 E5 E5 4E 30 AB
 15 07 22 3D 26 BA 0E C1 95 81 76 F5 F2 58 7D 8B
 8A 72 02 F7 FE EF D4 A7 78 A3 8C C9 FF 11 D0 15
 CC 64 48 AB 4C 22 C3 8B F2 9B DE FB A8 BB 1D 00
 FE A9 CA C4 2C 57 6C 60 75 AB 5F FE 9D 79 8E D8
 A8 36 B6 C6 47 43 22 D4 51 E5 82 28 8F 1B 9F 18
 20 D9 C6 4B 28 B8 4F 9C 95 89 D3 2A BB 35 0B 41
 0B 8C 4D 18 7E 64 11 16 9E 51 83 A8 34 CD 1F CA
 A2 DB ED 51 CA 16 73 E8 1C 85 82 D6 47 37 6C AB
 D4 84 89 B8 47 89 D9 ED D5 F8 2C F1 E7 73 B5 F1
 68 87 43 EA BF 91 FB 8C 2F C4 EF A2 E2 F7 62 F1
 F4 BB CE 79 5E 0F 68 3D E0 ED 76 AB 2C 3F 2C 7A
 47 E4 B3 1E 3F 82 50 4F FA BB DB 3F 19 BF 15 95
 AD FF 4F F8 25 5E B1 60 7C 40 7F D8 77 54 D4 3A
 59 FF 50 91 74 52 AF 81 C2 F6 63 43 EA C4 65 B2
 04 CF 47 8D B0 79 6A 98 F0 A9 34 EC D1 0E E4 B4
 EF 52 B1 D0 54 52 55 B4 00 92 25 E3 1F 40 8B 8E
 4E 0F F7 50 B2 E1 80 B4 6E 48 15 50 B5 93 DC FC
 84 35 AD CE 8E FE AC 1D 44 B8 E1 9E 06 85 9B D0
 1C 5D F0 8C 64 F6 B5 92 23 AB 87 7E B0 A9 16 0D
 FA 84 A2 94 0A 48 CA 71 2B 22 E2 63 D1 B5 29 49
 A1 D8 63 88 CD 2E 3A 53 DC DC D7 92 65 3D 67 42
 AC B1 4A F1 18 A8 42 69 C1 C2 CE E8 09 63 A6 0B
 63 29 41 36 DE 81 DE CC 22 7A 24 36 F0 A6 96 89
 17 FF A2 59 AB 50 CF C9 34 20 57 4E 18 5E 3B E9
 A4 63 C4 5C F7 6B 3A FA 4E 94 56 D0 1C 14 08 DB
 53 E0 19 BF EF A4 C0 1A 14 70 1C 70 4A 5A CE D5
 24 04 79 51 C5 0E D1 42 90 13 A7 11 BE 86 B0 01
 6E FB B2 B5 E6 B8 B2 12 1B 9A 6F 6B D1 37 42 3D
 53 39 4E 73 F8 A8 6E B9 0E 0E A9 5B 74 AE C2 22
 7E 3B 4A D9 91 FA 2E 77 8A A0 B0 21 E4 49 18 C6
 67 54 48 7E F6 E3 84 F2 CE CD 01 BA D8 58 C7 40
 14 61 6F 8A 7E DE 4C C6 96 7C 5F 3E F9 3F AC 48
 F0 CF D7 42 EF 17 55 DB 2F 90 CE 6A 08 58 BF 57
 5E 88 13 B6 5D AD 9A A5 63 DC FE BB 55 A7 1B FC
 39 2C 99 D6 F8 6D 2B 91 8A B4 3F 94 6A 52 91 28
 F0 14 E7 28 EB D9 78 00 53 3F 49 11 5A 5D 18 B4
 1C 43 60 E0 03 66 18 12 6F 93 3E 7D C7 0D F0 F3
 75 85 A9 AA FD 34 D5 3D 71 4D 1E 0D AC 4E 25 19
 A7 BA 25 FF A6 9B 7E C0 0B 38 16 66 E1 28 34 C1
 9B 28 17 37 E3 94 32 3D BD 0A 1D 68 8F 0A 83 A7
 D7 14 82 0B F1 8A 32 A9 0E DE 16 12 D7 6A 9D B2
 C3 48 DA 50 76 49 F4 D2 74 65 6D 7F 0F 65 DE AA
 77 2D 98 5F 33 B4 E8 64 5F 69 EE 1E 04 52 25 07
 5E 0C 61 BE 07 40 BC 03 F1 6E 2D 54 58 5F A1 53
 52 B0 DC 19 C0 D9 12 68 91 BB 65 2F E2 20 9C BF
 FC BA 70 9E 88 F0 F1 46 83 87 78 5E 2A 33 78 8D
 18 2F 54 0F D7 D0 27 9C 46 8D 68 58 70 54 7F 90
 DE BD 21 EE 3B 67 01 F1 10 29 0F 02 C4 08 C5 A4
 88 F6 44 44 C8 C6 81 20 D4 D4 58 C0 C1 2E 1C 62
 C5 89 CA 50 6A 26 5F AA CC 55 DD 43 2E 38 49 63
 C6 3B A7 ED 21 4B EB 5F 84 A3 BE 59 F4 DE 69 AE
 EB D7 FA 79 CC 54 B2 84 9D 04 D2 31 0B 9B CE C0
 47 BF 63 C2 2D A1 9D D0 F2 7A 51 35 37 52 B2 4A
 DD 0A 5B 1E AA 37 A5 E9 D6 0D 47 94 E9 28 2D CB
 75 C9 70 0E 26 81 6A E4 49 25 87 02 F9 E3 67 43
 BC 34 47 29 B5 11 6F 20 E3 DC 28 38 EC 81 FE 96
 DF 8C B8 5A 79 31 8F F3 A1 0B B6 72 E1 8B 8E 9B
 42 07 57 8D B4 78 3C 70 42 41 9D EE 30 94 DC 96
 F9 5E FB AC BB 4E 4B B5 75 6E AB 40 A0 0D 23 19
 C4 A1 37 17 D6 EB 44 78 49 D7 98 61 7C 17 02 C6
 D7 20 37 8A 6D 40 0D 92 51 7C 8B 3B 10 A1 00 CB
 61 A8 3C BD 13 D9 BE 27 5A DE D4 C3 01 A1 42 50
 F8 07 15 97 F7 C5 59 13 11 AB EA 13 C2 1A AE CA
 44 DE 95 3E DD DE E3 FA 66 51 DF 86 E9 89 59 87
 77 C5 78 09 CA BC 53 F2 0D 7B 78 1E 29 AD AD C1
 F9 22 9A E3 5B 25 AE B9 A2 CE 9F B3 64 6D 0A C1
 D2 FB 05 F9 BF EF 9C 6C 1E C6 80 0F 62 A8 B4 E7
 79 28 2B 96 4D 14 AB F9 AC 36 0E 0C 5B 53 DB 8F
 D6 70 56 1D DC 6A 2E FC FA 2C AD 78 8D A4 26 90
 14 64 0F AA 24 10 7F C8 14 96 9F 2A EE AD C2 23
 63 28 2C C1 37 8E C9 B5 8A 56 DB 36 18 F1 E5 F8
 BB 84 6B 7D 13 F2 95 27 23 EC CB C5 17 B9 D1 E4
 E6 0E 33 DD 78 F1 33 24 C0 3E D1 14 A4 AA 1C 5B
 1A FF 06 BF 9B 6F 36 40 E3 01 7E CD 24 12 71 24
 EA 06 45 EB 85 42 54 E8 96 0D 68 44 B8 70 12 42
 56 D7 06 39 04 7E 97 33 D3 7B F4 3A 74 71 08 18
 05 2B 17 A0 C8 46 45 CC 9E 78 3A BF EB 35 96 E5
 FF 71 87 F5 DF D9 D0 18 1F F7 DD 17 DB 28 32 98
 37 2B E8 4B 09 70 0E AB 6C 82 1F 57 25 B0 13 74
 ED 0B BF 92 BA AB 7B DF 53 55 3B BF F3 EA 3D DC
 4C C8 23 58 3E E6 6C 45 5E 12 4E 37 D8 8E A6 1C
 9A B1 79 A1 BF 59 F4 4F F7 EE 1E 46 44 25 9B 08
 64 49 C7 35 CB A9 CC 32 67 3A 12 9D 81 5A 0A C0
 FD 60 19 A8 18 AF 84 00 C0 4D 3B E1 95 A9 D8 A5
 B7 1E 9F 11 CF 5F 50 C4 C1 54 3F C1 14 9D 4A 69
 3A CB 74 23 AB 78 29 8B 67 25 15 1D 0C 17 AD 81
 45 E1 23 C8 98 E2 4F AD F3 AE 0F 42 CB F9 24 B6
 EB ED 2F 45 D4 05 63 3A FC D5 71 57 00 AA DB BE
 0C EE E1 30 14 67 1C 12 7A 7B E2 6F 84 2F C9 41
 4F 1F CB 20 F3 42 B5 A3 0D CA 43 D1 20 6A 13 A7
 8B 59 45 3D 19 7D FD D4 6F F1 B8 DC BA 89 37 64
 41 AB 84 98 32 51 EF 20 D4 BB 30 08 91 D6 E9 62
 30 1D 3A D7 12 CC 5F 67 CE 39 0D 92 C9 DE 19 67
 B9 20 55 EE 4F C1 34 D8 CB FA 22 C3 19 28 C8 8E
 A0 2A D6 4E 0F FF EF 77 3E CD 79 12 00 C1 3C 75
 4D 97 27 9E FF 10 C3 BB A1 2F 12 C4 CC F4 FE 44
 E9 A1 9C 29 3A 96 B9 C6 60 78 DF 07 28 52 FB 43
 10 8B 99 9E CF 9A EB A2 47 D2 E2 B6 6F 78 1B 97
 C9 1A E4 11 5C 11 86 FC 0B 40 8C 78 DA 43 42 D8
 1D 12 0E BE C7 B3 0E A9 AB C4 00 5F 12 07 52 CD
 B3 43 D9 EB 66 FB AB 94 B8 34 69 65 43 5E 82 DE
 9A 4F 74 89 2D 61 DD FF 7D C5 57 1F 2C E6 92 6D
 DE 09 C5 A4 6D C0 8B 0D C0 14 1E 8A BB 91 83 1B
 41 A9 DE 3D 87 61 FB 51 0B 31 FE 13 E4 67 CB 73
 15 65 69 84 76 B5 3D 5C 71 06 74 A6 26 D0 25 5B
 89 F5 44 6E F3 6F CD 27 EE 3E 82 06 5D 53 74 80
 6B 8F 94 2B DD CD B4 57 E0 9C 94 9C 67 F8 58 2D
 8A 29 BE E4 A2 96 07 04 6E 7B 5F D2 1B 31 8B 1A
 93 52 58 0A 97 91 D2 99 06 F1 33 FB D8 AB A1 43
 8C 3A 9A 0F 70 76 B2 DA 69 D8 B6 11 06 19 04 18
 E1 37 BB 45 80 C9 B2 9C 57 6C AF 15 E8 08 0D B5
 37 0E EB D2 80 F4 7F B0 B8 23 C1 5B 92 F5 98 51
 51 37 60 76 AE 7D 5C 9D E9 DF D2 99 92 70 9D 83
 B5 A9 76 5A 65 FD A8 8C D5 2A 9E 64 53 E9 C5 CB
 DD 54 4E 7D 23 FA FC 04 87 A3 BC 0A 89 B2 87 76
 05 61 95 A1 C9 38 08 3D 1B 19 71 BB C2 4F A6 CB
 E1 AB FC FD D3 E7 E5 3B 11 A7 5F 38 FD B1 29 12
 DB 38 CD 9A 12 1F 12 C0 EF E2 8C FC 25 D6 30 23
 BC 71 A0 B2 72 B6 77 36 94 38 4A 15 06 49 B4 35
 69 B6 2A 61 91 AF 73 E7 BB 7E 34 05 01 19 A8 EF
 63 81 2A 98 3D A6 BB A4 88 E1 5A 9C AE AC 0C CB
 9B 1C FC 8A BC FB 58 B6 FC D6 E5 BC 01 40 C6 5A
 60 81 EE 95 54 32 DD 73 0D F5 84 4D 3B C0 64 1F
 76 CE D6 18 2A 24 DE 6E 4E 2B 5B 46 7C 3C 72 AD
 27 89 88 06 95 3E 51 8A 1E B5 90 77 BD B6 11 8C
 AA 3F 34 C4 D7 0A AF B5 17 56 49 4B 00 F4 9A 9C
 BF 3B E1 37 20 B2 08 4D CE B0 29 BD A8 FC 38 4A
 57 7B 28 C7 C4 D0 E6 FF E6 81 1A F9 85 C5 4D AA
 88 40 7A B4 F1 11 0B 49 A8 A8 00 05 6F 2C 40 8D
 90 D1 5E 30 8E FC 6F 06 E8 03 6F 3C 37 DB E7 ED
 31 95 D9 12 8D 31 51 88 85 73 55 70 41 AD B1 D1
 2D 72 84 16 9D CF 96 EB 17 AC 9C 92 85 D5 F0 B2
 77 A8 E4 C7 53 4D A4 66 45 9D EF C1 1B 00 13 42
 EA CC 18 FB E9 D4 0D 84 C6 4D 6B 9D 32 01 3F CD
 FF 38 E8 26 F1 FC C0 6C 46 72 30 54 29 AD 2F E3
 CD D6 E0 27 A4 EE F3 86 AD 6A 40 98 54 AE FA 7A
 DB FB 0C BB 04 78 24 45 B0 DC BA 2F 80 B2 0D 5E
 36 11 43 A3 A5 64 D4 3C C8 0C 13 B2 4A 2A 00 A5
 0E F0 60 B6 95 89 3C 70 B8 16 09 B4 7B 6E 0F E9
 48 6A 7E 21 F3 50 C9 6A 63 10 8C 24 89 26 82 B5
 8D C7 30 A5 35 DD 01 27 F2 45 F0 92 FA 2A AA B7
 2A 49 0F 4A 4F 5A 14 DF 52 CD 08 27 7F 9A 3C 72
 76 9B EA 51 53 DD A7 2E 0A 19 BE D7 4E ED 75 87
 9E BA 3E 78 C4 66 9F 5B 25 8E 7C 2C 0F EE 3E CB
 76 54 C4 F4 85 92 E6 55 61 E4 54 1D F1 89 49 99
 92 10 D0 A0 90 E5 F1 42 A2 BC AB 16 ED A5 85 6A
 3E 3E D0 84 69 F4 05 6B 36 13 12 DF D6 B4 6F 0D
 8E AB E3 F8 79 B5 FD FA 01 DC D3 E9 2C 86 07 92
 FD 7B AA 5A 5A 23 46 8F AD 2E FE 78 76 49 FF 11
 04 A5 55 38 A7 2E F3 DC 23 44 B9 98 30 F5 A3 47
 62 87 2A 0F B3 4C 75 32 9D CB 4A 68 15 A5 66 11
 63 70 E2 19 79 78 B0 8C 8C 55 58 5A 31 72 03 00
 3D 79 55 19 E5 B3 6D 93 4C F9 8C 6F A4 3B 78 37
 31 0E 56 65 36 28 C8 83 94 8B 23 AF 19 E3 4A D9
 12 97 4F 99 CF 3E 09 67 3E 3D C6 10 F9 C3 A1 5F
 83 DE C0 EA 0B 7C 71 EE 36 BA 74 E5 D8 A5 C0 04
 BB F0 46 E9 30 23 C0 D6 C0 DF 4D A3 11 89 C9 E8
 24 B2 B0 55 D8 2C E7 3B 8C 40 D9 2F 6B ED 97 78
 88 E8 F6 78 18 5A 81 49 C7 84 9E 6B D1 20 80 3E
 87 0C 5F 67 90 62 74 01 8A C3 E0 61 D9 DD 35 73
 B1 F3 84 31 24 42 93 44 14 2A A5 C5 7A 59 B5 9B
 92 38 8C 4A D9 D4 56 8C E6 42 07 A7 D9 82 D7 69
 8B 85 89 05 7B 3E F1 B0 64 DF EE 11 F1 2D 3D BD
 C8 B4 8E 31 9A 59 34 36 10 B7 B0 9C 50 F3 D7 D0
 B7 85 DA 4D C5 74 ED FF 8F A5 24 BA 5D B5 28 F7
 11 62 CB 91 20 E9 D5 EC 5A 78 1F 45 B8 D0 CF 55
 90 60 E0 D2 90 40 91 3D B4 74 03 4C C7 5E 58 5A
 3C 4D C7 8A F7 27 7B 89 13 2E 31 1B 82 C6 DF AC
 2A 8E 88 74 B6 3A 09 D8 82 F2 1A CF D6 A3 88 86
 43 ED 00 77 9D 0A 98 EF B0 FD E0 78 B3 F1 C3 4F
 39 FE E1 05 BA DE BF 6D 27 3B B2 B2 A4 B6 EB 91
 BF B8 7D 0F 59 7B 85 39 8B 77 CD 97 16 D1 9D F3
 2E 48 C3 A9 2C 0D CB C5 D0 6A 35 7A 9C 8F 6F 73
 59 90 5D 71 40 9C 08 B3 80 D6 F3 93 C9 2D CA F7
 31 37 9C 96 3D 82 10 95 D6 EC 53 8F 21 22 1D 90
 0B 84 37 5A 3E D0 33 33 32 05 F5 BD A2 D7 31 20
 4D ED DF 5D 64 00 B4 7D 3D FF E1 28 6E 17 32 B9
 67 EE B3 A8 78 EB 42 F6 11 49 89 BC F6 50 D4 88
 C4 9B 58 4C E2 D7 B9 E3 99 89 C5 31 5D F0 4D D4
 75 21 D5 2A 74 E0 44 B3 E3 14 6A E1 0A 70 A6 BC
 9D 2B 7A AF 7B D8 34 32 E2 4F 4B B2 9C 60 69 2B
 38 9E AE 16 5D 76 64 0F 9A FB F2 23 93 07 FF AD
 82 9A F0 7A 5A 49 C0 8D 35 A3 90 75 FC AF 38 B8
 27 6D 57 B8 55 E0 13 0E 6D 8D 85 F8 F8 27 41 6D
 26 AB 1B DF 1D FF 4D D8 C8 7D 47 A1 ED 82 B9 BD
 09 3C F0 5D F5 DB D1 9A 54 BF 99 3F B6 EB D9 59
 08 8A 82 3A A1 2E 48 9E EA F8 18 30 F6 9B 7F DF
 60 39 EC DF CF B1 68 C0 D6 1F 56 8E AD FC C7 DA
 A2 2E 89 5D 6E 9C 07 23 6A 45 B4 D5 88 D8 19 DE
 2E 34 7C 60 0F F4 DD D5 F4 1A F3 EA AB BA A9 43
 A0 C5 E4 51 BF E8 65 65 41 48 FD 17 CD E0 C6 0D
 AD 17 FA 20 A8 C8 48 D5 C8 26 EB 16 46 DB CF BF
 04 EC 37 38 F6 E9 D3 E8 BE 73 59 9A 41 6C 2C 54
 67 BF 4D DB E3 A7 CB AF A7 0D 6A 4B 23 83 C6 8A
 8A BB D1 91 0C 44 A2 72 B3 D5 F9 2C C0 75 38 D9
 5A 4E 44 F1 BE D8 2F 6F 82 2C 60 70 54 32 76 16
 75 06 D2 76 FD 92 4F EF AE 23 05 60 C3 83 E5 AA
 34 D5 7D 0F 54 BF 09 79 5B 3F 41 9F 1B 43 4E A6
 CA 14 D0 B8 E8 D3 C8 BA 6E EC 10 B9 F4 70 6A A3
 2E 72 7D 51 4E B1 4C 04 7A E3 88 6F 69 8F B1 D7
 9D 84 E2 91 69 09 5B D8 A9 32 90 30 4C F1 23 FD
 F6 F1 A8 58 1E 67 C7 6B C1 6A AA 84 EE 82 FB 6E
 70 AD CA 1E B0 45 AA 8E 48 53 33 67 CB 07 7A 8F
 87 AC 07 C0 CD 39 B9 A4 FE FF C5 AD C4 8B 9F C4
 A3 BE A4 40 C4 DD 97 06 FF BC B8 16 A2 6C E0 49
 1E A2 AD FC B3 0F 76 00 B1 2D C7 64 F7 B4 E5 81
 6D F0 2E 76 1E 46 17 1F F0 3E C3 74 79 AC 40 B2
 91 C1 8D 15 5B B4 F8 BC 3E 43 1B 2C 72 B9 53 85
 72 EF AC F7 D3 A8 34 9C DE B8 0F EC 3C F5 28 FE
 C9 2D 6A 24 46 88 F2 BB 41 2D 7C C3 EE 16 D1 74
 E9 8C 59 D6 CD 0E 39 95 D3 37 40 75 84 75 F3 D4
 9F 0D 33 58 69 32 F2 84 64 3D B6 B0 E6 8E CC 45
 BC F1 95 3F BA AC CD 5C DB 66 98 0E 93 CC 4C 4C
 33 E6 8D 01 FB 4F B8 7E 52 91 C3 57 19 A3 93 B3
 BC 92 3B 50 25 88 F9 63 A6 96 BE E8 9C 1A B9 3A
 45 C3 1E 8D 9E CC 60 6C 2F 3A C6 44 46 53 FB CC
 46 C0 F8 B2 B5 7F 25 DD 19 8D 3E 1E 4F 49 CF FE
 AB 8B 00 ED AD 78 D6 74 E5 E7 19 1B EE C0 B7 8D
 13 38 48 7D 4A 9D B1 6D 04 1B F0 42 9E 99 EF 4B
 15 D9 4F 56 2C 58 7E CF E4 74 E2 60 90 6A 57 32
 73 FC 03 2E 5E B8 F1 88 F6 3D CA 92 6A 17 BF C2
 EA 78 D1 FD BE 0A 33 5A 60 E1 CF F0 94 21 34 AB
 29 55 39 13 71 B6 23 45 74 8D 6C D9 B1 7B 74 77
 BB B5 68 AF A8 53 0C 1F B7 3B FA FB DA AC 18 AD
 3D 02 95 8D 8E AB 32 E3 44 14 98 AD 07 D4 4F 7F
 50 C3 96 AB A7 B6 53 F3 BF C3 85 E5 55 B4 E6 B5
 55 B2 08 40 77 01 7B 5E F3 9E 38 DC 2B 40 CA E3
 52 85 5F 78 20 5B E2 B7 63 98 68 F0 B0 FC BA 1E
 E2 3E 38 B6 BC D6 92 B7 10 51 36 D9 00 C8 E5 27
 5F 53 02 CC CD E4 07 40 25 87 AC 26 F8 E2 C1 75
 C5 1E 3E 3D 3C 4B 00 99 AB 3B EB 7B F1 53 83 CA
 80 1E 19 0E FD 2B 0E 81 C9 DF 73 DD FA F1 3D 05
 89 AC 4A CC 96 4E 5C 18 FE A0 24 B9 2E FB A2 AA
 8B 65 DE 4D 0A B4 6D 0F 9B 26 69 66 1E 27 7C 43
 1C E5 69 ED A4 DF 92 B1 B2 15 64 1A 2F 5B C0 EF
 3B 08 97 9B DC 47 59 37 45 55 31 C8 A1 DA 87 8A
 1D B3 8A 4B E1 B5 C7 06 A3 54 E2 07 E5 C9 76 74
 CE 8F AF DC F5 CE 02 B9 64 99 C6 95 4C C0 59 7D
 58 26 35 BA 06 98 7F F5 2F 3A 0E D3 45 1A 8A 89
 8B 1E CD 02 AB 73 73 AF 81 58 5C FE F8 F8 07 7A
 C4 F8 86 7F 0D 9C CA DF C7 3C F7 11 B1 64 8D BB
 C6 FC 1B 9E 09 8A 96 EA F6 12 87 83 5B E5 05 07
 AA 72 5D B1 55 3A 61 53 2A B2 DA 81 D1 57 54 7E
 6C 4D 83 18 4E AE A5 67 7D 48 AF 8D 9A C1 D2 FC
 4F AB 42 DB E3 D0 F8 9C A7 63 21 B5 60 4C 33 8E
 7E 7B F2 6C E8 42 C6 B4 3C 78 3F 17 98 08 A6 22
 33 C2 69 6F C8 52 29 A4 9B C2 7C 36 6A 89 1E 55
 F5 8E C8 E0 E8 2B 68 2F CE 7A 82 E1 7A BD 5E B8
 43 AF 1F F2 85 61 0C 70 A2 84 6F 09 B8 F4 73 52
 D7 CD E8 04 58 B3 41 1A E5 DE 59 2D 38 3D 14 3B
 02 57 9F E7 1B 73 7E D9 30 26 25 98 AC A7 2D B6
 7F 03 D7 B4 6F 83 99 97 1C 00 4D 38 C1 E3 59 48
 49 F4 11 A5 19 23 EC 1D 9B 4A CC 1C 40 11 E9 DB
 01 77 51 A5 4C EB F2 63 28 2F 25 F7 22 3B D2 11
 3D 62 6D C7 72 D8 C8 6D C5 D3 2A 3B 6A 41 0B BA
 64 12 42 EF 90 E0 39 03 07 F2 32 E9 3B 4E 61 C7
 D7 FD 68 F3 59 E5 C0 A6 28 42 EA 63 36 E0 C4 DE
 03 44 21 19 6C A5 D1 52 DB D5 BA B4 62 7F FB 9E
 D9 A8 43 CD 32 8B AA ED 72 6A 37 C4 36 C8 FD 72
 64 68 09 99 B4 3E 93 94 88 4D 31 96 6E C8 BE B4
 7D F9 23 0F 75 AD 17 2E 42 21 47 61 BF A9 EF 66
 97 30 44 FF FF A0 54 EA BC DA 6E 5B CE 38 18 79
 30 24 FF 83 B2 5C 24 F3 54 18 39 FB 62 E9 B5 2E
 C3 29 5C BC F7 94 01 00 34 F1 DB 00 75 CF CB EF
 FA 26 1B 55 7E A5 D3 64 A9 FF E5 94 26 44 6E B6
 00 13 54 D5 93 43 67 C4 A5 BB A6 BE 6D 6D 7E 98
 FB 97 83 14 D3 85 04 F3 8F 02 10 F5 7D E7 CB 6F
 5E 59 D3 4E 5F 7E 6C 4D 1C B5 F4 B2 29 2C 75 43
 E8 F1 9C 0D 90 C2 62 7F A4 31 F3 B5 DA 6D 41 DA
 10 3D FB E2 99 B6 9B 1A 1E 9C AA 6F 5D FD 34 5E
 F9 D9 E5 66 E6 4C CC B9 DF 13 70 FF C8 46 0D 37
 A6 B9 57 ED 04 4C F9 DC D1 96 CB DF 26 BC E6 68
 B6 09 37 F2 A7 97 AB 67 09 32 CD 9C 83 A3 25 DE
 7F 8B 17 80 C9 62 2B 29 80 9A BB 37 23 EE 96 01
 1D E2 18 D8 32 28 F4 6D 79 98 1E 42 39 25 F8 36
 78 B9 7D 00 3E FD B8 72 10 3A D6 EA F7 7C A3 47
 BF D9 EE 09 4F D6 25 22 EF 54 37 39 90 A3 DB D6
 E9 D2 F9 EB 2E 2A 2D 30 B1 BF 46 4C 2F 34 27 E1
 70 8C 17 FF 7B 77 A2 45 8C 61 D2 E9 40 EB AD 2D
 D6 38 15 24 9A B9 A1 0A B7 EC 7D E9 3A D5 16 AE
 57 32 28 E2 CA 1C 72 62 30 D5 E0 75 9D 2E 49 40
 C6 27 41 55 C2 3A E3 6B 0C 49 D2 16 19 FD 47 43
 6D 52 A4 09 5C FB 1C 73 27 3E 2D 18 F1 B5 65 0A
 C1 98 91 4A 97 57 7D 3D 90 1F 65 A1 40 58 F8 F7
 60 00 77 C2 75 0A 32 B2 24 97 A4 0A 92 B4 CC FD
 99 EA D0 D2 95 30 76 3D 8A D1 1A EB 84 21 3E 87
 12 7C DC A4 E4 4A F2 9A D5 46 39 97 3E 04 CB 7D
 36 F1 B2 20 A3 54 0D F3 1B 44 99 01 23 B3 CA 8B
 3B F3 DB ED EA 8D 56 50 65 0B 68 67 3D B3 A6 C5
 2B 06 9F 93 59 F6 DF 16 4C A9 2B 05 98 83 2C 5B
 8B 5F 20 31 14 AD FB 3C B9 67 A7 32 C6 56 0E 4F
 34 66 0B 5D 6C 0F 39 61 BE 85 D3 78 37 BB 44 1C
 38 94 55 39 B9 DE 3C 87 7A CA 52 62 FB 96 52 CA
 E0 38 A2 77 1E DF 9A 99 1A 3D 64 A5 B9 45 2F 6F
 1A 83 CB 38 2B 48 DA B4 FA 07 A0 18 18 5D A1 20
 C9 85 46 7D BF 26 B9 4F 02 60 41 38 6D 57 FE 63
 58 15 CB E7 EF 59 6B 6D 91 03 1F F3 87 F7 16 96
 F3 0F 79 4D A7 B4 22 B0 91 22 79 41 DE 32 1D B2
 04 A3 6E 57 3A 52 FB 49 02 65 96 50 9C 1D 00 AB
 8C 05 B5 17 72 CF 2B 1F 0A 15 33 AB 5B 63 19 28
 6F FF 22 E3 C1 A5 D4 A4 1C 48 73 62 57 B9 20 A0
 10 EB 41 FD E4 CF 4F EC 00 B5 DE AB 35 DE 43 AF
 97 C2 69 10 27 79 48 AA 1F 0C 7C 66 BC CF 6E 34
 08 6D 45 6F FC F9 1A 62 2C 1D 83 E9 9B 70 46 15
 3E A6 E8 D2 F4 81 3F 61 12 47 6B 98 D2 9D 11 67
 B4 DD 22 7C 07 FC C5 72 BD 2C 6F 94 AD 3C 56 78
 7A DE D9 C5 C7 B5 45 66 D6 E8 78 CA 7E C9 8A 50
 04 9E A2 99 75 2A 32 18 60 30 BE 2D F9 E0 9D 51
 A8 C7 6F DC 78 9B 95 32 1E B8 66 11 FC E8 49 8D
 BB 2D CA 1A 53 AF FB C1 3C 0A A8 2F 02 BD 3F 33
 21 4A 3A C5 26 D5 6E A3 48 49 DB E3 9E 62 D6 F9
 0D 5D D0 0F 8B 68 F9 37 37 89 24 EA EA E1 13 9E
 79 4C BF A5 BE 4C B3 3C 83 46 08 AD 9D B2 B5 CA
 AD 78 D7 A6 0F 61 BA AA 17 D6 E1 4E 4C 3E 8D 35
 24 79 ED 01 79 32 05 2C BB A8 15 43 B9 21 22 6F
 13 18 64 11 FA 02 EA 34 9D 87 76 F1 2D 64 DB 76
 7E D0 AC 31 25 33 F1 A3 C0 6C 3F 81 3E 7A AA 70
 38 64 A7 DE A4 71 F9 56 55 BF 3F 5A 5A EE 66 43
 B6 BE 7F DC 44 93 6B D3 19 50 CF E0 9E 29 2E 94
 3C 37 77 93 36 AA 6E 4C 82 AE 87 22 8A 94 08 35
 FE 88 0E 1C D7 E9 70 CE 12 22 9A 8D 2A BE 89 36
 1A E0 D6 21 4E 14 BC 7C 9E 33 BE D0 1C AC 67 08
 45 D9 C8 5C E1 A2 0F 31 4F D1 1B 1E 60 50 CC F9
 B6 5C C9 D8 28 F9 8F B0 25 18 87 A4 7F A1 F4 64
 DB 89 62 D0 D3 CE 09 1F FF 24 C3 08 B8 EC DF 96
 C6 89 AB 61 1A AF A3 00 FF 3D 24 E3 16 61 58 C0
 3A 26 6E 73 A1 F0 1E 48 FA 43 21 41 64 97 74 80
 F7 AD AF 7C 37 3A EF 08 74 D2 04 E9 89 F0 C3 00
 01 1C F4 7C 3A C9 A5 38 60 81 46 B5 FC E9 CB D1
 C1 6B E8 41 14 D9 5B 49 1C 76 B6 D3 19 4F BA FF
 25 5A 3E 89 D2 5A 5A 7B 34 17 34 4A F1 03 2A 74
 8B 23 6C DC 0E FC 7C BD B9 86 C7 59 8C 26 A8 A1
 60 32 E9 C3 EA AF 69 00 84 C2 FD 63 F8 D9 1F 04
 F8 DC 1F 66 77 3C 66 78 63 F1 44 D2 C2 E5 E1 18
 60 67 1F AD FC 95 B4 B0 23 34 10 EC 13 C9 3B FB
 E5 B3 B5 B1 CC 83 71 3A 8B 74 3E BB FE C6 42 89
 89 F4 B6 04 9B 0E F3 F6 CB 1C 86 7E C8 82 26 27
 30 ED 64 35 CE 40 87 0D 24 FA 23 CB 00 51 EC CD
 D5 23 23 94 B7 50 55 A6 E8 68 D2 27 5B 4A FD 54
 93 32 F1 75 28 F8 44 2B 67 93 E4 22 11 41 B1 80
 D7 66 D3 EC 47 CA EA C3 9E E7 B2 73 94 49 E2 2C
 89 AA D5 8C 75 99 1D A2 CB 2A B1 4D 7F 7B DB CD
 47 E9 82 48 C5 3D 4B C7 8A B0 26 96 9F D4 B1 05
 0F 20 36 6C 52 65 90 50 92 BA 05 73 64 4D 3C E6
 B0 FC 10 DF 61 E3 D2 52 7F 17 4A 0B 7C FB 1D 4F
 66 10 0B B4 E1 4D E2 0E 4D 6A F3 5F DF FB 17 11
 8F 55 4D 9D 69 75 FF 16 5C A3 47 64 22 B4 52 B5
 A4 39 DC 02 EE 0F 7A 40 15 90 B4 EF 0A AE E4 B9
 5B BF DB BD A8 08 F4 80 7B 3F E0 80 41 64 49 4C
 92 80 FF 7B 3A B9 F2 24 28 5C 0A AF B3 3E 7C FB
 68 29 5E D4 5B DD 2E 31 DF 82 5B 07 31 65 F1 F7
 3F 64 5F 58 17 B0 01 3B EF 02 4C 00 78 0C AC 91
 36 98 FD 25 0D 63 5B 4F DE 39 D2 38 32 D5 FD 52
 68 B3 84 D0 72 A3 F5 70 D7 19 BF 2C 54 42 A2 1C
 63 D4 57 9B 76 0A DB 7C C6 0C C2 9E 5C 36 5C E0
 0A 69 1E 5E E6 2D 07 66 BD 27 9D 03 EF 23 A7 1F
 71 30 A6 69 6D 27 35 B2 EC DF 21 04 BE 15 8F 55
 1B D3 CD 2D 0E A6 7C A6 2F 4C 7F 4D F5 E8 76 17
 9F 87 BA A2 2D 60 30 93 A5 1A FC 72 25 E3 52 B6
 99 B1 74 75 98 41 11 53 21 38 A3 24 01 75 01 16
 3F 6C 42 7E DE 82 49 8D 9A 50 B9 4F BE 56 B0 72
 BD C4 05 0C B8 65 D5 D9 97 1C BE 68 BC 40 67 69
 81 E1 E0 5E EC 3B 27 F0 38 87 1F B2 86 7B 06 E1
 9E B5 FD 3E 10 B8 FC F5 B6 B5 1B BC 2F 67 5C B1
 77 5B 6C 95 20 D0 B6 9B 53 6E D5 CC 7E D8 9A 90
 EF 31 95 13 4F 10 76 2D 46 64 A2 75 96 91 5A 7B
 F7 15 CA 85 08 6A 8F 02 B7 D2 18 81 27 34 A2 2F
 35 B4 30 3E 15 2B 38 E5 B2 FD E8 F0 73 42 B9 07
 6A A0 A0 5F 51 E8 B1 B4 51 2B 01 81 66 34 BF 15
 E5 2B B2 C4 37 4E A8 D0 0E 6D 99 1A E4 89 F2 84
 AD C1 F5 73 7B 55 34 CE 8E AF C9 45 00 DE 15 91
 10 C5 3F 27 17 C4 5C BB 50 D1 8C 60 79 E9 01 6E
 37 28 0C 2A AE 8D 87 77 5E A7 4D 9C 4F D6 A3 75
 BF 97 1A 6B 99 52 12 4D 61 28 45 EB 88 08 66 F4
 50 12 87 37 82 A1 55 A0 FC BC 89 49 B2 E2 79 D3
 21 A5 61 94 66 6E 2C 7E 3C CB 6B 58 EB D1 2B D1
 EB 3C DE 03 F5 C6 92 D4 5B 3A E6 19 3F BD 43 89
 1C 5C A6 36 16 6C 02 87 5A 2F 71 FC 34 96 E1 2A
 92 6C 5A 26 DA 07 EC F6 D2 46 AD 7B 46 62 C9 07
 C8 17 35 B4 FF 8D 75 D6 A0 07 77 66 51 45 69 1B
 CA EF 48 7D DC 42 90 0A B3 97 84 F8 17 25 39 05
 74 B7 78 19 64 62 4E 13 E5 F5 D1 C5 5B A8 E6 0A
 2F 01 F8 48 D9 F3 8A 85 0E 66 88 AE 54 C4 ED 58
 2A 5C 16 A9 3D 4E 7F 93 99 6C 6B F1 AF 00 B3 9F
 19 87 E2 92 C1 F5 0A 31 70 55 48 49 FC 4B 6E 4D
 9C 4F CB BE 27 EE A8 7B E0 56 10 2E 8C 22 89 C2
 5B 8C AF E3 6C 4D 61 50 FD C2 B4 89 B1 F6 74 F0
 80 1B 92 F8 0B F3 12 E0 8A 0C CC 02 D9 EC E4 91
 2A 0F 6A 8B 2A 8A 6A 97 6B 3D BB 93 19 53 D4 8E
 79 0C E2 16 98 69 2B 4A 89 04 C9 58 18 BF 2C E7
 51 04 27 E2 72 50 E0 B7 B5 ED E1 48 67 2B 2C F4
 3C 61 4A 80 75 71 90 8B A0 2D F0 EF EB DC AE F7
 45 EE 24 05 F9 95 46 6A 70 A1 FF 7D 83 7D F0 6C
 66 7D CF 46 67 55 B7 27 94 13 4D 42 D6 BA 31 0E
 9C 68 CA D4 41 1E A7 E1 F4 30 1D FC 0D C9 EA 69
 6D DE DC 30 82 C2 B0 B3 EA 69 C6 4A 2A 90 19 9C
 E2 4F F5 E6 32 4B 49 82 B1 25 93 E1 D6 37 5F F3
 0B 09 CD 23 A2 83 AE CD D7 AA AF EB 91 B7 3E FA
 66 B4 C3 DD ED 6D 77 B0 91 1A 55 87 A1 3C 9E C3
 D6 61 99 46 FD 7A C9 F3 63 41 B6 B7 06 2C F8 1C
 8B 6E 21 F0 B3 BA A8 26 F5 59 AE 85 2B 72 E1 9D
 72 11 6A B8 CE 9F 6C 24 55 6D C6 F2 77 06 78 09
 02 FC C9 C8 7A 72 FA B3 9E B2 69 AC D1 4C 3D EE
 F3 3C 15 DC 18 01 0C 58 3C 68 A1 42 74 79 F8 54
 03 A4 D2 9A 7C 49 18 EC 07 FA 64 CD 55 5C 0A 0C
 CB E3 76 FB 5C 2B 95 F4 78 80 92 0F EA 80 10 E4
 69 65 6E CD 25 3B 3D 1A 55 9F F1 AB 5F 9B 8A 85
 1C 03 32 F5 C2 2D C2 0E EF 0D 43 DA BB BC 63 33
 ED 7B 62 95 BA 3C FE F5 C4 FA 32 22 A5 B2 BD 10
 85 19 92 67 D1 D2 70 99 C1 CF BB 10 FE 65 E2 43
 C1 77 94 46 9F 44 36 7D 9E 35 3B 49 CD 81 29 CE
 05 44 85 03 1D 00 82 11 7D 22 7B 09 2F 70 0C 24
 C7 FA 8C 78 B8 75 78 5B 6B 2B 2B A6 DE 67 BB F8
 68 25 69 60 E4 E6 4D 00 5F 30 60 10 D1 77 A7 23
 7F 83 0E AA 82 1C 00 7F 0C 42 2A FB 1A 76 85 6E
 CD B7 B9 6A 2F 65 B1 39 C5 A6 98 0F C9 C8 0A E6
 5F 8F 95 E5 67 E2 24 9A 7B 89 59 FF 96 F8 7D C8
 72 59 03 7C E3 7A 15 E3 3F B3 D0 2D 4A 1E 79 D9
 B5 FE EE 23 C6 13 D9 05 E7 40 56 51 9D 26 C1 C3
 2E 0B 82 2A 77 65 22 07 1E 44 FE AE 32 06 89 42
 AD 31 DD 16 D1 1B 33 1F FB 2D 49 8B 96 D4 A1 E0
 5C EE E1 1C FA 6C FD 39 7C 67 70 A1 AF 67 9B BD
 27 27 7D DB 2A 83 F6 59 DA FD AF 5A 26 02 CB 6A
 AB 20 AF DF FF 6B A8 40 37 98 40 2D 4C 99 E1 2A
 59 12 69 41 C0 EB CC 99 C4 10 51 C1 F7 B9 AA AC
 50 85 7D D2 31 DF 2D D4 2A 42 FF ED 90 7D 48 EE
 76 52 88 62 B8 63 F0 5C D4 26 88 4A 40 EB BA 59
 B0 75 A9 DF 0B 8F B4 8D 77 2C C4 F2 F0 65 40 EB
 75 94 07 1C AA D9 AE 46 2B 6D 27 0E 7B E0 DC 77
 5C 45 38 73 80 E6 AC E0 5A F3 E6 5A D9 06 12 EF
 10 0D 39 B5 AA 80 5A 7F 60 1E 92 BE BB 74 B0 0D
 42 0B 0E 03 B5 3F F5 76 7C E4 83 D8 83 59 D4 9B
 1C 5F 4A 2A 83 2E BB 21 F6 FB CB 43 BC 83 C0 34
 38 78 89 F6 3C CC 34 0B B6 AF B1 6E 91 2E 4C D3
 4A 6D 6F 9C 3E 85 08 35 BF 47 D6 D7 8E 01 68 57
 2A 5F 86 9E F3 41 24 BC F4 8B 39 2D 90 C2 25 99
 36 20 E7 74 ED C6 DE 51 4B 6C 40 45 36 F5 3F 00
 54 D8 A8 B3 C2 36 75 65 46 02 5E E0 4A E6 F0 A2
 7D F5 AE 27 FA 43 BB 69 24 16 13 3A 1B 0C 7F 00
 34 DD 2D 7D C1 A9 12 45 F8 34 01 97 07 21 7F EC
 A4 C6 94 00 51 13 85 9B E8 3C C4 69 39 8F D4 E6
 DB E8 EF 42 18 75 3C 51 0E E2 B1 1F 83 07 94 6B
 41 E1 32 C9 F6 DD A2 A2 16 3E 5C 72 F1 E7 85 88
 97 80 CC E1 0D 29 C8 B3 86 1F B8 F2 2A 83 9E A3
 84 F6 7D A0 C1 FB 98 E9 FC 5E 13 FC 07 71 96 4B
 60 C3 A2 2E 61 82 53 87 34 E4 26 5A 34 27 36 42
 4F 9A 56 45 24 BF 0A 79 C7 C7 19 24 50 A3 80 5D
 0C D9 24 84 5B A0 C8 83 C8 BB 7A 4F 6C 55 A1 BF
 6D FF 7B D7 29 DA B8 E9 35 E7 54 6A 06 D9 8A 10
 57 56 92 32 2E D0 E6 90 BB 58 21 53 24 4F DF 95
 2B D0 F1 B0 BD 2B 63 B3 45 97 A5 3B CA 23 AC 6C
 B8 BF 0B 60 20 98 12 AC F1 C8 98 C7 8A F5 23 1B
 05 94 F2 DB AB CC B4 02 CC EA 10 8C 49 E3 38 3C
 FC AB B7 CC 5C 5C A6 E1 98 8C 44 D4 90 5A 14 3F
 39 28 E2 DD 3B 7E 5C 73 EE D1 9D 87 E2 FD 03 3E
 63 0D 97 6E 52 38 15 0E 7F D9 83 26 23 BF 4E 17
 8D 5F 09 1E 1E A2 E5 42 FE 4E C9 F1 A4 44 CA F7
 34 5E 24 22 A4 1E 02 70 C3 F0 1E 80 B7 74 21 A5
 64 36 44 49 F3 6F A7 5A 6F 93 98 85 BA 6D D6 B3
 82 4E C3 F3 EA 8F 19 7C C7 2F 0C 61 5C 5A 67 43
 5E 13 4C 69 4A 0E 14 8E EA C1 E2 29 7E 86 CB 11
 A8 06 A5 B1 B3 4E E2 6A 83 16 55 DB 56 F3 11 E2
 64 EC FA 83 FC 6A 0C D9 A7 3F 1D 40 30 70 B2 2E
 07 E0 BB E1 6E A0 B9 CD 11 10 0B AE AD 56 1B 54
 1A F3 4A 91 26 E0 24 E2 CD CE 94 59 A1 D6 D1 B3
 0E EC 4C DB 8B B7 3B BF 71 7C F6 17 B9 12 3E 1C
 2E 76 FC 1A 01 0A BB 68 2E 54 57 2F 35 AC 1B 67
 17 09 53 12 78 71 CE 55 75 A2 58 EF C5 41 C3 39
 8C 3E F0 16 B6 F2 C9 03 1A 8A E7 33 34 90 A5 FE
 38 41 FC 96 CF 94 17 87 A6 E1 5E 01 2B 06 57 09
 CF 6A 18 07 DF 80 A7 D7 CA 8F B0 74 AA 2C 6F 4A
 71 03 BD 6E E6 D1 9A 6E 48 9B 4E 69 21 60 09 A4
 58 4A 3F 2B DF 18 08 2D 02 60 04 B4 16 31 4A B0
 74 D8 D8 66 02 F0 18 1E ED A7 03 01 49 0B 9C 72
 10 0C 23 AD 40 04 6A 58 EA 18 E7 48 AC A9 84 15
 F5 D6 DD B1 5E 63 EE 52 17 4C EB E5 A2 26 BD 3B
 64 D0 B9 F8 DF 40 FE 15 00 95 36 F0 83 92 2F 0E
 6C CF 57 0B 1E E5 7E 3E D9 3A 9B 55 D7 5C CA D4
 AC 9E 4E FF 85 31 64 C2 0D 6C 18 69 B7 71 43 0A
 79 06 36 BB 55 AB 22 03 60 75 42 AE 25 4F A1 7A
 3A 96 B3 A6 89 E8 F2 E6 24 FC 44 44 F5 40 77 A0
 2A 65 BB F3 54 92 16 64 17 E8 68 66 4F 4A 94 8C
 84 A7 42 92 2E B6 A7 F3 69 CB E3 29 62 AE 1F 5C
 3B 40 C7 26 C7 A1 DE FE 4A 0B 4C C5 8C 68 94 4E
 DD 84 D4 B5 69 CB 61 12 9E 8A 53 E5 4F E1 D4 E4
 75 77 22 F5 90 55 5A D0 8E 43 35 47 53 27 1A 5C
 BE 5C 7E 37 A4 C4 3B 18 A3 0E 8B BA 1F F0 CC 05
 69 A5 E8 0A 54 6A E9 B3 0E 1F A0 21 36 26 95 D1
 D4 E4 E9 D5 FD 1E 68 2F 13 DF D7 2A 22 F8 84 AF
 98 0B FD 55 A0 72 41 A1 DA FF B6 71 92 19 1A CF
 90 74 FA 12 03 1B 55 6D 3D D0 DA 43 45 09 31 6F
 89 7D 9E 73 6A 1C 6A 5C 05 72 27 CE 69 A7 74 67
 10 E3 E3 64 ED 7E D2 55 C0 B1 34 2C CA 8F EA F7
 2E AA D7 2B 6F 19 C2 90 1C 54 FE 96 5F 55 9B 18
 6A B5 84 8B EF 16 DD 37 7C CD 77 A5 E6 AC ED 92
 D7 64 F7 89 59 7A ED 8F 60 1C A2 CC 10 20 27 3B
 92 A6 A7 27 9B 45 12 A4 98 6E E1 91 61 5C 0C 28
 00 59 34 75 DC 5E D4 86 FB 58 55 33 8B EE E5 9B
 EE 90 B9 2C 93 39 D4 EC BA 7F 59 45 8E 0E 7D FD
 AC AB 5C EA 00 C4 4E D4 3F 14 EC 19 CE 07 AD 60
 5C 3C 30 AD 6C 2F BF 5D 14 31 B6 E9 F3 12 53 97
 4F 2F AA AC EB 9E CC 43 0C 53 B6 94 ED 86 6C F6
 94 CB DE 11 D5 75 CB 03 24 90 F9 67 02 E9 A4 50
 C0 D1 DA 9F 5C 37 19 0A 68 FD 7E D5 25 21 9D 21
 14 C8 5B 29 EB E1 94 0F D5 FD 6E 07 4D BA C8 F4
 4E CD F7 AD C8 52 3E 55 39 4C 10 39 9F 30 8A 29
 B6 D8 73 FB 1B 2B 1C 39 D2 79 B7 A2 45 20 A1 CA
 E8 6D C0 32 DF C3 6B 2F E5 39 E2 FE 09 F5 0B 05
 DA C2 80 BD 20 D6 F6 5F 25 11 4C 59 9D 0A 11 9F
 30 3A 36 E3 9E 4A 1F 46 A2 32 FA 68 F7 34 22 17
 6F 26 62 52 9C A2 E7 10 C1 BB FF 45 11 11 9C 74
 AD B8 92 7D B0 4C 69 92 33 2B C8 0D 87 7B 1A 68
 E6 31 DC 34 CE 22 46 4E 00 AE 23 0A 06 12 50 0F
 10 E5 97 7C 47 C3 3D EC 78 0B E9 33 77 BC 0B FD
 80 E3 13 9C 4D D9 DE F9 7D E1 34 6D A4 43 D3 F0
 52 A6 87 EA 9E 0E 46 09 F4 A0 3B B3 45 8A 47 82
 8E 68 73 05 BA 8C CB FA 3B B8 CA DB D7 6D 27 C4
 87 72 2B E5 37 D2 8B F0 49 DA 77 25 56 D2 15 44
 D7 22 45 DF 81 FF E0 5B EF 77 5F 65 83 F7 C2 8B
 6A F5 AF 40 12 51 8F E0 83 91 A5 E3 80 5C D7 F7
 0A 99 C8 5F 60 BD 4D 1B 33 D5 53 1B 2B 93 08 56
 10 3F 81 18 C6 1A EA 3A 96 F5 68 B3 33 9D D6 4F
 0F E0 A9 47 4A DD 15 76 66 A1 44 11 13 81 A7 D6
 52 05 92 D5 28 B4 97 C7 D9 49 A3 9A A4 19 86 29
 ED 32 12 1E 17 FC 47 2B 38 50 3B CB A1 E2 F1 36
 35 E7 44 49 A2 D9 FD 01 D8 4C AA 0E 45 7E C3 FA
 C2 D4 82 C2 66 02 A3 0E D0 76 2A 7F C5 5E 03 8D
 46 C6 36 67 38 18 24 8E FB 45 AE AF C6 6C D4 DC
 FA 75 32 0C E2 E8 0C 5D 2C 37 24 C1 60 C0 7B C7
 35 56 03 44 5D B6 96 45 22 40 83 E7 1E 69 4E 8F
 2D 67 61 80 6D 92 6C FD 71 F0 6F 88 D4 0E D5 56
 8C 43 B9 A3 DF D6 59 93 1E 9E BC 43 E6 4A 5D E1
 5B 2B 2C 32 AE 66 DD B5 DA EB 3D A4 97 E8 C9 E1
 FC 96 82 57 A2 D1 7C 7B CA 22 68 45 42 4F CC 1A
 30 47 0D 24 0D 41 7F B0 B6 30 8D A8 26 7B 5A 8E
 0B B7 B9 51 FB E7 43 17 F3 78 AB 17 5D 5C 95 E4
 64 94 B2 79 3B 31 95 6B D7 65 03 93 3A 56 FB FD
 54 F9 2A E8 40 82 FA 73 C6 72 1A 10 F2 81 E6 FD
 BB 8A EB 09 8C 30 07 B4 01 71 C6 5F 87 3E FC F6
 DB D4 ED AB 62 0D 58 0F 39 8B 92 0D 5B 96 9F 74
 02 69 0A 55 BF 0F A0 28 A8 08 EF E8 14 2F DA A9
 9C 5E EB 87 B4 39 77 56 42 EE D4 A6 7A 80 AA D5
 01 55 09 C7 33 DC 94 FB F2 43 6C E4 7C 9A C7 F9
 C4 05 3F 33 34 A6 64 C6 EB 5F A0 CD C1 FF DF 61
 5E CB ED EF 00 45 9A F1 C0 BB E5 82 AB BD 2F EB
 78 60 0E E4 61 71 95 17 8D 45 B1 DC 6D 22 63 B3
 82 32 E6 6C 7A D0 6F AF 87 FB 7D 2D 2A E2 3D 8B
 AE 6D 5E 49 F3 E2 97 8A 89 7B C1 24 93 17 70 48
 71 5B B1 98 17 52 C2 82 6D E3 5B 21 E6 00 B2 F7
 5B BE D5 C3 7F 81 1A 6A C7 02 1B FC F4 C7 25 77
 0B CC 8D 33 FB 5D 15 4E E0 56 B8 37 2F 38 17 CE
 D3 BC 94 CE ED A2 A2 56 B7 8F 4C 41 16 EE B7 5F
 D5 35 E2 86 43 50 54 21 7E 8A 18 18 E6 01 34 FB
 59 A4 E2 24 13 80 17 37 01 5F 0A C0 F7 29 01 A5
 20 AC 7B 3C 10 B7 5D 81 8E 01 C9 1D 81 B8 AB 81
 C7 C0 6E 2E E9 47 28 40 88 94 5D 37 13 0D 1E C2
 87 8A CD 16 6A EE 74 0C 6F 16 89 F2 27 83 75 10
 38 A3 08 B2 BE E6 7E 8F A0 94 4C A2 BF 17 0A 37
 F4 ED 86 F7 93 B9 54 44 F6 5C C2 FE 63 30 F3 EE
 3C 8A 9A 76 00 93 5D 6E 4B B6 82 5B 18 F5 A0 7D
 D9 EC 93 5D 79 EC 64 FA 66 19 F8 95 3E A6 15 21
 03 83 A0 4A 14 BF A9 D2 CF 05 4E 3B 89 18 76 1C
 B9 41 B6 48 95 4C BA 34 E4 F1 41 40 73 7D C5 9C
 6A 9F A4 77 55 F5 C9 8B 23 02 0A A2 C1 7B F9 00
 5A B8 CF 45 05 C8 F3 43 2D B0 BA B8 4D 06 4E A2
 65 EB 35 51 14 D5 08 13 5D 39 CA 4A 0C F0 38 4D
 91 15 84 DC 62 27 74 60 65 3D 7F BF 7C 3C A3 B8
 2B 8B 3F 54 66 70 89 EF 32 9F DB 6F 9C E1 E5 70
 E0 17 A1 F5 CB 10 48 88 7F 23 10 B6 89 DB 54 33
 69 56 CC F5 C1 D8 59 B3 1E 66 DB 58 31 EC 6C 7F
 77 8E 41 FE 7B 43 1E 7D 24 5F 11 5C F2 9A AC 61
 DD 99 09 08 DD 30 FC 13 F9 1A 18 EC E3 02 A2 AD
 A4 20 CB D6 D0 0A 39 40 61 AF 1B 99 73 46 94 50
 AB C4 4F B9 3A AA E6 D2 BF E0 3F 35 DD C6 4C 99
 4D 18 23 36 62 4D 3A 97 83 5A FE 91 99 1A 26 3E
 56 80 2C B5 9C 33 6C 51 6D 5D CA 5A 82 BE B9 FE
 9A 10 D7 FE 45 88 6B 9C 96 00 0F C8 2C 1D 2F 0C
 65 E4 46 2E BD 96 76 1E 5A B9 DF 08 B8 D2 57 FD
 20 58 21 C3 B9 D8 76 0D 4D 5D 9E B1 D8 EA F7 11
 83 1E DE 3D 57 E1 FE BD 8D 03 4C 86 C6 07 1B D4
 AB B7 0F EB 1B 97 9D 61 6E DB 4F 54 CA B0 E0 55
 AD AE 64 34 9D 5C 86 A6 AE 60 03 C2 BF 60 56 EA
 EB 97 3D CF AC D0 8C 9F F2 F5 F8 1A 69 04 D6 A9
 85 D1 F5 C2 CA 00 EE 3C FF 7F E9 1E 91 4C 8E 1B
 9C 5B E7 4C B4 75 64 CB 1D B1 C7 96 71 9B FB 37
 18 90 B9 19 72 4D FC 73 24 18 C5 90 07 BD 7F C1
 77 C6 5A CE 5C 1F 4B F8 30 C1 7D DF 1B B5 16 FA
 3B 21 46 35 8A 68 C4 A9 17 32 DE DA DF CE CE BA
 6B FA 63 D0 EE 21 4C 05 C4 B8 C5 9B 15 69 ED 69
 38 32 72 9F 10 9C 37 10 7C 5D 14 1E 02 49 8F 90
 EA 1E 32 5C 28 72 3E DC F6 A8 62 F8 9A 9C 86 B3
 7F AE C6 A7 57 C2 B4 2D C9 90 FD C6 32 4B 9E AB
 24 5D C0 06 CD A9 35 41 60 5F DA 2A BB D4 B3 3B
 9E 9B 8A 9E 1F C7 A2 67 8C 92 5C CA 42 F7 66 64
 45 40 4C 14 D6 8D 78 C4 8D B2 6B 89 9D 50 91 BE
 66 A6 E7 52 BA B6 B6 E5 F7 52 7B E6 E7 FD 42 F4
 9F F8 78 B5 AC 3C C9 B1 ED 61 8E CB DC 6B 7C 5C
 C6 57 05 6A 1E 04 23 0B 80 31 32 96 76 66 61 52
 D1 F6 9C 13 D2 6A 98 19 EC 15 A2 06 BE B9 18 56
 BC 1B DD E0 E1 04 CE 6F B1 72 60 29 D5 1B A7 30
 9C A7 3B F2 60 1C 03 F1 6F B3 A1 A9 6A 34 4D 1F
 6C E3 EC 01 20 B2 12 85 89 B3 BE 0D AB 1F E6 12
 52 28 4A 7A CA 3E EE D8 E9 66 57 D2 8C E0 E7 26
 14 D3 DD 4A F6 F7 94 B1 BA E3 FE 69 78 AB F3 4F
 C1 E6 DB F0 9E 8D 7F 31 93 C8 6B 0B A0 12 A7 60
 BD E6 A6 DF 84 FA D2 2B 2F 5E 04 D4 57 26 48 1E
 5D E8 1A 58 E6 F2 39 65 0E 37 22 C5 96 D5 D9 56
 C5 90 E5 D5 6B 16 09 27 E6 74 BA A8 32 E7 86 80
 6B B4 A1 E4 22 47 8B 0B 21 0F 40 4C 45 C2 E3 7A
 13 25 AB 07 C0 95 A2 C6 55 64 56 47 B3 8A DE C8
 E4 85 BC A5 2E 13 1C 12 C7 14 AE D8 8B 87 32 A6
 26 E3 F5 69 C1 08 09 49 F9 5A C0 E4 4F 00 8D 16
 D2 37 13 A6 F4 91 F4 79 D7 13 6B BB 0A 0D 90 0E
 1F DC 4A C3 10 AB D3 BD B6 5E 44 E8 D5 5A 6C E4
 3F 0E A3 3A A7 AA D8 E6 27 DB 3E 76 F9 C9 C8 82
 1A 7E 3D C3 6D 81 62 BD E0 98 33 88 BD 60 BE B9
 67 31 9D 4D F2 66 A0 04 08 C8 50 81 1A FF 45 F5
 18 2B 62 12 16 E4 0C B3 20 91 9F 5D 83 CA FD 76
 51 98 18 60 73 70 3B 8B 7E FA 3C A7 D8 14 9F 64
 F2 15 FC CA 6C 2E E3 9D B3 F4 43 63 1E 51 08 A5
 80 94 E3 9D BF F8 AD 92 D0 5B 6D DB 9B F1 EE FD
 B4 52 86 01 2B 4D 80 35 C7 C5 A9 AE 10 BF F8 77
 15 9C 2C D0 11 60 65 27 C4 D4 AB BF 79 D7 E7 B5
 F1 7A 8A 27 82 04 AD 9F 2B 3E F7 14 B0 85 90 A6
 E3 EF 4F A4 20 B9 8E 6C 2C F3 D6 C9 3C 17 E1 0D
 F4 8B C8 F2 6B CB 1F 20 87 26 06 FF CA 01 89 E1
 9E D6 5F B0 A5 5F B2 D8 57 86 53 0B 4E A7 15 DA
 B0 F2 4C D8 3C 68 90 08 1E D9 49 2C EB E8 52 35
 23 06 7F DC 66 51 63 49 4A 78 82 88 D0 9F BC EC
 3A 85 03 21 EB FA A3 07 2F B1 BA 84 87 55 76 94
 0F 56 C0 B5 E8 A1 E6 C2 14 46 BB 94 EC 4F FA F8
 CD 48 DF 43 76 EB D6 BE 69 A2 A1 17 6B 31 6A 89
 2B 42 F8 1A 6F 98 46 25 70 84 8A F8 10 30 E9 20
 01 1D 8E 5B 3A CA 43 05 C0 AA 82 ED 31 E7 D4 52
 D2 67 62 FB 3A 62 72 D6 37 C8 62 81 D7 67 4B 48
 20 CA B5 8C 95 98 D3 9E 88 82 04 DB 6C 74 C3 E8
 88 36 2D 35 47 93 4F 93 51 B2 81 AB 0A F9 A1 0E
 21 01 A7 78 C8 8F 46 98 45 7A 6B 52 8E 9E AB 2C
 96 8B 14 49 9C F9 18 BC 07 04 69 65 C1 54 75 00
 05 7E 5F 6C 4F 85 04 C7 32 03 44 3B 26 7B 5A 02
 D7 D5 F1 AB B4 82 9F 28 76 CB F1 96 37 03 4A 0E
 A9 0E FC C1 2D 6F E1 85 BB EA 0F 0C 45 0C 1C 4E
 D8 C6 E8 A8 02 88 EC EE 6F AE 64 74 83 22 92 F9
 69 89 BD 99 C6 E5 B9 29 FC 12 B2 02 2C A7 62 CA
 7D E3 D5 2B CF F6 99 DA C2 F4 47 B9 D7 6F 7A D2
 E3 47 71 D0 B4 43 44 49 DF 54 63 FF FA 28 11 72
 26 13 71 82 30 71 9C 35 4E 80 95 1A 29 9E C2 B5
 72 D9 4C 83 CA 69 01 FA 7D CB 74 D3 17 9C 16 0F
 34 D9 B1 97 0A 09 A2 D4 95 A3 12 86 80 E8 BF 99
 42 2F CD ED A5 BC 34 13 B9 EB 4C C0 F8 A0 B1 DB
 92 CA 89 A3 88 E6 CE BA F6 EB 17 58 6E 4E 7F E2
 F4 DA CD 50 E7 9A 91 DE 9D 77 CE 05 E2 73 60 60
 04 90 0D 44 06 5D 68 BA D1 B0 F7 65 A7 CC 61 9C
 C9 4E 9F 36 18 21 9A A8 82 DF A5 1B 59 71 74 48
 13 2D 86 6C EF C5 B9 60 44 9B 2D 97 30 71 E4 6F
 9D A5 4F 7D 29 65 38 4C 16 3D E9 B3 2A D7 3C 87
 59 0C D9 45 0F F9 D5 87 F0 D7 D4 49 7A 11 C3 CC
 39 57 07 75 2C CC A7 84 04 AE E4 03 E0 3F 3B EF
 3A D4 AB EC 5B 87 D6 3F B0 34 67 63 24 EE D3 4C
 A7 3E EB 80 89 3D 0A 25 C6 F8 D4 0A B6 8E 8A 6C
 6A 01 1B C5 95 D9 2C BA 58 39 01 A5 43 1E 98 73
 3C DA D6 06 23 84 C0 A2 E0 25 4D 5B 2B 4C C0 32
 73 D3 C1 5D 56 A2 67 03 9E E2 FB 6A 4B 4C 29 C0
 6C 16 32 84 B6 23 A8 90 0C 3C 86 DD 7B 84 D6 FE
 6C 0D E4 9A 8F 69 46 48 2C 7E 17 81 3C 7C E8 26
 97 83 88 CB CC 1F 3D 35 A4 F9 32 EB 44 C5 C1 5D
 5A 4D D2 9D DE E7 9A 3D 7D 06 20 E6 38 65 44 51
 5B EE 66 5D 7B 8D 2A 3D 90 33 31 55 DA 85 88 AD
 56 08 69 ED 65 60 FD 2C E8 90 43 2E E1 7F 28 9D
 A1 48 EF 04 D5 5C 2A F3 00 C3 4A 9B 10 5B EE 25
 94 16 E4 F8 75 3D DE 5E CB AB A5 CB 9E D1 07 15
 29 1D 1F 06 A7 86 7A 5A A7 2B 14 4C 46 7A A5 07
 F0 82 15 63 A6 B1 38 A0 89 9D 12 39 17 EB AC 16
 89 13 97 95 43 06 88 F2 60 D3 20 50 A1 EC 1C 4C
 75 A8 AB CD 8C 2C 33 DF E2 CC 7D BC E0 2D 2A 0F
 E8 19 D6 96 4E 8E BF 2D 45 D6 0C 39 22 D1 18 BC
 03 0D CB 64 90 70 C9 98 76 EE 61 CE E4 D0 CB A1
 B3 F2 C7 D5 A5 3F 57 0D B1 31 7F 6D 48 39 23 C7
 84 FD 16 58 31 46 D6 66 ED 55 21 F9 F1 5B F3 EC
 6B 4A 71 08 54 60 91 01 73 56 87 B8 22 62 D2 4B
 C1 56 99 C6 B5 EB BC 27 84 47 3D 4E 5A 88 7A D4
 67 8F 68 29 36 13 FD 31 A9 3C 7D D8 5E FC 3F 83
 D7 8D 25 E1 C8 67 D6 A2 EA 8E 5F 1C 07 97 25 BC
 52 0B BE 83 48 72 8E A1 85 41 93 54 1A A0 10 46
 E8 9F DE D3 2D 34 52 8B AA FC 37 60 14 06 53 00
 C0 15 93 F0 A7 5B 69 F5 89 4C 5F CF 00 9C 2A 15
 62 1E F1 DC 28 68 A7 F1 70 86 ED 4B 7F 8C AC E3
 2F 33 1A 05 17 30 9A C9 9A 13 6A DC D9 58 BC B3
 58 B2 32 5D F2 52 9A 8D 31 B0 10 D8 D6 F4 DC 5E
 60 0B D8 CB 55 66 EF 30 C0 47 94 2B 10 FE 82 7D
 48 FB 69 80 5E D1 9D A1 0D 65 BC 6C 67 11 07 94
 32 98 0E 60 EB F3 B7 C7 7F D3 C6 05 B1 53 C1 DD
 76 B1 32 44 B8 31 37 47 12 1A C4 47 17 DB F5 2B
 AD 77 47 6C CE D3 D9 9A 8C 72 0B 19 A3 1B 55 19
 43 33 21 34 17 49 2E 49 35 F2 FF CA A3 4F 72 93
 18 AA 89 5A 14 8B 0C EB 35 63 78 0D 2E BD BA 84
 3D 01 D0 A0 AB 6E 8D 55 5F 87 6A 88 36 D5 58 9D
 14 A3 2F 87 3E 89 25 CA 8A 41 80 F8 6A CF 4B 75
 CC 78 D5 75 E5 EA E5 51 25 70 03 01 A8 21 8E 25
 C1 9E A8 8D B7 4D 74 C2 67 0D D2 0E B8 85 82 34
 EC CF 6C 4A 6A 54 A7 AF 5C FA 43 60 A5 C0 79 CA
 5B A6 D1 E7 F9 C9 A8 C5 86 36 F5 E3 85 AA 4D 08
 C8 C9 4D 78 04 30 68 3D 3D 6B 8F 56 13 97 D9 FB
 F6 B5 25 69 3C 63 CA FA 91 9F 3F B8 D5 23 3B BD
 A9 27 20 91 B8 C7 DF 5D 88 A2 D7 6A CA 29 5E 81
 5A CF 19 66 C3 6D 9D 1A 38 4F F3 CA A0 68 7E 4D
 E4 8E 12 72 01 EF D6 5B FB 5B 3D 0E 7D A2 B5 2C
 E4 B6 55 93 CE 65 BD 63 22 A2 19 CC 5F 8E A1 15
 50 CF 7F 4F F0 68 36 A7 63 47 78 BF AB 63 84 4D
 5A B1 F4 BE 1B 28 7E 7C A7 3A 9B 80 3A 89 8A 48
 F2 14 9D 85 16 A2 77 BA 17 5D DA EE CB 3D AC 5A
 2C 1F C5 4E DB 7F E8 FB BB 6E 89 7D A4 8E EA F2
 F6 F4 FE 37 C2 6E F7 D8 28 32 53 DE 17 AD 2F 0E
 D2 4E 8D 98 EA E8 1F 91 16 A6 2C 75 1D 43 6C 8B
 67 7C B1 7F 1B EF 25 8B 25 A4 DF 87 FB 81 34 8F
 62 0D 9A CF F8 B5 7E D1 E7 4F 45 04 50 7C 82 8A
 D8 F3 EF F2 97 BB 74 3B 22 49 CF 2D 12 4C 3C C3
 48 88 DA 5A A9 9A 5D FC C1 58 7F A7 2E 1C EF 2E
 27 2E B2 AE 0B B5 78 89 60 8D F3 36 9F 14 FA F7
 05 47 5C CC EE 93 75 E9 D9 AA 4C 7B EC 23 62 FE
 3B 48 12 AC E4 61 09 E0 17 48 0E 90 F3 60 65 3A
 3F EB 9A C0 C8 51 C8 0A D2 C7 F3 87 44 D2 D5 E9
 BF 36 1B 49 A9 4E 3B F7 52 F4 54 BE 84 D3 F9 05
 6F BE 64 6E C8 B8 AA 07 D7 44 24 91 75 A1 B5 1E
 87 92 4C 49 1B C7 6B E9 4C 31 AE 56 1C 2E EB 0B
 65 D6 21 19 4A 44 5C 56 EB 4C 7F F5 28 C7 43 D0
 A7 08 19 5A 5C 01 D3 8E CC 47 B4 5D 41 69 28 2D
 51 79 10 0B 8F 21 DB A6 1F 25 E1 B9 98 61 AF 95
 42 64 D3 C8 2A 48 8F 62 3D 61 34 36 88 43 F4 E1
 FF C9 5C 03 F2 07 8D D5 63 C1 6D E2 AC FA 74 8C
 01 90 A7 53 35 26 E2 5F 6E 42 1A 8F 1D F1 0A 9D
 E9 BF 11 4F B6 AA 17 F7 60 BA 90 AB 27 5F 7C AD
 C9 55 90 4C 86 FB EE B1 4E 5B 59 71 30 05 F6 9E
 2A A0 66 BA DF B1 AB 74 F5 0C 32 A3 90 BD 0F BC
 56 01 9D 97 BE 0C 48 B4 70 CA 9B 89 96 A9 8A 8F
 0B 53 42 68 71 CC 7F 10 0F D0 09 AE 25 93 48 C9
 96 07 F9 DD A2 14 4F 98 7A 12 91 24 6C 10 2F 31
 36 24 06 BD C8 3E 80 BE F4 C8 69 4F 6E 4E CA 14
 14 E4 EF 9A 7C 70 D3 19 A1 44 A4 E9 8C 41 A1 19
 CF 32 0A 97 67 69 28 24 80 57 8A CA C6 1D DE 01
 A9 6E 05 80 41 0A 63 3C 64 58 1B AA BE 01 AE F2
 F2 9B C1 7F 47 13 7E D3 10 91 6B D9 0F 50 C0 8E
 FE 9E 68 E3 64 0A 63 4E E6 C9 F5 CF A4 39 79 B2
 65 15 27 F9 C0 17 5D A9 47 57 B7 07 70 7D 89 AD
 A5 5F 62 AC F2 BE 90 34 CF 65 61 37 F2 A7 ED 28
 67 56 76 2B 03 B5 36 A7 88 75 6B 69 3B 15 3B 02
 DC DC 4C 4A 93 60 4A 83 5C 80 EA 74 1D 20 12 71
 62 FD E9 50 33 C2 58 22 56 0D 29 FC FF 7C FD 95
 06 ED 9A 52 C9 46 05 C3 51 94 80 D1 16 02 6A 7A
 12 1A 8D 47 66 40 FC AB FE 8E AD 95 A2 79 48 4B
 0E 1E 33 34 C9 69 B5 A7 8E E2 B2 08 9B DA 30 6B
 E1 BF 9E 58 27 35 18 AB 86 40 AB 09 37 E5 D7 0C
 86 D8 8A EA 70 19 5F 6B A9 C1 24 CB D2 85 C3 21
 1D 63 3C 53 2A CC E8 44 55 FE 71 DB 63 72 3E 5F
 FA 7E 15 89 BA 42 FC 39 34 73 21 B4 92 68 67 85
 3B A1 59 96 E9 A4 EE 75 98 B4 74 F8 AA 36 34 54
 3A 35 1F 28 AC 35 AD C8 32 13 2C C3 36 C2 65 5A
 C9 E0 8F 76 60 FD 90 C0 BD 5D 03 81 E4 D5 B3 3F
 CA 20 75 76 1A 1C 41 D8 8B 39 DE 47 5E 0D 03 9E
 B8 D7 94 BD 80 40 8B 7A D7 0E D6 21 80 5A FF ED
 76 8A E0 B4 75 22 90 F4 8E 2A A6 20 EE 3F 5B 45
 D2 36 68 1B 86 80 19 F0 D2 C2 E7 CB 35 0D 52 19
 84 E8 25 4A A7 4B EE 05 CA 4D B5 15 B9 F0 10 06
 51 02 3B 89 B2 27 41 02 F2 8A BC E8 75 88 1C 54
 F8 73 2D 47 BD 86 8D DE C9 84 46 B2 DC 02 35 7B
 8B 23 7C 44 2F 41 E9 13 A5 0F 13 7C 69 4D 70 39
 9E B0 7E 1F CF 67 3D A1 4F 0C C9 61 12 45 9E A0
 F9 5F CD 85 DA 5A 35 12 19 36 8D F4 83 1B BD 28
 12 67 10 7F 48 9E 45 55 00 56 79 AA 6A 84 4C D2
 79 D1 86 5C 2F 49 AE 2B 01 A8 27 5F 49 CB A4 CC
 A7 FB 07 89 AF 9E C7 BB A7 98 BD 86 25 19 3A A4
 81 C5 07 9B 34 31 9E CC AF DF D9 06 EF CE 8E E3
 90 0B 68 5B FE 7E E5 88 01 06 2C 6E 05 DF 40 F5
 B4 8D 8A E7 E1 BA 4A 67 81 71 DA F4 B5 5A FA 02
 78 DE 9D 33 F8 86 4E 8F 6D A6 83 91 CE 47 B4 86
 4B 7A 13 D3 EA 49 0E 74 86 D4 AE F3 5A B7 90 02
 29 62 D5 06 92 D7 15 B8 D0 5B AF 68 C2 1F 23 69
 B5 BB D6 B8 AF 6D 21 57 C5 82 98 3C E8 D7 3A 95
 54 2B FA 1E 61 42 C1 17 68 87 01 00 5C 66 6F CF
 BB 46 04 39 51 CF 73 4E 04 28 8B 21 D0 B0 C9 AA
 64 E4 D7 90 26 68 62 4B AC 7B E4 6B 51 66 9F 22
 76 59 C4 FF 2D EA 06 F2 D0 88 BD 61 26 13 A0 7B
 8B 18 0E B9 54 AB 63 52 8F 6A 55 9C 68 F4 D7 2C
 0B F6 FA 91 F7 EF AD BA BB CB 3C 85 14 81 EE 1C
 96 A8 CA 92 C0 55 E0 38 EB CF 6F 75 94 E6 45 25
 94 D3 F1 86 57 E7 51 9C FE F6 07 9C 92 FD 19 15
 C5 48 5A E0 53 2E A2 FC 46 63 5D 42 0B 3A 37 75
 D7 C4 B7 D5 B1 ED 2D DF BA A3 F9 31 18 0E CB 51
 34 49 92 21 1B 6F EC 1C 78 CD 03 86 F5 40 92 E7
 DD A1 6B 72 52 76 29 30 7D 8A 4B 20 65 AE 83 2F
 F6 2C D4 10 7B 6B 05 D8 C0 EA 6C DD F4 65 B8 79
 08 D2 9D 3B DD 55 0D 82 98 86 1A 79 4C F9 3C 8A
 8B 1C C1 E6 AD A4 ED 88 F0 41 19 28 80 28 9E 0F
 4D 12 C6 D7 3B 46 FE F7 26 3D 08 66 F5 C2 9A C6
 5F 56 56 3F 2A 81 53 7A 06 D1 B5 ED 03 59 20 1C
 5E 32 DF 9D 98 D1 1C 92 5F E3 6C CF CF F8 6D 3A
 C1 2B 5F AE CD CF 2E D1 A1 82 A3 D6 BB AA B8 B1
 0E F1 70 9F 19 D9 4A D3 C5 E3 46 42 58 A7 FD E6
 5E E9 4D A1 1F 30 D9 C7 79 8B 79 A7 57 13 ED BD
 CD 99 D6 6A 27 97 46 E2 46 33 96 81 28 B4 A7 4A
 2E 0F 9D B2 ED A3 83 D1 02 BB FC 77 AC 6C EE 5F
 04 3F 7A 9F 93 5F F8 BC 94 65 24 B8 F5 B3 8D AE
 98 6E 55 D5 98 E5 91 E8 B4 45 B6 BB B6 16 12 62
 50 55 AE 13 AC 0B E6 49 43 F7 CF 78 56 F3 46 16
 88 DE C7 49 F4 44 87 4A CF CB 87 8E 7E A1 7B AE
 C2 23 22 76 BC 9A 3C 33 BD 1D 1A E1 F4 3D 1B 6B
 4C 6B FE BA F2 6C 13 15 20 3B 58 7D DB 1B F3 6D
 D2 B9 6C 0F 66 C1 B1 59 1A D8 4C 07 D2 70 1A 6A
 38 C5 6A 26 3B 99 8F 46 E5 7B 62 FD 67 C7 BC 26
 A6 EE 15 D6 4E A8 9E 1A 59 F3 40 25 57 64 A7 8E
 7D D5 DE D6 22 7D 5A F9 5C EC 37 3E E8 68 C9 09
 5C ED 22 56 C0 A3 44 72 0C 7C C2 0D 05 42 B4 A7
 D3 D8 C3 F3 85 30 A8 F5 AB 6F CB 5F 2C FD 91 B4
 A7 04 28 61 6C 5F AE 20 48 ED 66 7E 7D 48 A5 8F
 7C D4 35 C4 6F 23 BF 24 F0 6E BC 85 89 37 5C 40
 F5 01 14 F7 FE 15 D7 58 94 12 0B CA 82 C7 84 F8
 86 7F D7 62 83 E4 8F 83 72 1E 42 BE 86 E7 F6 A3
 A9 EC 4A 0E 45 A4 F9 77 4C BB 8C 39 9B C9 F8 A2
 51 C6 A5 DF 10 2D 2E E4 B6 FC 56 3C 50 78 93 04
 8F 52 29 64 0C 02 F7 B0 AA 83 1D 3C E3 C5 E9 C5
 C5 90 D8 A4 CD 9A D6 30 74 F2 2A C8 F1 F0 DE 7A
 1E 3D 81 69 CD 97 CE 02 9A 8A D0 02 F1 65 E8 8A
 9F 0D FC 09 3B F3 ED F4 23 1F 61 34 63 00 1B 26
 7C EB 98 E6 C1 EB 22 B8 14 C7 D1 E0 2E 97 B3 15
 75 19 90 91 4F 19 A8 01 C4 72 CD 7D 59 C3 9B 92
 01 64 AA 10 B5 45 7C 73 C3 F7 7D 6D B3 DD 62 6B
 59 CC EC 18 7D 7F 5B 28 5A 22 FD 22 42 E4 74 6C
 F0 66 82 88 4E 14 29 C6 E3 95 BF 4C 51 41 A9 16
 56 1D 88 55 ED 85 39 2D B4 1D A4 19 E6 38 5C DD
 9E B6 01 2A 54 AC 27 D3 80 F8 E5 40 55 96 75 6B
 05 A9 B6 7F 17 FD 67 6F FF 8E 43 71 CC A5 03 78
 7E B4 F4 AE 85 F8 59 5B 52 50 BB CE 01 F6 2B 49
 BC 6C 3E 00 09 91 C8 1E 5C 05 80 F0 C4 39 AE 2D
 7B 82 5C E1 08 B4 C4 2C 47 34 60 44 55 74 F4 B9
 79 72 97 3B B8 A3 8D 9B 0C FD 69 5E 23 67 4E 5D
 4A C2 F7 BD 25 43 06 8D 84 7F 55 86 EE C7 B9 2D
 A5 B9 64 0F E7 5B F5 71 B4 66 AA B6 7B 57 BB 68
 B3 4A 2B A5 75 4E 06 73 6C 0E AE 82 B7 B8 0A CA
 E0 B2 12 67 69 D4 D8 63 73 0D 86 AC 0A 1E 9B 7A
 5F 38 F4 98 AD A7 EC C5 D7 AC 6D 40 ED 86 80 34
 AF 15 A2 9E 88 A2 D6 07 9E 5D EA 7D 51 12 E4 08
 79 F0 07 C8 37 26 C1 55 41 B6 F8 5D 1D 4B B1 2D
 A9 47 EB F1 D7 B9 60 7D F8 97 6B 8E 17 1D 9A 85
 AF FA ED 2B E6 0D 52 78 8D D0 4B B4 0A 17 70 F2
 D2 0A A5 A1 F8 DD AD 1E E2 63 1D D2 97 85 2E 95
 42 EC 38 F3 AC 9D 5D 4B 45 C0 5D F6 33 23 E0 96
 C5 72 E3 9F CF 3C E6 CA BA 50 5F 20 60 10 9A BA
 AE 85 22 DA 53 29 EC C3 10 4E 68 5D 7F C7 B6 5A
 9B E9 5E 90 72 79 09 FA 29 B1 1D A8 91 C5 74 E7
 98 4D A2 5B 38 B8 51 D0 00 82 48 DD 0A C8 0C FB
 B4 55 74 D0 B8 77 0A 0C 03 9B 4D 1F BB 7C 3B 78
 CA 6D 44 92 78 AA D3 D9 05 BA 70 6C 0D A3 FA C5
 CE 1A 1B 3F A3 FC 55 11 B0 96 45 44 CC 88 6F 78
 4A 53 A2 87 88 E4 CF B7 33 EE 4C 9A EC 2B C6 61
 64 DB 31 3B F2 1E AF CD F5 2A 54 B9 1D 83 E4 57
 9B DE 48 19 60 7D 5B 78 69 E2 BA E2 6E E0 A9 9E
 76 D1 B0 29 B8 32 D8 D6 24 4B E7 ED FF B7 47 2E
 C1 3B 51 E0 B6 75 BD 23 61 F6 DE F1 DB 87 2E 6E
 61 E3 91 61 9A 7F 01 E5 48 28 9A BF 5E 71 CB F1
 DC DE B2 F6 F9 0A 3F E4 0F 21 3C BB 71 2B DD 5F
 50 40 0A 00 39 68 54 83 AD B0 C8 0B 9C CA E2 35
 E8 F9 54 A4 99 A9 D4 75 80 DF B5 13 B3 B6 59 EE
 38 B8 3B FA 8A 2D EA 0F 8E 56 EA A5 3B 24 01 FA
 6C B3 CC B8 0C 73 88 83 99 2B 5A 92 55 8C 69 69
 B2 C1 24 98 BB 50 E0 C1 FB AB 87 7B B6 BC B3 4E
 AF 93 8F 83 76 3E DF 0B 6A 77 97 B2 59 09 D6 B0
 D3 C4 11 B1 44 C3 14 A1 DC BD EE 2E A9 6A 5C 0D
 C9 32 55 29 66 C7 DC 9B A5 6B 7D 57 1D D3 E0 3F
 5C 17 52 A9 63 A3 D0 0A 3C 19 8E 05 B9 2E A5 7D
 5D 0C B2 B5 98 52 1A C5 84 04 D2 4A A3 D8 3F 39
 9F 6D DE 55 7C 3D BE 92 B4 63 68 ED 93 75 3E 3C
 11 C6 F8 72 75 26 2C 0D E8 A6 07 B7 4D 07 5C BA
 02 57 F3 C4 12 53 56 E4 EC 53 7B 67 F0 C6 EB 6C
 0A 09 C8 98 DD 77 02 93 4C 25 EA 73 0F F1 B7 D2
 B5 EC 58 A8 D8 42 7B 94 C9 EE 1E B7 86 70 0B 63
 F1 0F 56 B4 33 05 82 B6 C8 1B F4 BB 2E CD EC 66
 4E 2D 9F 36 49 F7 05 1D CC CC D4 35 3B BF D5 93
 CF AB C2 24 DC EC 06 9B 96 C5 80 15 76 9E 13 2E
 61 B8 EF C8 29 BE 04 39 2E 71 16 1C 97 50 16 2A
 E9 9C B2 0A 80 E0 B3 EB 15 3A EF 3A 6C 2B B3 45
 B5 48 12 2F F4 24 3E BB 96 88 DF E0 4A CB 9C D6
 60 62 32 F6 AE 3D FF B2 91 29 6E 16 2E E8 14 01
 9F F4 30 AD 57 5A E2 21 CB 62 D3 5B 89 F6 B4 2E
 5C F0 44 9E C1 40 C4 73 DC 93 B7 55 36 AA C6 D5
 7A 46 24 D2 8B 44 B4 6C 63 7E D0 DB 51 ED B2 92
 83 86 E3 06 0D 24 59 1E 59 80 91 DF 3C 7B 94 77
 7D CF 6B 99 7D 34 3B 8E F8 DD 0F EE 74 19 25 2D
 13 AD A1 48 0B FB 8B E8 74 86 44 7F C3 49 89 47
 0A F8 6B 83 97 FA AF 67 23 8C 10 BB B5 DB 1C 94
 50 38 1C E0 E1 79 2B 35 8A 5B F6 82 87 12 AD 75
 40 2A 22 D0 59 A9 58 6E 9F DE 3E DE EA 3D E0 36
 72 D0 53 16 A8 24 A3 3E 2E 0F 3F 17 3E 81 D9 88
 CA B8 C3 08 3A E6 AB A7 BD 64 37 80 AB 1F AF 59
 6B AC AA 11 93 8A 30 DC 9E 92 65 A9 F1 9B A6 42
 9F 4D F9 25 77 EB D4 E6 17 F8 8F 8A CD 6E AF 82
 1E 11 F2 AE D9 5F 67 01 F3 6E EB FD E1 A6 37 68
 93 55 0F A7 90 FE DA D5 5B E0 B2 F4 28 55 74 5C
 66 E0 96 8F 8A 0E 19 EB 1F 0F 98 CA 36 E2 54 F1
 1F 99 5D 0B 0C 28 5D 99 F1 3F C1 43 0C 85 B5 AA
 B5 B2 62 28 72 C7 07 A5 3C B6 A4 33 3B 2B 3D 00
 65 BE F5 AA 4B 09 33 81 0B AD D0 26 63 07 20 65
 08 A1 5C AD D4 EA 5E 60 AE 9F D9 FC 1D 53 37 0B
 2F 80 5E 0E 24 C1 10 7E AA 09 D3 2B 8A 73 98 70
 3E F6 4D 42 B0 FA 25 A2 85 88 80 B2 92 E7 C9 1E
 C1 9C 8C 16 EF BA 76 9F E3 B6 47 D6 AC E2 86 79
 A6 E5 2A DC D6 B1 C4 4C 58 77 A6 77 E2 38 84 E2
 7E 34 CB 99 43 EB 3E 0A 9C 19 C7 E0 32 DA CA D2
 90 E4 B9 A0 52 37 7D 07 7D 43 3A E0 15 BB A5 19
 89 46 B5 0C 49 A7 B1 A4 C2 76 60 E2 2B A9 F9 A3
 B3 B2 FE A7 90 93 DE A1 03 53 B8 FF 61 0A B3 7D
 39 F4 B6 2C 9C 0F 26 99 BE EA 19 59 A6 E6 E4 37
 46 C9 31 35 2F 5F A8 12 A0 40 C6 F2 BA BF 29 E7
 CA DD 6E 23 FE 05 5B 62 EC 16 4A 35 66 32 B4 17
 BF D6 1D 9D B2 63 0A A2 F1 D0 51 26 E3 AF 1B A3
 9D 43 D9 C4 3B 17 0C 24 12 61 70 D5 31 0E C1 54
 D7 0F BE 21 F9 1C 49 06 0D 0F B4 75 C8 05 40 F1
 A1 35 63 44 ED D8 81 96 5C B3 9E 88 34 44 1F BC
 E5 B1 10 9D 6F 63 0A A7 91 F1 B0 52 49 06 AC DC
 F9 9E A2 0A E9 4F 8E 8C 34 6B A7 1B FB 7B 0B 8D
 32 3A C1 49 0A EC 29 B1 4A 58 90 1E 9B D4 9E 00
 F5 43 7E 8C 9A 5E D2 F9 DA AC DA 29 09 37 F5 BE
 C8 6A 46 B5 FC AC 7D E8 0A E6 B8 7D 02 17 34 AB
 23 57 F7 06 94 81 EB E4 90 DE 2E 63 CF CC C1 8D
 1C 11 28 0C 55 D7 F7 D2 E8 03 23 A2 6E 7D 72 21
 3D 9F B8 CF A4 88 71 B8 41 E1 6D C0 FB 60 6A 07
 E6 09 C1 54 04 DC A0 18 79 BD 2E 17 80 6F DD 85
 B2 35 EE 8E A5 A6 60 3D C2 1E D1 F9 56 AA 4D C9
 AA 6C 15 71 2F 08 E2 2A A6 80 1B 6A 3F DD 8D FE
 83 4D 1B DC 59 4F 01 E3 32 8B 21 3A 5F 18 B6 08
 F6 F9 24 A1 8B EC 63 97 B5 EC C3 06 03 2E B8 1C
 3F 9C 7C CD C6 CA 06 D3 F0 0E F6 AD CA 22 AB 24
 88 12 0A 63 FA 60 8D CE C0 B4 96 D7 A3 80 7D F2
 B7 16 70 77 05 57 5E CE E7 5C DF B9 92 85 AB 12
 97 1E 22 2D B9 3E B0 32 65 04 9F E6 42 D5 81 C6
 6E D9 EC 8B 59 7D C4 25 06 50 10 34 12 0F 13 C2
 D8 CD C9 2A 65 B3 1B B4 6B 81 FF 1F 94 36 00 15
 73 09 F7 FF 98 CC 77 28 C7 BF 9C 68 36 6B CF EE
 48 5D 43 D2 27 77 73 39 0A 1C 0A 73 19 E6 B4 96
 F3 7D A1 FD 85 30 64 82 5C 9D 2E FE 0C 4F BC B2
 B1 4A 27 5A 76 09 A1 50 55 A4 EE 0F F0 8E 6A 6D
 4F 91 06 F4 75 ED 7E 69 D4 2C EB DD 70 0A E1 CA
 DD 7F 19 77 BB A7 2E CC 68 75 1C E2 60 42 CB 54
 C6 98 B2 66 25 CA 2B A1 A0 19 BE D8 F0 66 BD 74
 B9 91 DB 3D 00 CE 49 F2 A9 8E D2 23 C7 A3 3D 89
 F4 A0 10 50 B7 A0 2D EA D3 3E 0E 7D 2C CA BB A8
 9D 4A 0E 72 11 35 3E A4 70 F5 E3 76 BF 67 DE 2A
 93 C1 41 64 A4 29 77 BA 11 A7 35 2F 7F DB 00 73
 6A B1 EF 9B E5 C6 B1 05 47 A1 91 29 FE 82 01 7F
 BB 10 E0 C0 6F 2F E6 4E 8C 04 47 7F 9D 92 61 19
 0A 93 5C 6D 46 3E AE 46 2B 84 D3 BD 83 44 84 73
 AF 30 44 A9 FA 71 40 2A B3 3E 63 F7 0F C4 C4 42
 DE 29 1D 1A BE 44 C8 12 78 E3 AF BC 25 66 8C 14
 63 5F 00 69 6B 14 FA FA A0 63 77 4F F3 00 F1 B2
 18 84 13 AF 79 05 4E F9 4A F4 8E 74 F7 6E CA 6D
 7B 0D 4E 3D 51 9A 45 B0 1F D9 4E DF 06 DC 32 F8
 08 9D 2D EB 8E A2 65 95 9B DA 31 3D 60 FA C3 85
 60 99 DB D1 DE D3 02 DA D0 DF CA 89 06 31 97 0E
 B4 9E 90 9F DB FC AE 61 93 DA D7 AF 68 58 C0 1A
 FE D9 8F 27 88 4F 32 C0 9C BB 0B 6D 43 89 94 5E
 40 D5 27 DD 23 CE C4 78 16 FE EC DD 8A 20 69 87
 A1 D9 A5 10 85 C3 F3 8E AB 20 7F 1A 8D E0 A8 26
 2B 90 C0 C2 AB 3C 7C BA A5 E2 F9 92 74 68 39 0C
 C5 F0 6F F6 04 CE 98 F9 6F D2 EB D7 04 4D 54 CA
 20 A3 75 5A 4F 57 54 B3 06 A2 00 4D 7A 43 73 26
 10 11 49 19 41 92 D7 63 07 37 61 AD AF AA 3C 5A
 6F 5A 8A CC E9 7C 7F 43 6A F4 52 B6 95 C3 52 84
 2A 40 2C 63 8A 63 1B 89 75 1C 7A 55 A6 A0 57 51
 2D F9 77 4D 6F E4 84 F3 7D AB 4D 37 F4 12 92 ED
 49 42 A4 BD 22 4E B2 46 A7 9F 08 8F B5 49 17 3B
 EC 09 F2 F1 9F 66 EF 14 09 98 E2 C5 95 F3 5B 77
 EE 20 D8 2B 6D 4F A3 75 86 52 26 3A 0E 82 DA 4C
 0A 9C 1A BF 43 E2 57 A0 47 70 F1 86 9A EE BB 15
 85 52 F0 60 43 F1 BE 6E 71 CA 71 E7 35 BA 2C 9B
 D8 9C F9 75 D8 6D DC 40 15 C3 42 39 74 A1 1C 68
 23 06 8E 89 AA 4B 2C E5 97 6D 62 63 69 57 9F 0E
 BA AD EE 50 58 78 B9 74 0D 46 17 7C C9 43 AB 40
 FB FE 76 95 31 85 DB 4F 0D 3A 8B 54 13 9C F3 15
 1F 6E 33 71 16 01 6D 4F 95 88 3F 67 56 31 C2 86
 1E C6 1A 3F DA 60 F7 37 E3 14 45 27 05 DE FA CB
 D6 06 FB 4A C9 38 0F F1 A4 4B 90 E2 C7 B2 FD 21
 34 F8 36 41 C6 D1 01 98 32 B2 FB AD 58 13 7A 2F
 CA B2 7A CB B8 36 96 4A 68 6B A9 C1 64 9E 73 D7
 7B F9 73 DD DF 88 CF 31 50 33 13 81 30 51 CC 4A
 8D EB 03 2F 69 08 B2 AD 26 AD 7A BB FF 9A 16 02
 EF D3 EA 12 16 4C 27 C8 E1 43 D8 18 5C 6D DE BA
 36 31 E4 64 AF AD 73 F5 88 C0 94 A9 1F 74 6E F9
 7D 4C 77 29 BD 1C A5 DC C5 84 80 82 07 78 DA 18
 02 F8 B0 6F 21 35 6F 37 46 B0 80 07 1E AC 1D 62
 5E A5 C9 50 0E F9 06 5B 90 06 F8 09 80 73 A3 49
 37 86 ED 43 9D 4D 77 0E 4D 49 1B D7 68 D1 68 8F
 5E FF 00 57 C6 21 02 32 18 B2 EC C2 7A CD EF 11
 2B 6F 7E 47 D5 CB 94 BF 3B 5F 7E B1 56 C8 31 35
 59 71 0A 8F 74 CE FC 8A 4A 78 C1 23 CF E2 98 CB
 FC A4 F3 A4 00 59 97 79 68 96 22 45 FE 8D 42 01
 72 FC D9 85 70 05 28 FE 04 A3 63 A5 15 5E 35 74
 CB 92 91 2C 84 04 07 77 CD EF F4 24 27 17 E0 DE
 B3 B4 4D 55 4A FB FB 15 8E B4 D4 18 B2 C4 CB 88
 CD B8 81 64 15 DD 44 6C C9 9B C8 B1 A6 0F 00 E5
 BD A4 A3 64 0C FC 9D B9 85 E0 7F D5 05 B9 C0 F6
 DA 58 E9 6C 48 1A 63 A5 9E 43 4D 38 21 97 13 AD
 6E 15 12 9B 39 50 F3 2D AC 40 83 4A 97 3E 88 AA
 A8 BA B6 44 84 E8 11 8F 3F EB 70 27 D9 02 CC 33
 A1 23 47 F9 3D CC 8E F2 45 90 69 AE 53 71 DA DB
 EC 72 B0 32 72 F3 9D 4A 1F E6 F2 88 13 81 ED A5
 37 A5 98 86 FE C1 C9 C5 4E 6A 18 F9 5C A2 60 60
 DF 25 05 72 DA 56 C6 B3 97 F5 92 F3 94 4E 38 DE
 CC 1B DA 21 FD 25 9F 93 39 62 E5 30 0C 34 8E FD
 DF 8A 90 21 C5 D5 29 33 F3 04 B0 4F FD 48 88 24
 E3 18 B2 F5 94 FB 6F E9 A0 7E 56 75 86 2F 4F EB
 2D 33 C4 9D 21 6B 9E 2E CF F8 7A 8A 6C 0C DB CC
 DD DE 40 F5 64 B3 1A 6D FD 43 18 BF E1 FF 83 E2
 1C 0A 0D 17 1F 8A BD 81 3C C7 4C A6 99 4B D2 32
 0A 37 1E 09 94 42 13 33 4D D2 82 45 F1 45 D3 F2
 98 52 75 F3 EA AB 14 35 5E 42 78 3E 51 29 09 8D
 0C 13 AD A4 F1 29 CF B8 3D 21 C1 63 0A C7 AD 24
 39 4E 31 BF 47 84 3B 46 22 F7 10 7D 66 B5 1C BA
 7A 9D 59 EB 42 AB F4 12 18 76 AF 65 1A 33 FC B6
 CC 17 22 16 1E ED 40 1A 10 B6 40 B1 A0 B1 17 3F
 1C BD 98 70 42 BC AF CD C3 A2 7B 2B F5 F2 9E A4
 B1 55 B9 36 E0 5A 68 31 A6 10 B0 E4 96 10 9D 74
 59 B9 81 4D 47 6C 77 61 94 E5 FE 65 8D 71 16 32
 44 71 9E 00 BE 5D 72 16 FD D0 B2 CE F4 6F D5 26
 E5 A6 C6 56 D7 DE 51 63 1F 0F F1 8D C6 B5 35 16
 72 B9 AF 14 09 63 E5 80 B0 58 6B 0A D6 E7 5D EB
 C3 D0 A6 50 D6 06 6A 7F C3 A7 2F AF D0 5E 40 39
 E0 46 30 B3 96 76 4F 31 FF B0 03 3B 54 9E C3 9F
 B5 1F A5 A7 49 E8 9D 3F 58 1C 71 A4 E0 A0 5F CF
 72 51 3A 09 96 49 B8 DE D2 8D 8B 21 34 41 7F 82
 CA 41 06 6E 63 3F F9 9D 53 3B 00 D0 A7 1B EB 84
 DD 7E FF 31 37 22 2C A0 2C A3 56 AA FD 2D 81 79
 BC 69 E1 B8 F3 04 76 82 4F C8 AD F0 1E 4F 8F DD
 43 94 A2 05 6C FF 78 2F 28 74 D1 C7 86 B8 43 45
 0F 6E 2D E9 1D 5F 7B 06 12 FC 4C 50 B8 67 85 C2
 5E CE DD 08 FF 83 80 D2 DE 67 06 DB 6C 7F 73 E1
 63 C7 E3 81 6A 38 55 05 F3 FC 27 BD C4 80 F6 55
 BA 47 87 93 0A 71 74 B8 08 4E 61 8E 66 97 11 09
 3D 65 FE 6F 67 43 C0 DE 04 AE FE 9C 65 A4 71 ED
 05 8F 59 F2 84 F5 4D 78 82 31 25 52 C7 1E 32 75
 34 26 6A B8 5E C3 D5 10 C6 64 DC B1 6C 61 88 0B
 D8 FF 63 3B BC 38 CB F0 6A 40 E2 03 2E 35 B9 53
 46 D5 B2 56 C5 7B D7 D2 2B FD 6A C4 D5 BA 3D 37
 21 22 DE 26 94 3D C1 8A 64 13 8D 6C 90 0A 31 56
 44 52 0C F3 2F 63 F2 87 D0 02 49 9D F5 F0 B5 26
 A1 97 4B 76 A4 3F 91 F1 F1 70 FE CD 4B 16 8A 29
 C8 01 DD FF B5 AA 30 10 49 0A E7 CB F4 B1 DB 1D
 6C AB 27 7A 15 39 32 4B 7F B1 7E 19 6F FF 0A 2C
 E5 96 BE 28 63 A2 C9 11 3D 1B 9F 01 61 22 07 44
 4F 4B DB F3 FD 1F 2F EF BB AA 08 E8 2B F1 DB FE
 1B 9A 73 F3 DC 03 6B 3F 63 51 28 21 E2 C8 C8 0D
 9F 13 CB 92 39 C1 55 30 61 27 5C 13 5B 24 C4 38
 32 0C AF EB 40 51 69 3F B6 89 42 2F C9 88 2C 8B
 B6 3C 19 27 7B 0C 4C D7 2A 78 50 A6 34 58 84 75
 AC 31 56 74 F7 95 6A EB 03 C7 61 3D 03 E6 8F E8
 C8 92 88 DC 51 78 12 04 9D 60 9A 77 5E 4D D9 29
 67 6C 80 2C 98 45 28 DC E1 A8 51 7F 8A B4 96 0F
 CF CD 60 F2 6A B7 72 41 C2 95 88 78 BB F1 23 83
 24 4D CB B6 E3 E8 73 5F 52 9B BA 72 6A B8 2C 5A
 77 3A 82 15 53 4E E0 01 66 EC 36 FE 74 36 96 7D
 AC 1F 26 8D D3 67 F7 A0 62 6D 56 EE 12 56 A0 9A
 8C 2D 1B AA 2D 2E F9 E5 AA BE 1B 0B ED EB DD EB
 05 E2 11 DE C4 7E D6 B5 CC F1 4F 7D AF 2F D1 C3
 8F A9 BE A1 C2 C7 63 91 F3 C4 EF 6E 42 78 3F 0D
 BA 34 84 38 FC 25 F7 8D 25 66 AF 67 9D BB 1E A7
 8B 0F 58 9D 96 A1 74 88 7B 88 A5 AE 21 40 DC F1
 4F 16 C0 13 DA FF 4B 8E C4 3D F5 D0 77 5D 4D C4
 3F A7 46 37 F5 CC 0D 94 C5 97 A1 E6 E2 84 AB 21
 29 1E 3B 8A 8B 75 EC EB A7 68 4A 05 38 A2 7E 70
 A1 A0 5B 97 8C DA 14 A2 72 AF C8 52 20 D2 72 05
 0C AE A5 E1 74 18 BC 09 B9 3E 18 BC A2 92 0D 8B
 E4 44 35 4D 74 40 0D D9 A8 5C 96 CD E3 B4 8B C9
 94 06 7E D1 F8 E3 00 35 DB BE 57 51 5F CA EA B8
 46 C1 75 09 AD C1 D3 1A 73 F2 31 05 26 39 4F B7
 E9 BD 2F 65 57 70 A1 CD 31 F9 8D 0F 7F AF 48 9B
 6E 3E C4 CE A2 C1 73 CE 70 B0 D1 AC 92 9A AC 5E
 CE 92 B9 9C B5 51 7A 30 3E 2B BD 39 F4 27 EE 8E
 62 84 2F AE 08 93 EA 87 70 D9 9C D2 12 0A 42 AC
 50 7B 3A C5 8C C2 1F 6C 37 95 E2 65 EC D3 7A 23
 F3 BE E1 BA FA 4C A6 9C C3 77 F5 43 3B 09 F9 00
 C5 36 AD 25 51 4F BB F0 5B A4 CF 7C 0C 76 F0 07
 A2 BB 98 F1 92 68 78 7E 40 62 6B F9 14 FF DF CC
 2C E3 2F 29 C2 64 ED 9D 6E 67 B5 5E B4 2F 15 A4
 FF F5 F4 40 67 B8 BC AE 5A 53 2B E1 8E 14 8A 82
 58 9C 2F 3B B5 87 CC 3C 67 37 8A CA 88 B0 E9 58
 9C 1D 81 A2 51 00 4C 15 34 11 E1 57 DE 0A 36 4F
 9D E0 21 58 61 66 36 5C A7 23 0C 78 2A 60 74 1B
 F8 44 F4 75 1B 7C AD C6 11 F5 5B BD B4 C8 A7 2B
 A8 45 C6 62 BF 74 31 0D 43 B0 AB 52 E6 F8 3D 71
 4E CC C3 B9 05 67 F5 5E E8 2F DF 7B 47 EF F0 21
 DE E3 32 32 A2 D1 DA E3 51 C6 A1 ED 2E 5A E0 B5
 50 A9 AD E2 25 B5 51 6D 25 66 1D 60 03 83 60 30
 FD C4 ED 0F 67 5F 21 1D A7 62 FC 63 BD 31 91 11
 D5 56 3F 25 71 44 62 B1 29 8C F4 44 39 69 D4 2B
 40 97 E2 2B 4D E9 99 D6 A9 BD 57 A2 7B 5A C6 A0
 9B F6 B5 EA 3C 3F B3 EF 1F A2 3B E4 EE 91 3B FC
 7A 82 74 26 20 D8 01 EC 23 53 0B 1B 1A E4 D0 A9
 E0 55 EC AE 7A 3D 53 70 00 92 76 59 8B 32 86 0C
 8F EB AC BC 41 EE 60 F6 A8 D0 39 B9 F9 66 87 31
 76 FA 07 80 FE 16 47 85 72 DC C1 42 01 69 E2 81
 D8 D0 A3 91 4D 36 AE D2 31 F4 51 9B B1 B5 3B DA
 21 D1 56 72 3D 2C A5 92 98 C4 6E 76 BA 81 4B 4E
 ED 4E F9 77 6C 79 9F 9B 47 79 1B 2B 92 46 12 EB
 2D 3F 5A 4A D9 63 54 15 9A 25 9E 33 80 70 4E 66
 70 B2 75 88 A0 65 33 57 2A 4F 59 E9 62 F7 28 50
 04 71 C4 9C C0 23 BC 69 10 16 70 99 65 42 47 39
 42 05 1F C3 2A 7C 9E 32 83 68 4D 27 25 1B 67 DB
 34 29 5C A1 D1 39 D4 BE 11 29 75 93 0B CE 5C AC
 B2 5B 2E 73 A9 13 53 81 C7 04 59 8B 09 23 87 43
 7F 4F 64 34 08 9C 12 1A 8C 96 A8 A9 07 52 B6 CD
 DC 80 91 09 D2 76 72 5E CE A8 91 4D 86 DF E3 0D
 E5 98 84 58 2B 85 DC AD F9 F9 BD 82 85 A9 2B AB
 01 7D 5F B7 8A 4F 1B 77 79 3D D4 31 0A 0C DF 86
 C8 2E B5 EF 0C BB F2 E8 4D ED 93 D6 F9 1B F6 94
 23 90 78 C0 41 DE 6C 0A 86 9A CA 58 8C 59 04 29
 4D 2C B3 4E 02 31 B5 17 91 8C F8 C7 62 90 EF 66
 64 1D 28 A5 E2 09 5C 47 5E 70 9E 93 79 4C FD C6
 47 A4 DC 63 0C 98 69 A7 4F A2 A6 C6 1E DD 0D B5
 75 68 BA F7 4B 92 35 54 92 14 70 D5 82 DA 1D B0
 04 6A D4 84 3D B7 02 10 CF 18 E6 84 E0 BD C0 2E
 56 AB 4B B8 5E 44 78 74 09 A1 AD 92 3D 0A B6 93
 39 1E 9B 98 23 7A B0 17 BA C2 C7 2E 4F C3 5A 2D
 C2 8D C2 C4 FB B6 95 62 4E 84 96 F9 12 31 58 B0
 42 1E 91 09 EA C1 C1 EA 2F 93 2A 32 50 7B 29 9C
 79 2A 39 8B DD 18 6A 65 B0 80 AB 68 F6 9F 92 70
 AD 4F 45 4F 9F 4F 0D 76 2F AB 90 54 F2 B3 EF 26
 FF 2C 7E 3D 3C 37 98 72 E1 64 D0 27 27 D8 55 2A
 6A 86 48 D2 4F 8A 94 A3 65 77 F9 63 14 03 3B 73
 E2 84 67 FC F2 BE 99 BB 35 7E 52 74 A4 16 D5 8A
 B4 8B D4 2A 94 D4 48 02 C7 6A 19 9A AB 15 E5 D5
 AE 86 19 D8 2F 94 58 95 1C 19 7D F7 25 7B 72 1F
 C8 1A 2B 02 B5 20 66 97 62 2B A3 11 0C BB 44 46
 A9 BE 09 3F 29 76 EC A8 62 70 9E 61 6F E2 F9 87
 96 C4 39 9D AE 38 4E 9B B4 3D C0 31 A5 5A A9 5B
 2F E1 0D 05 F8 8A 98 1A 07 69 1B 0A CD 3E 9E C8
 26 31 26 26 54 BA C3 4C 48 B9 84 3F D9 EA BB 8A
 F8 EB 33 B4 9E 27 EC 05 00 0E A6 01 9C 13 67 DC
 C2 5F B5 E2 19 E5 49 45 F5 16 28 D5 91 61 86 2C
 C4 1B 33 92 45 D9 E3 A7 63 8B 15 48 CF 33 FB D2
 21 1C 7C 76 01 C9 BA 9F 84 8F C9 A8 F4 CF 46 DD
 CD 20 24 E5 AF 2D C6 C3 D8 F3 8A AA 18 1B 76 16
 78 DF 1D FC E6 48 98 09 EA A7 0A 28 53 08 75 73
 BE 1C 83 02 FC 34 EB BC 1E 31 11 91 19 BB 0C 7F
 6B 79 E2 AF B4 87 13 66 D5 3A DE 1A E3 51 C6 AF
 3A 65 E6 62 CF 73 8C EE 59 D5 C4 A4 E3 6A 49 1A
 71 03 F9 D7 04 40 68 35 C4 73 AB AE 0F 89 44 09
 B6 62 A5 C5 8B 55 06 46 C1 7B C5 CC AC E0 EE CF
 89 2D 61 67 C6 19 49 2A 41 02 8A E2 81 E4 40 52
 7D 62 52 C8 FE 93 3B 39 76 A0 E9 F0 27 98 B8 2A
 45 67 30 B2 E9 F6 4A AF BA B9 E2 CA 60 45 68 A7
 B7 55 6B 50 AB C4 D5 13 F7 2E 80 6D B0 21 EF E4
 93 42 E5 C9 4C E6 F7 17 EE E4 ED 45 69 67 91 9C
 40 D0 15 D0 34 BC 23 7C 1A 61 5D 9E 24 4C 4F EF
 06 3C 29 36 14 7B CA 9E 24 15 97 4F E7 C0 60 95
 46 EC FE AF 80 A7 AB 60 A3 35 97 07 16 60 28 2F
 46 2B F3 14 30 02 D4 3B 57 27 48 7C 02 3C 9F A0
 B2 88 67 8A 12 F6 8D 5D 88 C4 1E 91 34 7A 86 6B
 82 4A B4 5F AB BB C0 97 D2 C9 F7 DA 11 AE 4C DF
 54 C4 68 E1 EF 7F 88 16 C5 2B 9A 35 39 F8 44 05
 92 01 02 7A C5 EB 72 FE 46 9F 1B DF 71 07 01 D7
 94 88 DA CD CE 26 FC FE A1 D3 7F 9A 65 C8 86 F9
 7B 37 45 F9 8A 05 8C F8 83 D1 06 DD 3C C4 13 18
 F3 59 A5 63 A4 54 81 23 1D 6F 23 82 82 4F 45 1E
 DE AF E0 D3 B7 63 71 21 C3 6C 6C ED F7 CA 39 FA
 55 B8 97 B6 95 51 6C 74 48 35 B3 02 36 E9 18 1F
 2F B6 50 5D F8 FB 4C B1 FD 4C 28 03 EC F7 63 80
 08 04 76 B6 F7 48 20 17 45 38 93 5A E3 62 EA 05
 76 09 F0 D6 55 33 D5 F4 83 C9 40 31 4C 2E 67 B7
 D0 34 B2 69 F9 7A 35 5D 65 DC 35 6E 82 93 C3 30
 0C F4 64 5F 74 98 A8 C4 A3 40 79 5B 6D 3F A2 11
 BB D5 DA 7B 8D 34 19 5E AC 53 49 75 BB DC AD FB
 CB F4 D2 26 82 B3 F5 79 F5 87 86 01 0B 2C 07 DF
 89 98 BC 27 3A D0 8D 84 6D 20 BE 2F 6E EC 46 D3
 7B 40 FE 06 85 97 B4 DE 85 39 95 8D EF 40 19 2D
 01 B5 DA 2D A3 90 55 90 2F 38 48 B2 DC 38 EA 53
 44 C9 DC A8 0B 7C 68 DA 31 59 AA 5D DF 08 79 48
 5C 1C CF 17 4E 1A 46 71 3A E6 6E 77 05 E4 0C FA
 9A 6D 5E 98 3D DC 1B DD 49 D3 A5 36 2C 00 A4 6A
 A2 57 E2 22 DC 17 E2 14 77 35 A7 FF 2E DD 73 DB
 57 A0 2E 58 14 AB 2F 48 46 86 CA E9 8C 9D 90 A0
 45 55 C7 03 8E 8F 94 52 1F 13 95 33 2C E0 AE FD
 23 81 2C 79 AF 40 9C 95 68 69 60 C1 FA 30 00 33
 D8 26 F7 BF 75 16 F6 08 11 16 48 61 6C 38 BA A5
 EB 9C 88 85 1F 3A CE 20 E9 9E F0 E2 B3 07 F8 11
 14 FC 8C F9 F4 4C DD BD 59 F5 44 30 51 D4 35 31
 9F FA 95 9F 99 35 B3 A1 20 53 5A AE 37 F3 E8 D4
 05 66 A1 D9 51 EF 63 FB 21 08 5B 56 5C 9D 82 A3
 28 B4 10 62 18 F2 A5 C5 1E 75 19 5C D3 BA 85 1E
 E9 12 FD 5F AF 1B 58 FF 1F 17 A4 05 69 2D F5 1D
 D9 8D F7 24 87 4D F7 C1 EC 90 1D B5 D8 5B 4C A6
 9D 53 E8 32 EF 5A CD 5D F6 BF E3 10 99 55 70 9A
 4C F5 0E D0 B8 98 88 2E F9 09 9F BC 9D 5C 3A 88
 35 FF 0D FC D6 CD 36 5B 94 D2 67 DC 39 24 E6 A7
 3C 96 5F 49 7A A6 61 48 34 17 F5 78 F7 EE C7 82
 48 5F B2 3D DE 20 16 91 99 F4 2B 2D E5 A3 4B D4
 10 12 1B BE B6 56 F8 EA 73 24 B7 D8 1D 91 2E F1
 E3 20 ED 44 6E 1A 52 D0 A7 6E 23 A6 BB DA 5B A0
 04 5E C7 44 B2 AB A0 F6 06 07 7D 67 E1 15 68 0D
 63 25 66 CF 58 F9 AA CD 0C 0A 56 2A 85 59 E0 D3
 A7 26 06 AB 39 55 A9 D8 5A 69 04 EE 73 F7 7B 4D
 C7 49 71 F8 00 C0 54 B1 D0 DB E8 8B F6 5D 57 9E
 6B 5A 28 09 90 7E 81 73 8E 73 28 CD 87 21 0B 2D
 5E BE E9 38 76 A1 5C F1 50 DB 55 EA 2D 19 10 04
 D7 45 2E 60 87 27 47 2B E8 76 BB A6 34 4E DE D4
 AF 2D 70 48 5D BB CC AC A5 BE 36 CE E6 77 0C 26
 57 23 FF A3 5C 7A 94 AC FA 9D 8B BF C9 94 A6 79
 02 C2 51 1C A2 C1 57 0D 55 58 18 3D 8E F6 40 54
 0B 7A 46 20 CC 20 BB 66 A9 C9 1D C8 1D 3B 5E BA
 26 E3 D2 AE A8 5C 30 8A 31 CE E5 A2 AD 3E 75 2B
 31 F6 D8 0F 2A 37 C1 F2 F5 1D 57 85 B5 B4 9D F2
 80 94 0F 76 F4 86 D0 48 40 F9 26 A6 4B A3 80 BB
 28 FC B3 A2 76 9A 6D 4D 7C 07 D1 65 71 D8 6F AD
 88 C2 74 1C 16 E3 D3 1C 13 CB 17 39 3B 99 BA E0
 36 C8 58 75 F4 E8 0D 95 30 D1 49 95 66 0C F1 6C
 DF 30 4D 0A FE 57 FB 5D 10 A2 EF 27 43 64 8A B1
 59 84 9C 1A 40 C5 0B D7 AE 2C 54 88 D1 AE 96 39
 AD CB 91 50 03 77 D1 E2 8C 15 C4 EF 49 2C FC C2
 9F 13 13 78 C2 BB AE 9E 9D E1 9B D1 BB 3B AB E6
 B5 CE 80 BE 6A 75 2A 3F 23 E1 BA 89 B6 7C A6 74
 EB 32 5B BB D0 90 2A 67 9D 6F 1B 5C 84 82 36 C0
 5A 27 41 A4 D5 47 85 D7 2A FD 05 83 3F 72 4C BB
 26 45 07 F5 DC 55 58 51 CE 0F 03 3D 48 16 B3 6B
 F6 B1 6E 01 63 14 00 E3 EB 13 28 BF F1 23 96 0D
 E0 6B 62 FC B4 A5 2D A2 19 C1 05 67 21 C0 5A 71
 21 7B 29 59 E8 A4 DE 63 84 59 31 B8 EB CB 9C 7A
 84 63 B3 77 8A 90 9C 87 97 9A C9 2C C6 2B 1D 6A
 6D 0B 51 88 71 D1 D3 AB 81 FE 7A 78 F9 07 5B 70
 5C 03 5A DA 2C C8 0B 89 35 0D 93 70 47 F7 13 69
 16 2A 21 9D 0D 4C A7 2A 5A 82 1F FB 18 75 F1 1E
 02 6A 1F 17 4E 62 43 21 BF 51 94 B0 85 1C BB 24
 70 96 F3 1F 78 42 AC F1 A7 D0 EE 09 85 77 59 90
 DB EA 99 E2 C3 6B 6D 36 54 7E 40 34 AD D8 D8 B4
 4F C7 62 D8 DF CC B1 45 01 A4 54 B1 62 E9 88 37
 C8 1E 4F F4 55 DF 3C E1 39 27 B9 EC 57 82 1C 87
 98 1C E0 03 C2 EF 8F 82 2F 8C 1F B9 3F 86 58 6D
 4B 4A CA 03 71 68 28 C4 CE 60 90 07 0A 43 5C 6B
 BC D9 28 19 3D A8 DB 10 25 FB A3 D8 BE 54 D5 58
 0A 3D F2 3C 2F 70 30 F7 61 AB 91 EF AE E9 A2 72
 AC D5 AA AF EA 16 90 54 C6 F8 87 2D DE 24 1B E3
 F8 E1 22 C6 BF 3C 2F 85 45 9F 3F 00 27 BE 84 9C
 F2 F3 C2 6E 70 B8 E8 64 24 AB 7F 24 43 9C 78 63
 3E 53 04 30 15 60 3B 46 95 8E 39 F2 61 46 DB F6
 AC 57 6E 9A 5D C2 77 48 AE E1 87 4C ED 09 E1 04
 8A D2 50 77 DA EC B4 C5 84 AA 18 EA 45 EA D1 84
 57 73 C0 EB E1 3E 56 00 45 CB DE CB 4F AF 80 17
 F7 09 2E E5 D7 1E AE 55 58 42 37 77 88 75 3B 90
 8D 59 46 CF 5B E4 97 A4 8E 09 0D 40 CC 4F F2 51
 E2 13 CA 41 09 A1 EB 5B C5 DB A0 DB 23 1B 78 64
 BB 24 53 90 A7 34 CF 79 F9 DD D3 37 E6 8D C9 14
 46 D7 4A 6C DC 14 52 AD D7 62 AB EF D6 A3 38 52
 5A C4 01 E6 11 55 59 BE E5 B5 45 BF A6 30 74 44
 09 FE 8F 92 91 FF AA 0C 48 EB C9 7F 65 7F 2C 44
 03 7C AA 39 A9 B3 DB F9 7A BD F8 12 E4 03 23 65
 3D 1F 68 F2 9D EE 83 E8 81 E9 31 E3 39 56 B8 64
 6E B8 F4 C1 62 39 F6 C6 AB 5D 7D 18 F4 9C 3D C8
 37 6B 95 C0 C1 1F B6 3A EC 74 4A 29 B7 86 FB 6D
 96 90 4C D3 97 F7 68 32 C5 B5 00 1F 3B 45 AA 30
 26 E9 99 3D 9D 67 3D 1E 32 00 99 53 EE 25 7F 2B
 EE 9E 1B 82 42 4C E4 85 C9 06 F6 BE CF 51 56 A8
 58 93 09 EF F3 1C FC 6F 31 A4 78 3A A7 E2 12 E1
 D0 C6 53 AA 73 6A C3 80 C2 5B 7D A3 24 5E 94 00
 2B 2B BF BC 56 63 04 C9 FF EE A0 82 F9 02 FD E8
 42 23 85 5F 03 85 05 FF 3B 4A B2 A8 4B 57 F7 29
 CD 9D EB E5 23 6E D5 E2 71 FE B6 10 E1 50 24 15
 0B 0D D9 EB 33 A9 12 D1 EE 63 AB 9E FA 1C 49 77
 20 25 C1 71 FA 2D 26 73 30 90 66 A3 D5 80 AD A8
 CD 69 FA 49 30 2C F2 48 4B F3 EB 23 1B 75 C7 CC
 6A AD 18 7E 5E 49 7A 70 98 5C EB 1F D9 DA D4 5C
 28 C3 2E B4 2E 86 25 4B 76 03 4C 15 EC 5D CF AD
 3F 48 F4 77 A6 B1 95 85 87 E0 E5 0C 98 DA 15 BE
 EF 18 09 CD 4C E6 32 45 FA 97 22 24 F5 9A A2 F5
 D3 56 BA C1 35 75 A7 B7 11 B0 E0 42 9F F1 33 BF
 95 72 98 A2 B8 E1 2D C9 2D 41 F7 84 60 D1 BB AE
 D8 92 09 E9 07 F7 48 48 40 D3 09 CA 12 3A 37 83
 59 D0 00 48 51 E8 84 BD 4C DF 71 05 B9 DD 37 66
 FC CD B6 3F 65 C0 2B 82 86 E4 4A A1 35 9A 7F EE
 72 BE BE 07 E8 A4 50 D8 7D B3 99 B5 FD 3B C4 DD
 42 C0 94 A9 35 CF F9 AC D4 92 C5 C8 30 D4 72 99
 DD 94 2B 86 61 3A E1 4D 4F C2 C5 AB 34 67 6A 70
 86 EC C9 F8 C3 F7 02 E1 EC 00 56 5B 55 04 8D E0
 C5 57 31 13 78 7A D1 04 2F F4 8B 5B 74 7F D6 8F
 03 4A 6B 2E 53 68 76 C3 14 8D CE 27 C1 8B 07 BF
 04 9E 4B CB E5 92 F3 7F 69 CA F8 90 98 05 40 44
 E5 D5 93 C6 14 22 A0 08 1A 23 08 0C 01 A3 F7 D1
 25 59 1F 03 06 20 E7 49 0D 05 92 ED 36 9E 23 B9
 90 4E D6 16 EE FD 7C A3 69 19 97 44 24 12 EB 41
 A8 A1 25 40 08 3D ED D7 F4 04 92 02 0A F9 DD 0E
 0C 82 47 BD 4D 3E 16 55 97 F8 A7 2E 7F 03 3C 03
 49 D8 1A A1 D7 EC 78 99 02 4C D7 33 E6 ED CD 98
 FC 43 89 A2 19 D7 49 95 1E AE 96 C7 F4 44 8F E3
 A4 DA 0F B2 A4 E7 E0 55 FC 26 8C 1C AC 67 6F B4
 24 82 6E 27 24 41 AF 1C 64 A6 0D BF 48 BE 4A 1F
 A5 1A 52 D8 64 80 B3 BF 6E B9 64 F3 A5 9F 3C 4A
 24 E1 06 CD 60 EA CB 53 8F 15 F8 FD 2C 92 0B FB
 D3 2E DD 21 39 DC 68 F0 71 6D 51 0E 84 57 47 E8
 A0 08 28 7C BF 90 26 E3 31 36 4F 6E 70 F7 CB 7D
 EE B7 40 BD 0F 01 B0 06 21 D0 27 4A 3D 87 94 FA
 12 61 CE 8B 87 40 41 13 75 9F C6 3D F6 B9 05 C6
 47 A5 5A D5 41 09 85 47 3B 74 D4 34 57 26 C5 37
 25 F9 B6 49 1B C6 82 4C A9 9E 15 E4 79 C0 C2 05
 16 D2 50 F0 B5 7C 75 B0 81 B7 97 8F 9B FE 45 86
 88 15 46 AC 42 0A 66 6C 59 14 AB 9F 31 83 24 30
 1A 0D B0 C1 E1 83 4A 48 70 0B 51 FD FB 18 86 9C
 9A 97 EA 8E AA 11 65 5E 5B 6A 99 B1 9D 53 C1 20
 FD 38 71 9E D7 61 16 8E 1E 99 67 22 DF 7D D6 3C
 4A 4A 12 0D 28 43 89 01 55 9C 8E 3B B2 EA 23 89
 3D E6 56 05 3D E0 45 20 C3 D3 11 1C B1 BE 93 62
 98 BA AA 4E F7 EF 47 A7 F1 D3 E4 3D 6D 23 B4 0B
 10 DE 7D A5 F3 40 8B D3 47 42 0F 12 2E B4 C1 F8
 5E F8 7C 17 2A 81 0A 65 01 B5 9A DC 40 8D 28 4B
 B2 03 43 70 9C 59 20 7D 00 EA D3 F6 87 B2 A3 51
 8C 6B 05 B3 9D 23 5B 60 B1 BD BD C3 40 64 B9 89
 0E 0A 64 A6 2C 16 7E AA 40 DF B7 47 FB 8B 5A CD
 8B B0 3C F8 4C 1F 79 F7 C9 3D C4 E8 17 62 2F 57
 2E 3B 08 D6 40 6E 5B 20 98 70 74 75 94 16 73 6C
 D8 72 2A C2 94 FE C2 DE 6A 00 93 41 A8 A7 25 01
 D7 C0 BE CA 80 DB B8 6A 7F 1E F4 C2 1D BF 20 BB
 0A A5 E0 CA F4 98 11 26 11 3A 45 48 F7 07 FC 12
 5B 45 96 2C B7 72 49 60 1F 1E DD DF BC F1 5D E7
 5D A7 6E CE 36 D0 E0 BB 07 96 52 06 8A 7C 74 24
 6E 26 BC 2D EC BA B2 4C C5 1A A4 01 A5 3B 60 EB
 1E 2A 11 24 1E 3D 79 ED 26 AF 0D A9 80 71 C9 1E
 D8 72 AF 45 42 96 83 57 18 32 52 BA 71 A8 2E 4B
 66 92 59 F5 C7 D6 4B A2 C1 C8 5C BB 41 1A F9 03
 47 03 31 B7 C8 43 E3 B2 E6 DE 46 91 CD 69 FD 3E
 16 83 CD 40 42 CE 0D 0F 67 75 92 B6 62 02 5B 93
 FF F8 9C 5E 7F FD 1F DA D3 C1 A3 0B 74 8A 87 7F
 9F 20 A9 1A 86 7A 46 62 FD ED 5D 92 11 92 8C 13
 B3 74 8F F7 73 35 7D 71 FA 10 37 59 9C 10 90 DE
 19 13 8B 42 A9 26 B4 D5 7A B0 F4 83 CB FC FA 3F
 38 80 80 09 13 21 6D 4C D0 3B AB B5 86 20 AF 39
 24 F0 50 21 39 E0 BF 23 7B 23 5C C6 92 DE 04 FA
 91 21 8F EC 9A 74 F1 E4 BC F1 8E 7E 6A FE 8D 43
 44 47 1C C3 B9 93 7F DE 73 50 71 AF E6 E6 97 21
 F7 7B 2A 36 74 8A B9 A7 14 2A B2 98 A0 5C 23 8B
 72 D8 A5 13 CB 21 C1 E9 E1 ED 6B 7C EF B9 48 D5
 74 30 7A C7 FE 84 7B EB 11 8C 64 E5 67 07 47 80
 1B D0 4E CC 0F 98 A6 BA FA B3 43 46 2A 38 0F 2A
 1F 95 62 0C 21 D4 4D 01 3C 88 86 24 06 54 A0 0F
 58 D6 F6 17 EA 58 02 E9 9B 0C D6 09 70 85 53 67
 5D 15 38 3C D5 B1 9C 94 14 E1 71 4B 76 42 59 F7
 0B C2 9C 6A 14 F5 65 73 6D 94 DB AA 34 88 DD B7
 AC 92 9F 74 E1 95 08 81 AC BD 02 05 AB 5D DC F4
 28 E8 B1 FB C3 F2 F9 6A 51 A5 37 E1 9E 92 7E 7E
 56 CA 39 57 2D E3 33 28 41 71 6F 69 35 32 77 50
 09 AC 8E 1A B7 FF AE 02 2C 75 8C 2D 7A 0A 84 84
 BC E8 BB 94 9E CC 80 43 13 2C 72 4C C1 4C 83 B3
 03 E7 BF CB EC F4 E9 32 2E E4 DB 7E A9 B1 48 61
 FE C3 D2 67 E8 90 AA 84 DB 89 64 AE 98 2A 03 54
 D0 8B EE B8 1C 1C 0B 79 24 0C 87 DA 9B 4F DF 87
 07 74 4A 10 69 5D 7F AA 7C 32 0E C3 AB 85 B0 5F
 54 32 86 24 5F 02 17 C3 EC 09 BD E9 57 47 36 13
 E9 52 FE 82 DD EF A3 B0 95 F5 00 85 92 11 3F 09
 9A 5E 13 B3 9D DE 06 AB BC 65 09 7D E8 CC F3 68
 C4 FA B7 66 44 71 62 D4 D9 54 9B 34 C2 93 DB 89
 BC 0D FE 12 FB 95 63 14 9B F1 17 E4 7E F8 C3 9A
 2E B8 4F F6 3F 32 C6 53 A0 63 6A EE 3B 78 5E 77
 C2 7A 9C 6C 39 75 70 03 D2 71 4E CC 34 98 A5 80
 05 EF 71 AB 1E B5 F4 A3 CD 7B D1 D2 1F 9B 0E 2F
 7E C4 46 57 32 9F 85 D5 72 E3 50 FA CB B5 B0 76
 ED 0E 89 DB 4E D6 EB 58 21 C7 84 C7 30 1C F1 6B
 B6 5A 31 19 C6 EA 96 FC FB B8 C6 F6 99 33 E2 55
 FD 72 36 24 3D 2B 7C E7 AC 05 58 A8 4C E7 E3 7A
 A2 3B FE 78 2D 07 9E D1 31 3F 55 E9 E4 33 DA 61
 9E C0 F3 0C 40 82 82 70 A6 DB 3C 38 3B 4F BD 2B
 F5 1D 0C 35 5E 45 2E EF 9D AD 91 3C 5F 47 7E 89
 98 93 8B 08 B3 74 79 80 94 A7 A4 B5 55 2B 13 8D
 26 F0 F1 C2 1A 17 3B 90 98 96 80 C8 05 41 0B 29
 4E 33 BD 7E 9E E1 BF 07 9E 79 71 63 2F 7F 74 A6
 B3 76 E4 15 BB 2E 46 3E 06 92 EE 73 18 91 D8 36
 BD E7 F4 22 34 06 56 30 2A 41 51 5E D6 5D 44 97
 1B 00 0C 76 D6 B0 1A 52 86 B5 23 C3 45 EA 60 73
 CF 5B CD FC 83 12 2F 34 E4 56 C9 C2 2A B1 59 B6
 99 47 63 E0 53 11 3C 50 8A 91 D6 07 DB 87 52 73
 8E 7A 4B 92 A4 C4 BF 71 65 3A FC A7 56 17 9B 7B
 C6 72 9D 9E 12 EA 1C CD 12 87 06 AF 09 0A D3 F0
 D5 05 E3 D5 29 FD 6F CE 8E 04 22 45 23 6B 4B BC
 F0 95 5B 37 BB 98 34 49 49 A0 77 69 26 B5 24 EB
 A5 AC 28 11 FF FC 03 B6 F0 1B F0 DA 37 7E CD 67
 17 C0 F9 90 35 C9 5E 9D 17 FE 2F 2F F4 54 3D D4
 5E 29 9F 7D 89 02 79 23 D2 22 DB 4A 6A 17 F1 42
 A2 B3 F7 9B 4C 72 B6 80 C9 AD 27 56 7B 79 23 43
 41 96 6C F2 B5 0E 26 ED 83 C0 6F 17 B4 C6 CA 24
 D9 C1 D1 0E F5 A7 53 2D B7 C2 E4 D3 5C 5E 94 FD
 4E C1 5C D0 CF 68 D6 A2 E3 FD 3C 2F 0A 9F F6 9F
 19 B0 2E 48 05 4F 18 BB D8 A7 09 DE 04 BB E7 28
 03 13 12 36 E2 DA 8B DB C8 C0 6E AF C7 D8 54 F3
 10 2A 37 CD C4 37 12 CC DB B1 3E CC 1A D6 E6 E2
 9F 1A 47 A4 6D 37 BC BF 62 4D 7F E0 DD 06 E9 81
 69 F2 A1 DC 46 99 37 B7 E8 B0 6B E6 9F E9 55 47
 84 7B 9D C7 ED B3 DD 88 D8 47 4D 79 78 E4 6D 41
 AC E5 38 B7 53 8A 72 FD C1 8A 9D 0A 5C D6 23 01
 B4 BC 45 C2 1B F9 EE F9 58 4F 16 A9 E0 E9 A4 6A
 40 28 D0 05 DC 0D C0 D1 FA 48 FE E9 BB 79 70 C8
 33 94 47 FA 30 7A D8 25 80 8B 1F FD 81 AF BF B4
 50 3A 2E 80 2F 53 34 4E 3A 4B 6A D5 41 69 67 B2
 E0 17 1E B5 3D 15 34 FC BD AF 99 82 C2 52 72 F1
 6E D7 AB F8 2C 9B 9C DE FF A8 C7 5A 53 60 47 31
 B1 E3 08 D0 92 1F 28 DC 25 56 AC AA E7 95 4B 55
 CD FB 64 F1 16 38 04 F3 0D B4 C6 9F B9 8C 36 C7
 A6 D2 10 60 1E 27 A0 E4 5D 6F 61 62 EF 08 CD 9F
 E6 D2 08 3C CC 58 07 8D 83 DF AD F1 D7 CC CC 13
 99 4A 69 E7 BA A2 78 C8 9A 1C 46 2C 96 C5 96 BF
 82 5B 48 26 4F 35 4C FF 30 B6 30 C7 0B 92 50 F0
 0B A6 CC 1B A2 CF 63 75 1E 5A 77 4E 35 8A 73 90
 B1 F3 85 BF 5F 4A 7C 1E EB 77 56 4E A8 B6 C1 D5
 A7 01 46 18 85 C8 F5 6A 71 DF 1C D9 67 EC DC E8
 3E 2B 96 09 59 A3 F3 27 51 EA 26 3A F7 56 FB F8
 C1 E7 CF 20 3B 49 BA 0E 0E 24 4A 5A 7E 75 18 C7
 9B D4 58 8E 28 58 C4 2D 38 1D 6F A9 F3 B5 99 92
 F9 DC 41 AF 5F AD CA 86 62 E6 7B 55 00 17 95 31
 0F 93 29 BD 7E 5F 62 1A AE 4F 46 5D D7 2C 2B BD
 CF 28 3E 74 50 8B 4C DA 70 5B 29 EF 46 77 CB A1
 1D 5D 4B BF 17 4E 5E A8 77 55 11 9E C6 E1 48 DD
 D4 25 99 B6 CD D4 AB ED A0 79 41 78 C3 84 A5 E5
 78 65 0E B5 E7 26 C5 86 D9 EB 51 A9 AE C5 2D 4B
 0A 02 99 83 6F 4A 42 C4 55 82 16 A2 04 F4 F5 DF
 98 2C 25 41 03 97 08 9B 79 58 C9 D7 8A A9 9E 55
 FA BB C1 E0 44 09 AC 20 ED E0 5A 5A E6 67 43 10
 5D 64 B6 46 F5 2F B4 D0 CE AE C9 D5 95 6B 9A 27
 37 ED BC CE 89 D9 37 DE 22 4C 20 B7 13 DD CF 4A
 ED 76 C7 5F 89 2E D6 3C A2 55 0B 9D 2F 80 CC 9D
 F6 7C 3A A8 3D 12 1D EA A3 1A E8 AE E5 12 D4 22
 AC 7C 28 72 03 47 A0 9A 7B 40 F6 54 CF 4A FA 99
 B1 61 5A 0C A1 5A 38 C1 B7 F6 1E 50 AD 11 A0 95
 60 27 AD 4B EB 0D 01 0F 36 56 6D BC B9 14 CA 75
 F1 A1 ED F5 3B 51 BF 5C 03 65 8F 58 6B CB 77 03
 9E 2B 3F 19 27 3F 73 49 51 C3 20 59 01 65 74 E9
 2F B2 1F EF EA 11 F9 6A 90 22 37 A8 98 4D FC F9
 8C 78 6D 60 02 A1 09 D5 F0 70 C9 13 9D F4 13 72
 18 64 7E 9C C9 2E 5A CF 9C E1 BF 0F 15 03 BA 2E
 76 AC E8 D4 97 98 7C 0B 9D 14 93 C0 8F 7A EB 81
 65 56 32 DE 9E B5 BA 51 A2 5F 0F 86 FC 24 6B 26
 59 52 F2 6A 4F B3 FE 6F 74 64 F7 73 C4 5A C1 36
 85 32 42 3E E3 10 AB F6 19 0B 28 AA BD 6C F5 E1
 07 C6 8E 50 E3 28 A9 29 87 3C 19 D7 D4 58 E4 8A
 82 75 76 AC BD FD 75 25 F0 1C B3 D2 AA E1 D4 1B
 69 4E 76 9D 48 C2 78 F5 EC BF 4D DB 85 8F 18 69
 1C CC EE BC 6D 44 C7 95 0D 1B A1 E2 53 3A 31 2E
 71 9E 71 11 0A F9 1F FE 85 2C 9F 05 03 B1 BF D9
 60 CA 5E 89 C0 56 D0 6B F4 74 11 B0 F3 96 A3 34
 49 1B 91 35 4F 25 00 F3 C2 6E BE 35 5F 35 74 C1
 76 AF 6A 9E 32 EB E1 B0 10 40 96 FA A7 BE FC 92
 67 23 9C 17 41 D5 CD 88 A1 66 13 6A 5C 56 FB 36
 DC 27 FC 00 17 4F CC 2C A0 65 80 61 8B 08 6C 52
 49 09 6B 75 BF 3E 64 E6 73 F0 ED FE 91 45 86 32
 76 9C F4 FC CA 24 54 31 0E 13 C5 69 71 D7 83 75
 A7 0B F8 6A E9 E4 CB A9 44 D1 70 8F 45 A7 B4 28
 FE BB 7C 43 2C B2 E8 B3 37 7A 77 EA 9B 2D 37 79
 15 76 22 EA 1D 0A 66 81 01 C6 6D F0 00 F2 36 AB
 91 65 74 23 6F 16 D9 CC 5C 91 DE 14 02 0B 3B 0B
 AA C3 F7 72 49 B3 A5 C5 4B 37 74 73 E5 32 A0 A3
 66 4E 0E 9C 6D 43 4D 87 CC CE 8C E5 FD 27 AF E2
 04 22 76 64 41 43 B4 31 CA F0 0E 35 B9 F0 57 58
 91 C2 8C 98 36 1E AD 2E F1 AC E5 9B 64 29 E7 17
 D1 5B 16 7A 73 2C D7 39 FF 6D 69 CC D7 55 88 AD
 39 16 E9 58 41 0E 70 69 81 11 C4 A5 D2 A5 61 3E
 C5 FF 9A 2B DA AD 84 A3 E0 6A 76 66 DB 29 41 15
 1D E9 F6 6D 03 83 04 70 94 84 17 0F F9 DE C4 8B
 70 D5 33 07 8F FE 59 9F DB 79 A8 CC A2 C7 73 95
 42 72 05 A6 DB EC 3C 52 72 EB 23 E9 E6 C6 5D CD
 A8 7D C3 B8 B9 4E 49 8C DB CF 50 56 93 B4 CC 34
 95 83 D9 78 28 17 06 F8 0D 7D B1 CA 6B A2 40 53
 66 C7 63 1D 46 A0 B1 6C 98 C5 AE 8E E0 8F 16 DF
 E4 2F 2F 05 95 81 B7 61 EF DE F3 2B 9A D4 6F 68
 7B B6 8E FD 84 62 0E 35 09 01 9B 08 28 92 F3 EE
 7C 3F 5C 3B 3B 4C C0 4C 98 A1 32 F5 16 5B A8 51
 74 00 8C 4A 2D 68 02 BB BE C2 4A E4 2D 01 93 A8
 EB 1C 08 AC F9 80 D2 2F A8 D9 03 12 2B 51 3C 54
 5C 0F 19 CA E5 61 42 9B 32 C4 71 B8 6C 44 9D FF
 A6 CC 33 1D D1 34 A8 2F 55 E8 29 93 0D 56 83 25
 AA A9 B3 1C 79 15 62 10 D0 5D 65 92 D9 F4 0F 30
 70 38 43 E7 04 4C A0 CC A0 40 3F BC 41 FE E2 88
 3A 67 84 39 08 9C 11 E4 5E A3 2F E3 2D F2 84 6A
 6F EC 64 13 82 AB B5 B1 FC B2 23 BE FD C7 96 00
 84 79 2A A9 0D CD B1 6E 0D DD 6B F4 40 51 C2 DE
 DA 95 BA 4A DD 6F F8 BA 48 4B 2D 9E 1F 12 E3 CD
 68 94 79 1F FB 26 27 6D A8 A7 50 ED C0 60 23 9D
 BE AB ED 86 FB 53 01 8B E0 3C 5E 8A 86 27 4A 24
 00 D3 02 07 F0 7D 5C 95 8E 8E 5F 5C 4B 4C 06 1C
 2C 5D 48 DD 86 E9 6A EA 43 37 D7 1D CC DC AA 20
 FB AB 31 2A 1E 59 59 E5 88 53 9C 6F 4D 8F ED 7F
 B4 86 93 C1 9D 74 C6 AF 03 AA BA 54 BB DD 23 B1
 36 50 E4 B9 9C 4A B0 67 20 26 DF 88 4F 57 43 F8
 E4 B6 32 29 27 AA 13 85 39 EF 26 13 9C 0C 73 E1
 6F 16 D9 BF A1 49 91 96 1B 7B 68 F2 9C A8 34 9E
 00 E9 1F 53 37 3D 0D C6 E8 CD 90 EB 8B 17 10 95
 F8 DA AE 11 FC C7 0E 7D 68 3D A0 17 67 22 BA 56
 CF DF 32 26 AE 99 89 01 30 A8 EC E7 FF 94 92 59
 5A 3C D0 53 65 62 AA CC 87 10 A3 E1 CD 97 31 74
 14 DB EF C4 13 DB F9 A4 FD F0 E9 3B 62 AB C3 02
 C4 DD 25 4D 44 8A 69 5F 2A A0 69 8B E3 7C 29 0C
 60 CB 8B 2D A5 C0 31 C8 1A 42 F5 8A B1 BA 44 7E
 34 E9 8D 51 72 26 B0 0C 20 36 F8 2F 47 AE E3 22
 2A 56 7F 01 A5 6E 68 EE A0 3C 2C BA F1 B8 9A B2
 52 A8 BF 79 F6 A6 A8 85 00 63 30 8E A0 32 70 1C
 5D CC 30 2C E6 2C F8 BE B2 83 62 0F EC 36 9A 70
 B6 D2 16 33 B0 75 A6 86 6B 48 FD F0 76 48 7F 45
 C4 3E 89 D2 7B DA 40 4A B6 D4 83 0C 0B A4 5A A4
 54 21 42 2F EB E5 95 46 9A EC 0D 77 DC E7 84 A1
 02 B3 10 88 8D 15 58 8F A0 26 A5 AB FF D6 6E 0B
 35 A6 38 A8 F8 9D E9 10 5D B6 2A 00 F2 B5 F7 B5
 54 E5 99 98 9C 28 12 BB 7B E6 BE 77 77 97 FC 94
 EF 82 94 E1 4D 91 DB 9F 63 52 14 A3 76 0A 33 73
 5D 63 80 0C 44 CA 45 EF 60 C6 80 A4 39 BC 21 A5
 DF F5 00 75 33 9F ED 60 89 84 BA 6D 56 DD 45 C3
 9C 5C 36 F5 D9 F3 12 DF 32 CC E7 E9 4E 4E 42 D4
 14 9F 94 C3 6F B7 64 36 AE 1F 38 6E E3 9B 46 4D
 CF 93 D2 C1 5C 72 71 96 3B EA 0B 7B 11 AB 7D 0C
 87 08 A0 5A B6 0A DC 83 C5 8B BF A0 70 5F 12 C6
 C8 C2 28 35 24 9A 5D DE 4B 4C D1 E6 0A 0C 13 3F
 6F 21 CF 45 31 11 DE 10 98 C2 D6 83 27 90 31 62
 94 2E F4 E1 B6 3D 8D 38 A3 49 ED A2 68 03 75 E4
 8C CA 74 23 AF 7E E9 E2 1D 17 48 01 65 D1 B9 82
 8F EE D6 BA 29 1C D8 16 82 97 6D 2C 65 E3 1F 7A
 5E 10 BE E9 CE F2 E7 EF 2A 5A 77 89 38 7F A7 DB
 35 A0 80 C3 9E D7 F0 87 04 0B 0B 82 70 92 D1 1E
 9B 31 7A 33 C3 13 F8 1B 30 44 9B 11 24 87 34 B5
 4A 32 14 6E 2F 18 E7 1B EA 6F 62 B8 41 3B 40 47
 DD F5 A6 38 D8 CD FA 6F AB B8 4C 84 39 92 1A 4D
 54 4E D1 83 AA BC A4 F8 C9 8F 48 9F 8B B5 32 CE
 74 A8 73 86 17 B1 A8 83 EE 1E 59 2F 12 F4 4C 1A
 90 E6 B7 33 63 54 F7 D9 35 03 20 A8 FF 10 72 7A
 46 20 FD 97 AD 23 0A D8 61 1C 02 11 2D C8 69 1E
 B4 FE 69 9D C1 46 AB 73 82 24 D9 44 D7 AD A6 A2
 D0 AF CF 59 4B AB FE 0D 73 6E 35 F5 2A B7 0F B4
 71 AD AF 46 B9 9E 8B CF 3C 6F FB 99 BA 03 54 7B
 A3 8A 4F 32 31 67 87 60 8B 5E C4 4E 15 8B CA EF
 5B 93 44 6C 3E E4 30 18 08 C2 90 38 FA 3D BF 2F
 28 91 9E E4 4B B4 E2 34 09 35 36 83 D0 05 DE 04
 C5 09 9C 19 6F 4D 73 90 4B E1 D4 1A 94 23 76 4F
 25 AD 23 67 D7 A3 0B 96 87 65 EB DD E8 82 40 96
 CE A8 08 65 DD CF C8 A1 A6 20 8E 73 ED 87 2E 6B
 E0 9A 70 03 4D 79 68 53 09 EF BD 44 FC CC BB 00
 79 C4 BF C4 9E 63 1E E7 46 E3 24 F6 1A 2B 11 71
 C1 C7 85 D3 60 26 85 8A 2E AB 48 18 38 B1 74 DF
 C0 B1 43 8E 4F 8C D2 AB C5 39 EE 4B 89 6E CC 0F
 17 93 E9 94 19 B5 0A 58 09 F4 C7 95 C2 A8 74 A3
 87 54 16 4B 34 79 7E 0B D0 51 DB DD 7C 69 2B 21
 32 E8 63 D8 25 FF 63 05 93 4B 1F B2 FC AE B9 A7
 47 03 6E 78 28 C2 F5 89 A9 FE ED 74 1B D2 07 44
 B8 C6 FC 9C 91 86 4F E4 88 AA 89 36 7E D3 76 7C
 31 9C 1C 4D 2E B4 D1 41 95 AD 71 28 24 2E 0F CB
 D1 86 79 07 4F AB F5 4C 62 67 86 73 4A 76 A1 34
 19 66 F8 EE A8 16 61 66 72 88 80 8E 1B 88 34 D9
 7A F7 B3 11 24 C4 3A D5 F9 2E C4 00 18 EE 58 48
 53 96 35 38 AC F2 9A 65 4C 88 D2 5A E8 35 76 FC
 AD 4B 26 72 7B 41 7D CF 67 05 A4 FF 5F 33 68 1C
 9C D6 56 B2 40 B6 4E 89 A2 0C 24 F1 D5 32 8A 6A
 8F AA 01 60 CC 06 B7 3E 2A 5E EE 62 E7 CC 01 2E
 95 09 FA 7C DF 6C 6F D7 3D F7 D4 E0 2C 37 23 EE
 27 EC 27 37 BF 43 F8 B8 42 EC 9A 92 70 94 0B EB
 D0 E2 90 6A 65 C4 23 F4 EA B1 9A 29 9E F1 C5 CD
 31 D0 21 AB 09 1C 14 30 62 0C 46 B2 94 31 CD F2
 CB 45 04 39 C0 11 6A AE 35 B7 CB EF 34 B9 3F 9C
 71 E7 B4 90 4D C7 0C 85 EB 12 70 F8 CC D7 00 14
 87 48 F1 E0 0C 0D CB 51 05 E0 CA AB C3 DD E4 1A
 AA 14 AB 44 E7 17 9C D5 96 C9 D0 D5 02 0D 08 7F
 B6 C3 9C EC 1F F5 DA 0B C0 5F 19 1F C0 03 D3 50
 D7 D9 4B 5D 5E 25 BA 04 F5 CA 73 E8 84 0B 5D 72
 E7 1A 65 E4 19 A3 E5 18 F8 A3 30 98 95 C2 8B A5
 83 40 D6 6B B1 94 6D 95 F1 7D FB 97 7F 74 84 9E
 69 4B 6B 55 5F 29 05 7C F5 97 EB 2A B7 E1 F7 8A
 8D 2C CF 5F 4F 32 7C 4E 48 5E 60 C5 DA E2 C4 4B
 EC C0 95 7C 0B CE B8 2E 1B 14 33 AF 3E 50 A3 02
 94 EC 35 9B 26 F9 84 E1 A2 4B 8A F9 9C C1 8A 0E
 51 01 9F A6 F9 1B 84 8D 0C 6A 13 28 4D EF A4 4F
 C0 4A 79 3E DC 5D 35 3E 95 CB 61 4A 60 A1 CB 88
 18 F5 CF 58 30 11 DE 37 86 25 74 F6 B4 35 74 3F
 23 CE C2 92 52 61 10 B1 B5 24 57 DD FE 30 53 B0
 E7 A0 75 30 84 22 5F 8C C0 EA A0 64 96 12 23 0F
 43 F5 69 97 EA 68 8F B7 C4 D9 D5 8D 4C DA 05 3C
 7F E9 B3 1F 56 42 B7 B5 FE 3B FD AE 5E 79 BD 97
 31 08 E2 4E 12 E7 77 AA 71 4C 0F E0 29 20 BE 37
 CB C1 61 63 32 66 C2 A8 AB 8E 2F D3 E3 92 F6 57
 F0 56 C2 A1 D4 1B FC D0 CD 58 98 F4 6C D7 42 A6
 55 61 15 A1 FF 60 E7 95 F0 52 F1 03 A1 8D 7A B7
 8A AF 76 72 89 70 8B B5 CB C1 04 44 F0 3E AC 9D
 01 52 FB CB 43 94 B3 A8 69 84 BB C5 26 3A 40 8B
 76 9A 82 B9 2E CA DD 4C 11 0F CC FB 05 87 5A B6
 95 7F E5 9E D1 E6 74 87 C0 8B A4 D7 1F 65 3D 6E
 03 B2 62 CF 5B 5F E1 BF 58 23 74 89 47 CD 06 7E
 1F 17 43 40 DF A8 BF 57 E0 AA 01 6E 57 E3 F8 3E
 EB F2 63 D4 9C DB 5A 44 71 C1 4D EE 5A 64 02 6E
 0D 8B 72 B3 76 8A BB 6F CD 33 E6 14 7F CD A1 E8
 92 22 4C D7 8C D0 06 AA 1D 4C F4 94 D0 4F 01 67
 BA 4E 1D 14 2E 31 44 BA CB B1 87 AF 34 92 04 1C
 FE 5A 02 B3 05 5C 1A CD 5A 2E 5E 1A 94 BD 71 D5
 27 EC AB 37 A8 44 BB 29 5C F6 CF BF 82 76 49 CD
 8E 7D 35 45 5F 19 88 36 44 6E 3D 15 BD E9 04 D5
 8A 4B F2 D7 C8 B8 72 DF 04 E3 CE 50 B0 33 AE B4
 E8 29 C6 41 D9 7B 24 41 5A 31 6A E7 43 A6 E7 17
 03 30 6E 90 C6 5C 68 B9 5A F9 B1 3C 06 F6 CA 44
 F5 BA 85 B2 9E 83 D0 12 06 A7 FB 44 BB 29 B3 44
 69 AC 84 49 F7 2D 04 91 F8 DE 0C 68 1B 45 3D 01
 6E DC 46 7C A8 14 E2 7E 18 2A 84 76 BE 63 6E 5A
 BA FE 09 C4 3B 72 C0 2C FA 5D F1 82 F7 E2 AB 64
 A7 68 7A 25 80 CF A6 5F 1B 0B 62 E4 9E 59 70 4B
 CA C4 75 57 73 32 57 E5 CF D7 30 A1 9C 88 57 62
 39 D2 D2 CB 4B D0 96 C7 12 12 68 0A 97 BB A8 63
 15 B6 94 9D AD E7 65 18 79 B2 78 3E B5 59 A0 E2
 BA FB C8 CA 07 A9 BA 75 A1 88 FF 65 17 30 28 E1
 67 29 82 76 78 D8 3C A9 76 58 1A 83 0D 00 E6 4C
 46 D8 9B 89 3C 6F EC 68 53 BF 71 D7 A1 CC 70 54
 CE 53 CD 8C 4A 71 54 A5 32 C1 1D A4 DB BA 81 34
 55 E4 B0 C1 42 C2 2D 93 2D 77 17 1F 94 2A 60 A8
 D3 01 DF 03 EE 52 D8 38 11 54 F1 B8 37 A1 C9 43
 33 36 60 90 4F C5 3C 27 74 0B 0A 8D 2C CF CA B4
 6D 78 23 6E E6 AF E2 76 B8 08 6C FC 0B C0 35 4A
 90 B9 12 82 7A D9 F1 7F 08 70 2C 72 6E 09 B4 C5
 A2 95 85 69 FF B5 6D A1 41 89 9C C0 55 4B 3B 6A
 AC 59 83 AA 8C 99 E5 30 91 40 43 B7 67 C8 12 B8
 31 CC F5 E1 F6 88 B9 96 CE 40 34 A7 F9 98 8B B1
 15 0E 1D BC 7A 35 76 79 9B 15 66 87 14 86 08 A3
 5F 80 61 6D 9C 42 CF D1 6F E2 EA DB 54 F6 1A BF
 7C D8 EA BE 26 73 7D 8C 0B 82 53 71 D8 40 10 66
 05 77 A2 DA 76 CC 97 3E E4 F6 D8 42 E2 13 86 D3
 1F 6A 89 E3 D2 59 50 26 FD 00 4C C6 B6 E0 CF D1
 6E 6C 16 DD E3 52 B3 2F 0E 77 82 4B D5 E7 FC 68
 66 7D 12 3F 87 C0 53 9A 7B 09 CC C5 D9 B6 39 0F
 37 05 07 8F 32 E3 8E FC 15 02 1E 89 0C EC C5 8A
 49 B4 DE 51 36 DD F5 41 63 74 17 5B 0E 5B CD 73
 DD F7 08 CE BF 05 83 8F FB FB 9E C2 54 9E 32 9F
 75 09 79 0E E8 C1 57 C8 CD 45 01 1D 03 62 72 D5
 40 B1 28 9D FB 08 0F 14 98 72 2C 2B BC 4E 78 74
 91 07 B7 E6 41 65 E7 01 8B 43 ED 75 BB D2 81 DC
 86 69 D2 54 B8 1C 84 6D 20 D3 59 84 00 41 96 A0
 56 8A 5E D1 35 C4 1D 2A 35 F6 B2 C7 80 DD AD 78
 85 8F 8D 8A E8 D3 95 EA 05 48 BE 18 F5 74 BD 2D
 A7 C0 08 00 C3 AB 1F FC EB 29 97 1B 16 33 4B 00
 D5 67 D6 40 CE 94 D0 AA 68 6D 6F F8 EC 99 5B D7
 2F AF 2F C2 79 B3 2D B1 9A 26 E7 2A 2C 5A C0 87
 D1 BB 2D 40 42 64 D2 14 79 C1 31 05 9D 53 5A F2
 90 AF C9 A8 CC A0 98 14 0D 9D AA 84 58 8B 22 DD
 48 6D B3 4A F5 99 02 5D D2 EC 7B 4A FC 25 E9 B7
 F0 A2 F4 A5 32 D2 31 31 10 D4 37 C3 B0 71 36 DA
 EE D5 82 FE 9F FB 41 84 89 B3 14 14 FA 9E CB 97
 F9 0A 26 D0 BF 23 01 77 1D 90 64 00 F1 C4 78 4F
 3F B4 7E 77 A6 88 64 4A 9B BD 1A B1 C2 4D F4 3A
 B5 43 54 37 74 5E DD 7E 1D 27 21 9D CE 2A B1 B3
 07 65 AF 1E 32 E5 C9 0B 44 A2 C6 BE 73 23 36 1E
 CC 8D 21 09 3B F2 45 AF C8 B1 8B 6C FA CC 9F AD
 DA 79 A6 E3 21 59 15 BE E1 7D 70 8C F6 8B 0B D1
 49 DA DA B5 FA FC 26 91 BC 8E C8 09 D3 95 48 C0
 B1 DE BE EE DF A8 0F DB BF 34 4B 80 0F C7 13 C9
 FB 88 DD 41 53 DD C2 0C 8B B8 FD A6 CC 12 84 4D
 82 2B DF 0A DE 80 71 39 F1 FC 88 28 74 A0 88 09
 32 37 96 F5 E2 51 A7 4E AB 91 B2 0A 33 8E 1C BF
 E0 DF D1 51 D1 4F CE 75 48 97 5E 4E AE 9E 45 B5
 7F 25 5D 31 1A 7E 0B 50 8E 98 B1 E8 70 E4 6E 76
 78 3F 97 72 2B D9 80 43 6D 35 62 0A 79 D8 18 06
 33 42 F0 D5 FC 2B D7 0F 23 66 48 2F F7 3F 87 03
 F7 E6 02 F1 DA 4E 4B 37 A0 56 D4 F1 C9 A6 1E 32
 C2 65 FF AF 65 C3 8E 2C 01 46 86 05 4C 99 F3 C9
 A5 A7 A0 66 1E CE D4 9B 12 E1 27 E6 EF 0D 29 4B
 AD 45 24 7D 5D ED E3 D2 E2 9C 21 68 59 86 C3 51
 A7 83 5D 0D A3 B5 17 D7 69 DD FA CD 30 90 51 16
 8A 3C 02 4C D1 19 96 6A 2C 7A 8D CC 73 94 C6 68
 D1 DF DF F8 E9 DC 1D 73 D9 99 C4 C4 BF 5D 61 12
 8B 1A 75 99 0A 8E 86 E6 25 18 E3 23 84 2F 8E 2B
 11 87 5A 73 E0 88 7D 23 2F EB FE 60 0D 43 DC 82
 9E 28 48 09 87 FE E3 96 DF 7A 7D D9 50 B5 2E 53
 DD DA 5C 28 28 71 95 2A 2C 84 9E 0E 1A 84 DC 44
 20 04 22 96 95 08 48 9E A2 AE C4 65 B6 96 5A 0E
 81 5E 85 E5 5C 11 3D 4C 60 72 9F 36 15 B8 F4 5E
 AF 36 2F 12 57 84 DE 18 6A 3D 1E 60 02 F7 5A 5E
 7B 60 C4 FB 38 E5 12 7B 20 48 8F 91 51 C1 3B 66
 C0 74 DF 0C D3 B3 23 EB 06 28 C7 AC CA 5C 91 05
 98 93 2A F5 15 EE 7A 34 44 11 2F 8A E8 95 B4 54
 A4 FC 6F 7E F7 2C 0F 20 18 BB FB ED 7E 3A B0 7C
 48 EF B1 24 13 DE 27 27 20 9C 1E C1 D9 B1 79 D1
 F6 EA 34 C0 5F B2 49 59 61 4A AA B4 89 4A 36 FE
 DC 4F 19 16 15 5C C5 B3 3C C9 87 E3 FD CA F1 EF
 9B F6 CE 4C 4E AB EE 35 AE 05 39 F0 32 7D F4 BE
 61 12 4E E4 0C B8 3E A6 84 7B 56 2C EA B7 89 60
 DB C7 E6 9E 99 0C 2B 68 1D 81 F2 77 30 30 90 59
 86 A4 94 08 4C 8C 42 07 A8 C6 4B C0 0B 97 2F 90
 C1 06 BB ED 69 97 87 EB F6 55 DE AE A4 C0 E4 55
 69 56 E8 FE 2A 81 59 C8 27 93 53 EC 07 14 1D 89
 42 03 0C 90 4B 74 F4 A7 B9 FD 4A A0 EE F2 60 48
 06 91 FB 24 C7 0C B4 28 AF C4 75 6D 45 B6 F7 E2
 DB C5 6A F2 B2 E0 34 B0 20 81 66 C1 79 A6 D4 0A
 43 04 A4 77 BC 28 7A AC FA FC 66 43 66 84 B0 D0
 CA 2D 19 B2 F0 2E 60 4F 34 0B FD E6 28 40 94 AF
 F5 62 68 E2 86 13 06 80 29 B3 1F 70 18 96 A4 7A
 0E B9 9A 90 25 53 7C CF E2 04 58 84 BD 1D 89 4B
 E1 79 70 02 41 75 92 85 23 61 80 71 F5 FF E3 10
 A9 9B 79 CB 88 1C B3 68 EE DE 6E 1D C0 90 1C 98
 E9 B8 60 C2 A0 CE 30 AF 23 7E E6 58 9E 90 78 94
 B1 0C 69 6B 0C 91 53 FE 41 4F 76 B2 6A 54 DC 93
 DB D9 12 D1 01 7E 27 2E F0 62 13 33 1F 20 72 A6
 D3 4C 50 01 55 A0 38 7B 20 75 AB CA 4E 15 B1 C3
 6C 14 EA FE 06 11 9E 06 EB C5 82 A0 E2 4E E1 7B
 38 DB AA 6D E7 B6 58 8C A6 B1 C9 38 50 AA B9 6C
 C5 5C 09 D4 A2 50 A4 E0 CC 4E D7 58 F6 14 54 82
 50 15 C6 CB F5 38 18 BC 09 8B F8 1D D8 58 23 84
 D2 1C 54 77 E8 49 78 D3 D8 DC A9 CF 90 95 33 8F
 02 25 10 89 7A 94 D7 A2 AA 92 7D E0 52 9F 48 47
 D1 E0 03 06 9D 56 04 EB 7C E5 78 4D 0D C7 10 94
 7C FA 3D 5C F8 3E 39 64 7A 92 1F D7 42 47 48 59
 BC F6 B9 E1 22 B0 01 49 DC 60 5D 2D 44 78 B1 BF
 6D 79 D7 C9 67 8F 39 AD 85 3B B6 84 E4 0C 39 5D
 5D 02 62 C7 73 88 5B 95 60 F6 71 85 13 2C 5D 35
 D2 83 4B 2D E3 80 C3 AB 0D B9 8C A2 DD 9F 29 65
 EF 94 B9 7A 3E 80 12 52 4B 91 C5 51 DF 1E 9A 29
 A0 CE 2E E3 69 69 81 24 68 69 3E 7C 66 7E 48 A0
 DF 2F 38 F7 CC D2 4D A6 94 02 84 2E AD 96 B8 22
 93 25 AE 3E 85 3A 78 3A B8 62 F1 9E B9 8F 4E B3
 F5 38 55 A4 B5 8E 0C B5 6E A5 08 53 32 61 19 8F
 0B D9 0B 84 D3 B9 F6 79 DB D1 A0 29 70 8C 9A C4
 1E 4E 82 1C F1 46 7D 1B A1 36 F2 18 8B 24 C0 D9
 28 E5 9B F1 98 AF 77 71 AD 46 BD 01 3B 02 DE E6
 38 93 B1 C9 B3 7F 28 72 A6 3C A3 24 AE 9A 56 26
 5D 58 43 12 C5 AA 41 8F F9 3A 51 85 A8 EA 09 E5
 CB F9 1E F0 20 D3 7F D4 6F 59 2A CA 2D E5 00 53
 3F 6A 50 D2 88 93 F6 71 DF B9 C2 DE A5 51 E3 CB
 4F 9D B2 6F 1F 15 97 30 C8 C8 DC AE 74 DD 75 27
 EE CF 59 50 EB 00 2B 62 CC BD D5 EF DE B7 00 C2
 E7 6C 46 32 4B 19 04 67 C9 FA E4 02 7E CD 12 E8
 DC A9 BC 71 C3 61 7D 6C 92 FF AE E9 30 AC 4A CA
 E4 E2 96 EE 31 4A 42 05 89 20 25 AC 8E 36 B4 F4
 D5 1B 96 EE 3A B4 3D 8F 37 16 4C 79 82 63 6B 9B
 44 4A FA 3F D7 60 64 60 35 DC DB 78 4E D7 02 05
 3C 6C 59 18 61 C7 19 1F 29 8C FA FA AD F9 07 F0
 9F 64 11 2C ED FC CB CE 38 4F 56 72 CD B9 15 2E
 79 87 22 61 B8 D0 DA 7E 98 C6 1F 66 AD 03 6F 28
 01 27 05 30 8F 1E 05 35 1F 27 CD 51 61 43 41 96
 A3 11 C6 C6 7E C7 25 10 C7 40 8E AD A2 D0 27 76
 0C 81 BC 13 3C CB B1 77 36 59 ED FB 78 31 6E 89
 80 03 31 23 3F F9 55 36 CF 2D 28 91 69 17 EA 60
 E6 8E 8B F8 B6 D0 2B 88 17 FE 07 90 3F 75 3E F5
 54 B8 C4 5F 7A CB 1F B6 35 64 6D 2A 89 BC F6 21
 C0 AA 80 49 4F 30 7D 3F 86 C5 29 88 B7 36 B1 B5
 5A 15 31 24 BF A0 12 F7 DD CE 9B 32 BA 90 F5 97
 31 C0 FF EB 49 F9 16 BE 5B 89 AE 83 6C BB 23 B8
 2E F9 CD F3 F2 9C D2 9B 8B 73 2F 8A 28 C4 31 01
 FE 18 74 35 AA 59 03 DE FF 85 5C 18 93 15 3F A4
 A8 D0 E1 6E D6 82 FD E6 ED 3B 76 B9 29 6E 76 10
 C6 16 84 EB 39 42 CC 74 F6 36 65 53 37 9E 76 73
 9B 5C EA E5 B7 E7 29 05 A3 AE 9B 8C 5F 59 22 D5
 1B 18 CF 9E 3D BF FF 90 5D C2 05 99 2A 25 20 5C
 B9 B0 83 09 41 DD 8C 63 C9 88 71 63 81 12 04 64
 BF 63 F1 CD 12 E9 4C 44 3C A0 64 6D C8 D1 2A CB
 E7 37 18 C7 7B F1 12 72 36 D3 CC A8 4C 85 2D D5
 02 2C C2 C5 48 F3 CC E3 8B FE BA 3D 47 D8 85 F3
 07 27 39 C1 7F 5E 2A 1E 97 6E CF E1 EC 73 8D E1
 06 40 44 A6 52 E8 C4 C3 DB 56 13 17 7E D2 9A FB
 AA DF 09 92 E3 34 14 33 4A 72 A8 69 AB 72 FF FD
 8A 53 4E 0E D9 41 6B BC BD 1F 0C 27 AB 24 34 F7
 85 51 42 81 54 4D 60 A7 32 97 15 57 F3 7A C2 9B
 71 1B 81 2B 30 B5 CA 5A 47 E7 AB 24 DC 66 D8 AC
 1D 8F 34 B7 D1 6E 29 93 E8 15 36 3A CC 33 55 65
 4C 9D E9 75 F1 81 F2 36 66 B4 78 42 4D 43 C3 1B
 D5 AB 93 71 99 34 28 1B 2F 14 1D CB 1D BD 7F 4C
 93 83 0E 35 42 53 03 2D 36 CD 01 8B AC A6 73 5B
 BF FF 6A 9E 2A 16 AC FB FB 86 DF 27 EC 7F C8 54
 F8 79 06 4E 47 EE B9 A5 A0 4A 68 40 DF 9B A3 FA
 F4 B1 C6 76 8D 58 A4 6B 14 4A 91 E4 EF F5 E7 27
 7C 3A 64 09 0F 9E 7C 1B 17 A1 FF 31 12 64 FC 60
 10 42 27 7D 7B 5A 4A 6A 28 19 F8 58 B5 4A A4 52
 8C 12 91 07 76 B2 70 FD 41 46 34 CC 0A 72 E9 58
 E5 2D 91 D0 78 67 73 D9 38 AE B7 DA D4 6F A5 54
 18 89 10 49 D6 D8 25 73 B3 59 B0 7B F3 79 E1 CE
 C1 05 C2 3E 42 E0 41 12 02 94 5D 42 07 56 C3 13
 0D BA F8 16 BE C1 9F C7 DF 29 34 52 DE FA B5 A1
 AE 2D 85 A6 51 FC 91 16 5D DF A8 8D 70 78 00 91
 E8 56 BC 2B 0E A8 8D 27 A8 56 B9 5D 79 8A BA 20
 46 A2 48 92 9F 3F ED 1C E7 45 A5 27 3A CD 6C 89
 C8 24 76 AB 38 7B 75 17 71 84 20 EA 67 DA 2C 0A
 61 A2 9B 84 D6 66 D3 FE 13 41 32 4B 70 E0 1C 52
 C3 3E 2C 8C 8D 64 6B 71 34 A0 67 56 19 9D A7 4B
 86 17 DB A6 57 2A 88 A6 F7 C2 59 EF B1 02 A5 78
 13 BE B3 9E F2 D3 EB D4 AA FE 73 12 29 9B 85 44
 7B 4E E8 7F E9 A4 B8 56 A2 F0 89 5B 01 78 19 C3
 43 04 D6 16 F5 17 1A 47 A8 1D 60 2D 7C B3 46 F0
 0C 5E 51 BF 58 19 DC 90 76 5D D9 3A 20 F3 AA D5
 2B 70 51 46 B7 5D C1 C5 03 B9 B3 30 5B D1 44 4C
 B9 16 0A CE 5D 2C 77 62 59 09 F0 40 FB F7 FC 7F
 D2 A8 1C FA 9F F1 24 0C 86 90 27 64 41 DE 71 32
 CB 74 F5 1B 67 57 BD CB 3D AC 29 3F D3 5D 88 E3
 D2 CF 55 14 A7 58 2E FA A3 37 64 07 B6 3C 27 FE
 6D 5C 78 0A EB 9F 95 B3 19 52 98 CE C5 E1 19 12
 43 83 CC 97 3F 0E 49 4F 79 AF 89 6F 7D F6 F5 59
 30 AA 2C 4E 39 B5 4E D0 CC E7 FD 97 95 4C 5C 3E
 83 B8 3E B3 96 9F 42 3B CC BD 7D 65 DB D7 DC 0E
 EA 44 D1 31 02 80 EC A6 8A E0 DD 8F 23 E7 B7 0D
 72 44 7E 2F 12 1A 0F 63 04 70 85 C7 72 D6 A3 89
 60 68 31 DC 0D 93 28 3D 59 7B C0 DC 0D 9C 94 27
 E5 D1 6F FB 3F 3B BA DE 5C 40 AB 12 62 61 62 A6
 01 6A C6 A6 5C 62 CB 7F 7E 29 26 10 EE BB 11 3D
 9A 76 F0 84 4B 0C 18 E9 BC 1F EA 25 81 48 0A 39
 B1 F5 03 94 5C 93 39 28 D6 78 A7 1F 96 89 97 58
 C9 A0 ED 0A 82 38 CC E3 D1 45 FE 2F B2 4D 82 63
 DB 4D 72 28 D4 1D 2B 16 5C E7 DF 0D 5D 0B 46 3A
 32 FD 0A A7 10 0C 3D 06 32 65 51 F7 CA 66 3B A8
 BE 4C 37 56 23 6E 03 E1 99 89 1F 2A F4 4F 2B 3F
 6B 08 8D 12 ED A9 A7 95 1F 26 2A D0 54 DE B8 F8
 36 13 7C EB 77 C0 A8 65 A8 25 FD 63 78 85 36 6A
 46 FE B3 05 68 8E 28 AA 00 99 E6 DE C4 23 87 5C
 7C F9 C2 F4 A3 43 BA AA 0C 38 9C A9 FF 9B 6A 6A
 E5 88 09 42 CA 88 B8 BC 21 D0 BC C2 3D 63 18 25
 98 7E 67 2D 67 95 19 F5 5D 19 AE A7 92 0E 85 D8
 15 25 9C 6B AE FA 65 0B 68 E0 CD F3 7D E1 43 0C
 DE 29 AD 93 86 42 89 C6 FD A0 1B 76 43 8F CA B6
 97 F7 23 EC 4D 08 21 80 9E AB FD 0F F4 03 BD 60
 28 B0 27 BB 23 C8 BE 5E 24 50 A7 A8 5F E3 77 FA
 D6 F5 68 73 67 BB 7C 89 FB 19 DD 32 C7 72 C8 44
 4D 9D 1F 37 9E 5B 56 FF C7 F1 DB D4 15 C2 E6 B2
 4B 5D 0E 47 45 89 26 53 7A 2A A0 14 52 F0 7D FB
 9A BA A0 BF 91 5B 30 A0 3B 9E 6C E8 50 FE D5 3B
 4C 01 B4 DC EE CE 34 4D 14 CA F4 FD A8 35 19 C4
 49 71 F0 37 79 CE 31 5D 98 D1 19 37 D0 43 A4 7A
 19 A5 F4 05 CF 97 B8 67 2E 87 21 59 53 AA 46 4C
 46 F7 88 E2 E0 D1 15 BB FB B7 AE 5F 43 6D 54 D0
 7C 23 34 FF 17 8B EA DB 83 45 52 8F 5A 02 5B 0A
 DB E4 89 C7 27 61 50 98 61 85 A7 C0 4B 43 C1 C6
 BA CD C7 36 76 41 ED 1B B5 56 1D 1E 15 6A 4D B7
 13 2F 8B 84 98 78 58 AA 3C B7 34 5B 5B 7F 77 35
 50 7B F1 2E D6 E7 13 AE 17 D8 F5 28 09 6B AD A8
 2B C3 B6 C3 C3 8E 9E 75 B9 00 59 C9 1E CF F6 79
 01 7F 43 6B 24 F7 29 8B B9 65 15 77 CD F1 F9 44
 C2 D6 A7 B0 30 2B C1 D7 75 92 9C CD 90 85 DD 0F
 D2 EC DE 0F 51 F6 54 C4 50 C0 D6 9E 76 0D 94 81
 27 06 BD 34 0A 72 73 53 F4 7C 48 D1 7C F5 8A 70
 D2 CE 66 63 DA A7 96 6D 82 B7 31 90 B7 95 AE 14
 18 99 BF 9A B4 F8 68 3B 1B 86 46 DC BD BD 17 58
 FA D0 D0 4B 87 B6 22 86 59 5F 10 8E B7 7D 9C 48
 90 38 76 87 FA CC 09 FF E6 63 9E FA 6A 2D 95 B4
 24 41 66 37 8A 05 95 D3 5F E5 34 6A 77 7B 41 5B
 A8 6D FA E0 D7 65 EE 1F 34 0D A9 DD C7 F5 68 29
 8C 2D 02 D6 2B E1 11 6B F5 8E 97 BB DA BC C1 2B
 5A 81 4F A3 E4 F4 15 12 AA F3 35 F8 81 E7 20 99
 58 F5 5D 06 B7 E8 91 B3 75 91 50 D3 0D A8 68 CC
 A3 72 E7 99 F2 0B E8 5F BB 99 31 EE 4A 99 7B F2
 9F E6 B1 E7 2E EB E1 22 AA CA D1 F2 0F CD 20 B3
 94 12 73 6B 43 D4 B4 1E F4 EF 25 F1 CD 86 5C 36
 BE 3C 83 1E A3 FC 6E 0F 0F 36 ED 1C D7 D3 A0 0E
 3E 96 62 76 ED 98 BC BB B7 C9 5E 7B 5A EA BF 5B
 7A 6C E9 EF 9F 7B 72 32 DB FA AF 67 56 52 16 D8
 5F 5B 81 17 BA 15 EE 46 F8 71 50 47 6E FD 53 5F
 48 33 60 DD 61 D9 36 F2 D2 52 3C A0 23 75 A1 56
 DC 56 AE 0F 50 8A 3D 93 44 2D 36 56 CF 5C 71 23
 01 FA 00 14 A1 2E 80 4F 69 E5 09 07 47 C0 05 D3
 A4 A9 6B AB 8A B8 1C B4 1C C7 E5 5B 10 9A B0 4C
 13 CF FC 14 13 4A 7E 8A 1F 96 D3 A3 90 21 FA 5D
 C1 9E 40 89 0B 7F 3D BE E6 EE DB CB C0 BD 3C E2
 A7 74 65 5B 96 32 6B BB 17 5E DA EE 02 8A 30 79
 22 AC 16 41 0B C1 D6 39 CC 39 9E F0 E2 3A 39 B1
 67 35 C1 02 06 9E AC F6 B6 C1 CA C3 F2 7A 9A 78
 D0 E0 43 F4 86 C3 9F 1D 3C 96 A8 64 79 A9 A1 7D
 7D 54 95 ED 78 CE 59 6E 41 70 B7 46 9A 29 44 AC
 02 B8 5C D3 F9 82 53 DA 77 4F 21 00 EF DD F0 9E
 AB 7F 53 76 C2 B2 C7 CC 1F 72 1A 35 CF F9 0B D5
 7B DC FB A7 EB D4 FD FE 1A AA 36 B5 42 A8 C8 9D
 D2 01 A6 8A 69 01 CB 40 B5 92 E2 26 94 51 DE F9
 4E 61 3D E9 38 CD 5F 4D 91 A2 BD A3 BF 2A 82 18
 3C F5 99 36 2A AC 26 2E 5F 84 B1 A5 60 C9 3A 71
 26 09 8D 78 97 3F 4D E1 1A E3 43 BA FA BC BB 40
 DB 3C FC D4 AE 1D 98 3F 84 0D 47 23 40 3A 46 6C
 C0 A7 B3 A1 0B 40 2E 39 83 31 04 25 66 44 28 F5
 C4 1F 2C E8 B0 F4 B8 8D B3 CB 9F 2B F7 1F F6 B1
 5E 6C 71 C1 71 83 2E BB E7 FB EA 56 FA 68 DF 90
 BF 1E 39 79 60 A4 A1 8B C4 9B 1E A1 1E 2F 4B 1B
 30 BD D6 76 0D 40 70 25 A9 38 4A 1F C8 10 F5 B2
 76 DE DA 87 7E 9D 24 65 21 57 A0 B2 B9 72 78 55
 0E D0 32 E1 92 C6 88 8F EE C3 69 2A 68 A7 AA 08
 92 1F E3 F5 35 4F 03 28 56 B2 40 4A EA D9 AF 14
 D0 F4 56 90 AB 07 78 33 80 62 50 24 29 3D C7 29
 62 D6 C9 64 51 D7 5C 5C D1 77 7C 06 09 28 A7 74
 95 ED 2D EF FC 9D 5E 75 61 D3 F6 DD D8 C3 2C 00
 24 30 08 2F B5 97 50 24 00 9A 2F 69 EE 58 6C B7
 7D 94 C0 C5 AD 4F 66 86 71 E9 88 60 81 30 E6 1C
 EF FB CC 1F 87 88 32 F4 E5 D3 B0 88 15 6D 8A 83
 26 9D 9D 61 E4 38 DF A5 DF 35 40 ED 1A 43 0E 22
 A7 55 19 78 17 C3 8F 96 E2 6E 73 D3 AC 67 43 31
 D9 9B 76 CE 75 EF 23 14 81 91 27 8D 86 05 58 41
 BF EC 6C A1 75 83 EA B3 CD A3 DD 87 6E 2D 03 EB
 2B 35 EF F9 F8 B0 ED 0B E1 99 81 F9 56 70 1C 2C
 CE BB E3 E3 A7 C9 A0 F3 98 BC 63 58 87 0B AE 96
 34 69 AA 8A B3 6B D2 3C 2B B2 8C BD A6 E6 BF A1
 4F B3 7F 68 7D 3A D7 43 E5 64 A8 ED B3 52 BF EC
 C4 A3 7D 51 EA C2 35 E8 FA BB 2E 85 F0 4B 81 12
 A9 47 B3 71 D5 FC D1 DF C4 29 20 E4 EA 5F 02 29
 AD D1 72 42 A3 36 BC 5E D6 8E 3F 30 33 92 56 C2
 BC 54 19 DC 27 11 0D 66 CB AE DB CF B6 C4 8F B1
 29 AD 15 82 5D B2 1C 63 FD 86 C3 11 FB 19 0C 86
 CA CC 94 ED AE 63 1B D4 88 77 0F 60 41 E5 D9 1A
 8C 96 C8 56 5F F3 9E D4 F3 D9 87 66 4D 27 35 6A
 4F 5E 2A 5C F9 22 A2 87 AD 9E DE ED 94 CF 4A F0
 1B 1F 7E 8E 0B 0A AD 1B 96 13 43 AA D3 B5 8E A3
 93 65 B4 53 DF 4D 39 2C 08 44 27 41 28 CD 14 78
 A1 DE C3 F0 5C 3C 31 C8 4C 22 E8 51 ED DE 8C 4D
 61 E7 F7 16 3E 27 24 93 4C E0 86 C6 8D 7F 57 72
 21 40 1C 21 2A D3 E4 69 CC CE 1B 13 35 C6 E8 B5
 6D 57 B7 87 79 6A 58 66 2C 18 2D B2 CA 4C B2 3A
 00 9D C1 9C A1 15 CA 89 C3 64 1B 32 7F 8A E6 80
 6C 05 0C 1B 6E C6 6B 61 8E 4D 0D 20 9B 51 90 A7
 45 B0 29 48 95 10 F0 73 19 02 23 6C 6E 9F BF 39
 3E 4B 33 7C D8 A1 D7 25 3E 6A 41 9E 81 17 D7 7E
 A5 19 95 B9 91 6C A3 B8 59 FC AF 4A 23 A4 21 66
 9C 16 AE 79 EF AC 2D AB 62 FC 51 40 AB 7E 14 A0
 ED 93 16 72 F8 76 3F 16 6E 0D 2F A3 71 F1 DD 26
 22 2D 1F 57 C0 48 23 93 89 45 45 E5 9C A6 6C 92
 91 C9 04 26 62 50 0C F6 79 35 A5 E3 58 5D 3A 53
 A0 58 2E 80 34 5D 5E FA 0C 65 98 62 3E 15 6C 59
 EC D3 AA EE 0F 4B A2 3B 74 60 C1 C8 C6 4F D7 E0
 18 8D E5 03 4D 31 99 92 BE AA 2C 79 8E 47 68 2E
 4F 72 E5 BC 5B CB 71 AC 19 58 C3 03 BD 68 44 18
 9E 9B 3D D3 EE 11 87 59 85 F6 AE 56 36 81 9F CB
 75 6F 02 09 62 1B BF F3 60 DA BE 40 F1 3C 6F C7
 6A 4C D1 A3 69 78 44 27 94 8B 41 CA 15 F0 48 B2
 62 9D 15 1B 36 74 9A 1F C7 BD BA C3 30 2D 3E A8
 BF C4 94 6F 2A 7A C5 14 C6 ED 1D E7 33 6C 8C 6F
 78 51 D0 27 80 D5 7A 5A 9A AC 5A 10 21 81 24 3C
 B8 20 CA 56 82 3D 51 F0 D4 40 2C 08 CE 92 0D 20
 96 B1 56 FA C9 FF 12 09 4F 94 9F 64 77 34 00 75
 16 70 42 61 BA DF A3 49 47 47 92 B4 1D D6 58 9B
 5D BF FE 34 71 0D 9D 33 5E 8D 7B 0A 09 60 2D 52
 B3 E6 F5 D5 08 6E 36 D0 8F 0A 42 C0 24 EE 22 97
 16 2A 8C A7 98 C5 14 B9 48 0E C7 7A 3D EA 07 09
 5E B9 67 DF 88 95 2D 8E F7 66 4C 1E AC 76 A8 18
 CA 8C 36 AA 1F 3E 8D 70 A8 39 EE 01 86 1B 42 84
 92 9B 62 28 AE 3F 80 B9 AF 3A D2 97 75 2D 46 5E
 C6 13 54 1D 12 3C D0 D0 36 BB EF C0 32 54 2F 83
 34 1A F6 B2 8E C0 6A 0C D8 81 FC 4B B3 DC 64 3D
 FC 1B 06 87 F5 1D D5 5D 76 38 BA F3 B2 40 4D 90
 AF FD D2 6A C1 8F B7 D4 76 DC A1 DF CF F5 53 FA
 BE 59 52 13 67 B2 18 B3 0F AD 41 4A 81 F8 DD 70
 FF D0 03 AF C2 5A 3E E7 A0 7A 58 B4 D9 DC 3C F5
 D6 14 A1 C5 A5 8D 71 6C BF 1D 77 70 46 BB 86 09
 B3 81 F3 F0 19 DC 14 D4 19 F5 F4 78 5F 6A B1 1B
 2B 0D 17 F7 DC 94 EF 57 61 75 9A DE AA D8 15 AC
 4C 20 52 8C 95 D9 7A 5A 4C 2F 4D 8B 2F 61 2D DB
 5E 1E 3F 50 4B B2 25 84 58 43 8F 3F E1 AC B1 43
 FA DF 50 56 D0 06 2C 18 59 99 B0 A5 39 0E 20 E5
 03 5D DF 00 02 33 FB 63 58 8C FD B3 9E B0 74 1C
 BA 53 B8 8A 8E D0 2C B3 2A 6C D4 86 B9 33 87 8E
 C0 E6 DC 26 F4 A3 0E AF 81 90 DB 3E 5D F8 25 6E
 A3 F4 61 43 F5 80 0F 84 C2 73 B3 52 EF 39 9D 1B
 A5 BF 7B 70 A9 1E 96 72 C7 6B 9F 7D EB 7E 26 9C
 F3 BA 54 1E C8 B3 2D 45 1A 01 3F 95 FD D5 2D 71
 DA 3E 95 40 9D D4 2F 8B 15 8A B2 CC 4D 5B D7 A3
 57 3D E7 A0 CC 8D CF 53 57 AC 23 BE 94 80 7B 23
 41 4E 21 84 EA 9C FA 02 0D E4 E5 8E A4 37 9C FD
 FE BC AD 12 FA 6C 94 7E 53 98 30 2D 91 6E FA 7A
 FC 3E 3D 22 5C 49 C3 BD 89 37 00 4A B4 A8 86 6C
 44 F9 26 EB EE A8 B1 F9 FF 46 11 B2 E6 93 97 F5
 4F 3D 7E 81 53 06 7C 1C AE 17 3C C5 88 5E E0 8A
 C1 AC C6 D4 6B 6B 7C 01 8F 9E 89 4F 80 28 69 35
 37 F1 2B 3F 8D BB 03 37 38 A0 7A E8 2F 1B F6 BE
 17 63 48 CB 7C B5 BE D1 6A 11 41 24 96 B4 81 C1
 60 B5 F4 2B 2E 09 E0 2E 03 38 CB BC 01 A4 2E CF
 58 82 52 74 B3 B8 8C 74 5E AC 93 53 E3 8E D7 A0
 55 02 C1 73 9B 2C 06 97 8A 57 B7 18 CC 40 A9 05
 96 28 E0 21 4F 26 BB 95 57 46 90 D4 6D 51 AF 74
 50 41 A4 13 45 5B C5 4E DF A1 96 11 4E EF A5 67
 44 A1 79 E3 97 DE 5B 86 99 DA F3 E7 06 9A AE 5C
 DB D2 20 28 DC ED B6 8D A1 28 89 0F 6A 18 0D 49
 DB C9 2E 82 E7 A4 34 E1 C4 07 24 FC 27 95 F2 47
 4E 5A 81 EA 9B D1 52 4C 04 3A F9 E3 AD 6A 53 50
 E4 97 DE 07 35 51 FF 1A FF 0F 84 21 57 06 CF 45
 A3 5E D6 D9 6C F9 59 4A 16 98 94 74 05 A9 89 E4
 7F A1 44 76 98 AC EF 17 0B 62 D2 0F 50 9B 6F 27
 AF EB AD E4 10 53 2C DC 3D E9 A6 5D 77 A4 7E F6
 B7 07 CE 9A 70 19 1F 33 69 D9 F2 8A 58 DD B5 15
 88 4C D8 A4 BC 2E 82 44 92 E6 2B 4E 44 40 AB CC
 F2 DF 96 01 80 3F 33 62 26 14 D7 55 CC 57 F6 83
 E4 7B 08 BB 75 D3 B3 24 DC 31 5A 10 A8 0D 1C 55
 92 8E 0B BD FB D7 6C C3 67 8B AF 4E BF 37 4D 6E
 7D 9C E8 07 1A AD 4E 43 50 9F 55 32 C3 E3 70 B4
 EB BD E4 8F 98 23 9C C3 45 09 8E 3D 85 72 6A FF
 82 CC 1A 4B D2 8F 2D 03 9C 0E 94 87 19 D6 6F E6
 E1 5C 92 1A 4D CC 48 01 68 C0 6B 65 AB 96 CC 7A
 ED 5D 53 32 2F AF F1 D4 78 5B 56 A8 28 01 82 39
 CC 57 77 25 63 59 EA BF A7 AE 80 5C F6 60 F6 F3
 84 43 23 6F B2 8E 7E 86 4B 2A 93 20 AB 3A 35 54
 7B DC 9E 15 D5 90 C2 D7 7F 3B 1E B8 FF 58 81 F9
 3F 65 B0 A7 A3 34 87 3D 07 97 2D DA CB D7 6F A0
 15 6D 1A 2D 3C 4F AC 61 69 5F 3B E6 6C E9 E8 0C
 F8 D7 9B C7 56 FA AF 68 34 8C 49 D9 D8 4A 77 E1
 5D 3F 84 89 55 16 B1 FF D9 F0 63 0A 4F B3 82 44
 56 DF 5D 98 3A 6E 2C CB 86 FD 63 60 AD 8B 49 5A
 75 44 B6 36 0D 36 84 00 D3 8D A7 6D A5 2B 19 A8
 2B 14 D6 6D DF 27 EA F9 0F 68 5E D3 5B 30 92 9F
 CD F2 1C 70 1A 72 D9 DF 60 32 DB 06 0A 39 CF C9
 C8 9E AA FB 24 7B 4C 9E A5 A9 AD 77 21 29 92 BC
 1D 8F 1D D1 15 7D 95 88 9C 63 59 C7 9A BB 11 09
 23 8F CC 7D BE 0A 8A CC 24 E9 1F E9 40 52 64 E1
 C1 BA 01 51 C3 4B 75 D9 14 61 95 4B 8C E3 0E DD
 29 97 AD C6 AF A4 7E 28 7F 71 07 68 2C 3B 26 21
 86 F1 C1 D8 04 F4 4B 86 69 61 56 D5 7F EF 33 63
 44 A3 45 29 D3 9E 18 0B 6F 4B E1 66 E3 2D 37 55
 A1 7F 52 3D 57 D3 7A 86 28 FA 7F A8 86 C7 16 1F
 9B 90 3E 62 87 39 6E 36 D9 9B 8E C1 4C 98 CE 6A
 12 9C FE 3E 7E 38 00 1D 60 1B A5 20 56 C5 6C 82
 58 66 81 03 54 99 DA A1 A7 EF 01 B4 69 26 C6 74
 4E 56 E7 97 47 C3 05 13 A3 A5 D3 D0 F0 D5 2A 71
 D7 17 C4 67 FA 36 50 1A 04 EE 03 AD 2B 25 C9 83
 8E 02 AC A0 30 73 83 90 16 43 CD D2 3B 82 A9 81
 58 AA F6 DC AD 95 22 C2 DB 3B F4 48 A5 8A 10 65
 62 1C 0A D9 F2 40 2E 4F BE 5F AB 23 08 24 00 73
 24 FA C9 6C BF 3F D8 F9 50 D8 84 9C 72 9D 62 7F
 90 85 9E D5 2B 19 8B C8 DE C7 2A DF 6B 52 A3 94
 80 DE 2D 32 5A 18 C8 7B 9E 52 0D 7F CA E3 A6 88
 D8 45 B4 F1 55 45 DC A7 9A EC 87 27 BB EC 21 5F
 C1 F5 88 80 20 42 D6 B1 EC 8E B8 D5 CC 0B 9D 06
 B2 7D 6B 61 5E A5 00 70 5B DE 4D 79 2A 1B C6 2E
 FE 9C 9C 53 12 E4 00 D5 C8 79 12 1D 24 C7 53 06
 5D E1 E4 F2 78 B4 7B A3 CC 5E 5B A1 B6 CD 23 B8
 87 42 97 89 38 F0 DD 20 3D 37 DE 45 DB 2C FF A9
 A1 EC CE 81 FA F0 D1 07 3F 04 16 68 7F CA 4B 1B
 D4 25 4E 56 97 30 AA C7 0F E9 4D 34 93 0F 02 68
 C1 B4 8C 7A 8B 45 6F 7D F2 9C BC 5A 52 2F 4B E4
 4F 4D 49 86 41 5A 19 42 0A F2 49 0F 65 6D 00 DC
 09 DA D1 4A C7 74 33 BF 56 E1 F8 8F F1 B8 92 AB
 D2 5F E6 CC 98 32 42 1E 48 F2 9C 14 6E 9E DD EF
 42 A9 53 B8 D0 2D 26 E5 ED 64 85 01 F9 59 C6 A8
 DE BE C5 EF 93 AE CC 0F 7D 2A 34 39 A8 71 42 3E
 E4 91 1C F5 3C C6 21 1A 72 46 DC E7 40 05 3E 61
 EE 48 72 DE 99 54 F4 31 69 1D 11 7A AD 29 FF D6
 60 38 92 17 BC FB 4F 1D E6 54 BB 22 77 A6 CA B5
 25 11 0A A8 2D E0 1D DA CF 94 5B 80 E1 10 3A C6
 FC 6C 62 BF 94 32 53 C1 74 31 71 BA 28 72 38 F2
 CB 41 7A 4F EE 9F E9 C0 1D FD 62 36 09 96 2A C2
 B5 F0 A6 FF BC 8D BA B3 27 0E 7E 79 40 19 3F DE
 F5 C9 60 5B 0D 95 76 AA AF 26 8D C9 06 28 80 8B
 D1 0B A6 02 87 25 ED C3 8A C0 F3 9B AA AC E8 5D
 4E 9A 7B 94 A0 D1 4F AC 2A AE 63 28 0F C2 38 66
 0D BF B2 07 C6 C5 60 73 83 98 FA 78 13 77 E4 EB
 F2 43 F4 5D EA A7 98 11 52 91 04 CC 77 F6 EF 04
 DB 98 9C 55 5A 0F DD 13 04 A3 AD E5 A0 C5 53 EF
 F5 8D AB 52 CE 3F 1D 91 84 0A 69 B1 86 82 5D D0
 24 8E 3C A8 16 7C FC D9 8A 09 27 D4 62 12 DE 19
 F5 6B 99 D8 37 20 AA E3 EF 3B AA 41 06 E7 37 5E
 44 2C 79 DD 46 7F E9 2F B6 9D D6 3B 40 E9 3C 34
 A8 EC BB A3 17 55 86 98 C7 E2 AF 06 5E 58 99 A4
 38 AF 30 0E 3D E0 E2 C5 A8 4F B7 69 DB 14 D0 AB
 5F 4B E1 A9 72 62 56 7C 44 F2 67 26 7D 51 95 93
 25 6A F9 A9 46 EF 5A 6E 8B F3 82 92 F9 36 10 24
 E9 F7 D0 62 CB 10 00 D9 D7 C7 ED 7E 6E 2D 0C 84
 B5 40 2E B8 9E 9D 9E E6 BA BE FF 83 DF 9A 66 6B
 B9 10 2B D9 DD 90 E8 7A 5F 9D 44 98 0D B5 DE AE
 0D 44 3D 71 9B D6 23 F0 7E 37 CE 82 6C B2 0C 3B
 55 4B 34 70 80 6C C7 33 C2 E4 4B 5D C9 D6 40 5D
 49 03 1A 0D D8 9F 4B 66 1B FE 63 45 08 41 A0 F9
 9A 72 8E DF 74 0E 4C 97 A2 9C 36 1E E8 0A 0A D1
 22 65 E5 67 FF 78 36 55 75 9A 16 08 7D 2A 87 7B
 E6 56 BF A9 16 DD 31 DD 21 6A D9 33 3D 37 64 AC
 F9 23 69 05 0D B1 85 E9 92 3D 91 A3 E5 A3 19 43
 4E 22 62 7E 90 00 F5 E5 E2 45 87 9F 49 5D 06 19
 5F 19 8E 97 FE E8 F0 F5 E8 72 57 F2 D2 47 BF 02
 EE 96 12 6A 1E D4 00 34 79 AD 51 63 6B 6E 55 B2
 54 E4 E3 BD 0A EB 07 68 AF C4 31 5A 09 F6 7F EA
 46 58 86 F0 88 FD 0F B8 AE 0D 79 10 FB 29 5D 4C
 5C D9 85 2E E6 E9 26 0F DA 3D 41 7D D4 1F C6 D7
 66 6A 3A 08 D5 79 FD 73 DE DC F4 AD 91 9A B5 52
 83 93 D4 7A AE BF 6F 4C 23 79 FD C2 22 BA 74 0C
 00 2C CC 3B C6 32 12 82 BB B8 5D 83 D5 71 36 64
 66 2D 0D 11 E6 BB C1 FC E8 D3 AF 0D D2 A6 E8 EE
 E1 C2 22 3E C5 13 28 AF 18 EB 6A F1 11 C1 F2 85
 E7 41 5B 24 DC A5 A6 2E A4 CB A0 AF 8E A6 5F FD
 25 4A 0E 2C 3A 32 0D 5E 8C 0C C8 F4 AB 3F F6 BC
 E6 3A 1E B9 56 A0 54 8F 2E 20 62 63 9E 6F F9 83
 0C 53 1A 21 AD E8 BC C9 36 5F 33 92 B1 8B D7 9A
 AC 44 06 00 C7 E4 F8 BB DF 3C 82 09 06 D7 65 5F
 A3 3C 21 D3 F4 3A F9 2C D6 73 B0 AD D1 FA A2 20
 21 B4 9C 02 4E BE 90 19 B2 26 22 B8 47 9D 5C 19
 DF 4C B4 14 DF 1F F7 DF D8 F6 E2 EE 22 E3 DE 38
 15 D1 D5 8F FC 1F 7C 0B A1 F4 42 E0 88 66 71 89
 59 82 CC A7 B5 8D ED 5B 3C 4B 16 10 6F 89 C8 EA
 7F 7D C7 B9 C3 2E 01 00 AE 38 7F 81 09 E3 19 69
 CF 7D D0 C5 1D 6D 68 12 46 ED 27 D7 38 87 B6 66
 15 90 F6 37 8F 48 CC 7A 04 56 91 86 27 B8 4F 71
 DA 69 F7 37 B5 A8 D7 21 2F EB 39 A9 D7 95 09 A6
 84 C8 40 33 36 74 2F FD 19 54 14 2E 76 F3 E8 8B
 1C 65 96 65 2C 94 84 06 C7 91 71 46 81 66 D3 44
 4B 41 82 B7 24 5E 25 3F 98 1E 20 E7 9D 64 B6 61
 3D B0 ED 5E DE 43 3F EF 5E 41 B0 3D CD 98 81 EE
 64 59 35 12 A8 4C 33 FB 1F 52 46 1B B4 58 CB BB
 18 B1 2D FC D1 88 7A DB 88 91 A5 5B 6D 98 68 71
 AB EA BB B0 1A BF DE D6 C7 D0 33 22 A6 E9 31 A8
 44 B8 A2 43 A2 11 8D 7B 2F C7 5F A3 E8 57 5F D0
 97 C4 EC 81 36 7E 0D 84 E0 27 D8 C0 99 93 7B 4F
 2C EB 1B DA 71 4F 76 46 55 5B 42 E2 E2 DD A0 42
 5D 45 3D 9C C7 84 14 FD 1B CF 71 69 9C 2F 49 FA
 77 CA 58 12 0A B9 21 6C 9D EA 67 A3 55 A0 4F B9
 97 73 81 0B 7A 48 6B A5 38 45 3C 33 AD 02 70 7B
 29 0E 5D 94 3C 91 28 A0 73 2C EC 39 DD B8 98 73
 7C 3C 7D B6 A0 AE 82 61 03 7F 66 95 7E 0C DB 09
 27 31 78 FC FE 2C F7 48 16 9D 00 0B E1 37 B9 0A
 39 E8 4E 72 95 7F 93 72 18 03 B0 62 5E 43 FD 8C
 9D B8 58 64 36 B6 6B 0D 3F EF AE 60 B7 B3 39 D9
 7A 46 FE 30 7D 27 E0 9C C3 8B 67 81 8F 22 BF 14
 0B 1E 2E 27 DC 32 6B F9 2B DF 4A 89 25 15 36 2F
 54 EF 71 E3 4A 32 D8 50 26 72 0B CA 9D C8 EF 4C
 C5 67 29 B8 17 6C AD 8D DF 38 6C 54 2A AA A9 42
 E2 CA F2 42 5C 9C BA FB 0B 78 D5 A1 A5 ED 81 7E
 D9 2F E8 62 42 8F 47 9E 2B 54 A7 5E 29 20 7B C6
 17 FC 32 0B D5 70 AC 71 9D FB 1C D3 CA D5 C2 E6
 45 F3 21 75 BE A6 37 B5 C3 6E DD 10 C4 67 89 A8
 FF D9 76 51 AF 54 71 F6 FD 52 EE B4 3F 1B 0A AA
 57 EF 76 33 17 00 18 D7 3E 50 14 25 C3 0F 65 88
 A2 65 D0 C8 C7 F6 7A 8C 50 B8 BF DA 67 A6 3D FE
 0C B2 C0 E8 18 40 3D 77 0F 47 B6 78 E6 5D 19 AF
 11 DE E6 05 51 39 F1 7E 07 8B 85 A2 0F 15 9E 29
 5D DC 74 D9 30 8C 38 80 F8 2F 37 F8 1B 77 C4 EB
 55 C8 44 86 9C C5 D4 79 9F 02 C1 84 E7 0A AA 0D
 64 3C 3C 62 24 5C AE 99 DE 1E 4F 16 16 34 0D 1A
 8D F9 A2 4E 40 DA 90 C3 0B E0 D0 3A 32 00 62 8E
 0C 69 0E 0D 5E 7A 25 41 CC 14 E5 DE 3A 8A 74 E3
 C4 44 A6 9C B9 F7 89 82 F5 A1 EC 48 0E 7B 6E C0
 6E 29 E2 2C 9A 6B 57 B6 DD C9 B9 AD 3C 89 12 83
 AC A5 29 FB 3B CF 89 51 5B 19 9D 48 C7 8F E0 7C
 52 C9 17 2D D9 11 02 E0 1D EC 02 22 36 92 F7 3B
 84 28 6D D5 18 32 A3 81 DE 98 80 18 6C 33 8C 0A
 C1 39 C5 C8 FE 3D 22 2A 09 90 1A 21 31 37 C1 FA
 DF 59 D1 20 B4 1D 1D 51 8E 9C 2B 15 C8 20 B7 96
 81 59 38 D2 F0 99 73 82 1E 5E 44 A6 CC D5 A4 9F
 A0 9D DF 0C F8 65 F6 BF D2 F9 F2 42 8A 0A 7D 0C
 C2 56 09 44 A7 30 4C EE C6 7E 87 14 C6 93 91 38
 DC 33 72 7A DA B1 14 70 19 78 1C 9B AC B1 DF 9E
 13 DC AE 77 71 5D 73 19 5A CA F3 3B 47 3A FE 79
 92 E2 FA 1F F2 4C 0E 78 BD 29 3E ED 4B FE 61 0C
 EC 59 58 1B 44 52 E0 CA 8E 27 27 A6 25 26 DC 40
 2C BC 86 4C FA B3 3E 82 28 7F CF B1 C5 74 7C DE
 7C 9B C2 6F DC FC E6 06 9A 82 82 99 A0 B1 8B 61
 0D 11 1C BF FC BE 9E 5B 7D E0 05 40 45 04 AA 56
 97 B4 F9 D3 6D A9 BF 25 54 EF 5D 89 56 A9 C3 57
 3E 47 A0 3D D2 2D 3C 9D 01 19 6A C5 1D 54 40 9B
 E3 41 D0 FB DE AF 3F 10 5A A1 CA B6 F3 BE B1 25
 79 33 25 6C 2F 36 BD 08 A2 F8 2C 44 43 87 E0 EB
 FF B0 34 F5 9F 8E 3F 19 B4 42 C9 DF 9F E2 EC FE
 CA 6C B6 43 C6 87 A1 7D BC 55 9C 70 13 C3 97 FE
 C6 7B 9C D1 11 78 5B 13 7B 3F EC FF 7D C4 BA 0D
 BF 31 38 E1 18 FE 16 73 08 3E 54 FF 49 37 28 6C
 6B 5D 94 18 71 B3 C5 57 A5 85 89 19 E6 1F 0F 0B
 F3 8B 00 26 59 36 83 67 8C AB BE 1C E1 11 79 18
 D1 02 61 7C A8 7A 0C 33 7A DA 1D D6 22 5A 7D DE
 77 C6 84 C2 CC DF 31 F1 D7 4D D2 0F B3 D7 91 32
 BF 07 74 EA 32 C6 56 3C 2A 63 23 BC 24 F1 67 30
 60 3D 09 A8 F0 8E B0 41 0A B5 54 D9 FE 14 8F 29
 63 F7 04 1B 85 A0 A6 3C 49 D8 E5 DD FE 51 A9 45
 52 11 8A 9A 11 61 5E 5B 7F 90 96 05 DA 29 8E AC
 7F 3E 7A 5F 2F 26 BC 4E 11 E0 6C 5B BA 0C A0 BC
 EA B6 DA 0B EA A5 A9 41 11 84 46 F0 5A 63 40 9B
 3B D6 B1 83 78 A6 9C 02 C2 C0 7D 25 97 26 D3 8F
 B3 2A A1 9C EE F8 0B 99 54 3F 8A B9 22 FC 0D CD
 BA E0 DE 58 69 1F D0 84 43 28 F0 93 8B 79 05 A4
 A5 9F 39 1C D2 1E 15 5F DC 66 AA 4E AD 68 43 28
 19 1E FD B0 8A 2B 55 1E AB 82 4E 77 0E F0 AD 9C
 37 6A 84 07 2A 01 A2 02 94 D1 88 E1 D6 21 4C 63
 AE D4 32 F7 16 61 E6 E9 E5 9D F2 CE A9 2C 69 88
 DD AB 74 83 ED D1 BA 3D 66 EF E9 F8 25 62 4F 62
 18 90 4E 24 99 9D C7 2E FD 53 04 72 AE 0E 16 0E
 09 8A 68 7B EF 61 99 E2 DA 0D 1A F5 E7 0F 86 18
 F2 5B DE 7E F0 7F C2 09 4D 78 89 01 7B EE 4C FF
 4D BB CA 26 AF FF 4F 4B C2 27 07 4D FD 14 3A B2
 09 83 FA 3C B1 30 77 22 01 2A 5D 7D 68 07 99 C3
 B5 24 A8 49 75 C4 2F 43 AC 47 88 8D 29 AB ED 89
 AD AA BB CA 6A 1C 99 90 A6 14 7A 88 7D 54 E6 B7
 BF 05 4B E2 9A 22 0C 5C 2A 8C B0 75 CA E2 2C 07
 22 24 AD 69 03 2D 89 78 80 34 BD 85 42 43 BA 65
 09 21 43 45 0E 0A D2 13 B2 CB 5E F9 68 20 BD 2E
 B5 69 98 AC 6B 1F 8F AD 0A E1 E7 B3 65 08 C6 80
 4C 33 79 E5 B0 28 22 A8 8C 12 1E 78 7D 4A 9B 5F
 08 88 DE C4 39 72 C9 41 DD 31 E2 D2 22 A9 38 F1
 63 BF 2C 16 D6 1D 93 74 95 79 0F 95 22 D5 49 6F
 10 31 DF B5 4B F2 1F 98 51 B8 AA A1 2A 2E 1D D6
 A2 9C FC 04 56 10 D8 C5 58 CB 1B 04 7C EA 04 12
 C2 81 E8 7C 29 2A E0 B5 1E 0F 09 7C 25 43 5A 7C
 74 4F 73 F8 B8 E7 B0 73 2A 36 EC 91 01 90 75 EF
 75 DC F9 7D 2F C0 10 8C 99 C5 76 EE FA 4D 20 E5
 A8 05 C0 BE EB 77 8D 88 1B 2B A8 1E 89 13 CF 22
 E2 30 5B F1 C3 95 F1 59 84 A6 90 5B BE E4 A9 A9
 C3 A3 2A 0C 19 07 9A B0 E2 7B 5D DA CC DF DC 34
 C6 4A 12 F9 9D 91 5A 90 78 2B C2 E2 92 19 2E 8E
 E0 A9 1F 74 A1 A9 64 1A B6 A5 07 C6 44 01 42 5A
 61 7F FB EC 20 17 29 08 6B BE 59 62 97 6D 74 50
 2C F8 09 78 41 47 71 83 D7 A6 41 CD 05 2F 57 13
 B8 97 48 BD 1C 36 AA F2 5A 86 5D B1 5D B7 3D DE
 FB 39 31 DE BB 87 0E 23 58 00 FF C8 FD 89 CE 45
 45 9C 1B 25 32 D4 17 24 58 CB 37 CF 66 0C 5A 6E
 C8 21 5D E5 40 54 83 BD 2E 4C 06 26 88 1D C7 86
 0E 3B FF 4F 60 D8 14 FC 0B 08 09 C5 D0 B6 54 7D
 39 CE 3B 1A DD 42 D5 64 CA D3 CF D2 57 BF C8 D5
 68 99 8A 4A 36 B4 47 6F AE 49 67 4A C9 F6 1D 5E
 D7 50 12 6A 51 BA 49 B6 B8 78 57 A7 15 D7 5E 4F
 93 38 7A EA 41 55 B0 82 22 93 E5 86 B2 1F B5 A8
 90 E0 51 75 33 51 87 90 A9 43 19 BE 61 10 FB A0
 80 37 F9 B6 17 8C 7E EF C1 91 6F BF 3B EB 53 67
 9F 4C 87 74 DA 8F E0 0C BE 43 C4 AD D8 B9 A2 1A
 2C 1A 47 78 40 AF 73 92 52 5D B8 4F C5 1C ED D4
 1D DC 67 6B 6A 3D 72 75 A1 20 06 79 8E 58 70 36
 66 D1 FB 33 37 5A B4 78 14 76 D5 F8 71 BC 33 D6
 63 5F B5 CA 0E 08 B5 C0 ED 72 1F 8E 67 4D 9E FD
 9B 59 14 16 FA E3 F5 DE 02 0A 70 C1 25 AD 50 EF
 2A 8D 98 9D 30 D9 FC FF 4A 33 EC E9 E4 05 80 DC
 2D 8C 2E 0C 9B 07 91 7B 8E 10 50 10 03 45 27 51
 68 6B 44 12 4C 92 BB A2 2B D2 5A A1 68 F1 6C DF
 57 B1 F8 4B 02 0E 06 89 DB 5A 68 27 D7 2A 61 0B
 6D 84 34 98 5E 98 2C A0 18 D7 BA 64 9A EE 36 2F
 B3 1F C2 6C 36 F4 69 93 BC 44 7D 4E 50 18 DA CA
 50 60 FF 09 D5 B4 59 8B 2A 74 20 57 CD 46 0C 7C
 EF 4B 98 75 5E 53 3F 8F 1E F4 B2 07 D5 52 BB 80
 35 DF 98 8E 58 B7 24 D7 1C 63 C4 A5 FB 27 A8 7A
 BC 99 C6 73 B6 86 CD 25 2B 9E 3D F1 B7 E7 68 0A
 53 4B C0 49 76 58 66 8D 8D 37 98 36 CB 5E E3 BD
 DC 7D 92 33 C7 DE 1E 8C 74 13 95 B3 FD 9A 41 A2
 E1 A1 8C A8 A2 D4 17 39 21 46 0D 29 DE 2B FF 2D
 88 08 CD AF 40 D6 84 15 5B 02 2B 19 DA 89 AB A3
 66 1B EB 6B F7 F3 42 DC 0A 5A 03 1B E6 C3 B9 46
 B9 88 73 C1 26 96 74 5B 37 57 91 95 FB 6D 0C 8B
 12 50 30 F0 B0 CB 62 F3 67 33 63 B0 65 48 D7 08
 BE 83 77 07 41 5E BA C5 5A CA 5D C9 BF 04 1F 0F
 05 22 DF 69 B4 02 8F 69 E6 AF C9 A1 3B 5C DC 0F
 A1 47 46 41 25 39 38 57 AA 41 08 F8 41 51 40 AC
 3B D6 F0 08 7A F3 A2 ED 65 EC 8D 0D 77 CB 99 C0
 09 B4 61 D3 F0 1A 9E F2 E3 58 76 08 6E 19 8F 42
 B8 56 6E 66 D8 85 3D C7 C8 1B 7E 10 4F DB 98 E3
 77 58 34 C8 09 F5 55 3B F4 A1 D2 95 6A 0B F5 05
 59 42 1C A1 B1 E5 A1 CE B1 C1 FA D7 0A EC 17 78
 0B DA 5B A8 1F F1 4E 4E D8 26 BA 8A 01 86 D3 00
 87 D0 8B 11 26 25 39 76 30 5C EC 7E 65 E4 DE 3B
 14 13 3A 9E 3D 42 DE 59 52 68 2F B1 C2 BD A4 2A
 CD D2 56 70 9C 97 70 53 8F 13 A6 44 6B 91 12 96
 9E 81 B4 50 1B 6E 75 E2 49 6A C1 D3 0D DA A5 CC
 8F 88 11 16 1C 04 63 97 C1 5D 2D 0E F8 AA E3 92
 E9 2F 55 A1 35 A8 E4 C1 43 EC 58 08 1E F6 30 BA
 97 04 1B B9 D0 8B 6E F6 3A C4 34 8A A8 D7 79 55
 00 0F 89 0F 98 3D 9B CD 32 91 44 1F BD 04 25 CB
 77 5C 79 5E 0C B9 69 0A 2F 54 BC 01 12 88 91 E0
 37 86 54 30 EC B4 05 B2 B6 90 AA 3D 04 C9 60 35
 6F 7F 7D ED 94 3B 39 F2 3F CB B8 B4 0B AE CB 20
 75 79 CB DE 1A 42 8F 4F B5 28 65 35 21 40 93 54
 C5 DB 4F 61 3D 50 A3 3E 3E 40 A5 5D B0 C4 2F 23
 A8 CF 2D 40 EE C7 1B 91 FF A0 F3 5D 3D F0 04 BE
 73 BE 19 17 AA BF 03 76 2B CD 76 93 26 E9 B0 A3
 84 EB 50 26 73 A7 D7 58 2E 4B 3C 1E 23 0B 68 19
 F5 DB 40 0D E8 67 B2 3F 40 12 C8 CC EC 12 0B 94
 1F FA 88 9F FA 71 02 FC 37 CB CC D8 D2 C0 C7 69
 14 07 74 8E 71 6E 1B 57 0C 21 79 2D 59 7D CC FA
 91 94 60 45 D4 45 2A 0E 00 FB B7 E1 9F 40 49 64
 10 5D BE 04 EC F2 4F 37 70 CE FD 8C 5B 1E 78 1E
 03 62 EC C6 1F AB 71 21 3F 84 1F 83 E5 1F 9B D5
 8E 9D 8F A3 2A 4F B6 A4 C9 F2 48 81 72 91 A9 F0
 83 F1 6D 52 FD 63 41 3D 82 5D BD 4B 40 5C 29 82
 D7 40 9D 87 EE DB 14 7C 61 2C 7C 8A 5F FE 37 F5
 52 4A A2 AD 87 A8 22 08 12 03 29 3E 66 47 83 5F
 7C 29 CC B7 0A 83 9B 55 39 F8 A5 19 E9 93 07 82
 5C 2D 15 30 D6 AA F9 91 61 72 50 43 A1 68 62 B0
 59 EE 0D 94 3E D3 9A 2C 77 F1 DB E2 2F B7 1E 72
 56 03 15 4D 27 31 3C 28 6F DC 73 72 C9 1F 29 E2
 C6 6E 4C A3 A7 7C 46 B0 64 B7 0C EC E7 9B C5 6E
 6A F0 4F 59 3A F8 40 2E 33 3D 0F 4A 24 1C 71 81
 2B 19 E8 6D EB C1 43 36 D6 AF BF C4 40 2B 04 07
 27 33 E9 3D 7F B1 AE C6 EC C7 BE A8 A2 58 AC A6
 51 73 AC 50 1E B0 D6 DA 5A 73 F4 41 04 37 C5 6B
 FD ED 8F 78 93 CF 38 3E E0 94 E8 DD 4C C4 61 FA
 21 F1 1D 70 7C 6C C8 BC 70 B7 C2 8C 2F 9C 8B 9E
 AF 7D F7 64 05 D8 CB BA E9 4B EC D7 0A F0 38 05
 61 1D 2F 15 55 20 75 82 7A 26 4F C2 39 A2 13 0C
 61 D2 41 CF 8D 0E 73 62 5A 1E F6 4C F2 A8 E2 EE
 71 E2 36 70 95 09 38 86 D1 9F F8 0F 55 AF F1 18
 FA 4D B9 8E 3E A4 77 92 A1 C8 E8 45 44 10 AB 17
 0B D9 C4 FA 5C EF 1F 25 55 C6 E7 06 90 05 7F 61
 B7 4E 5E 67 D0 DE DA 22 8F 51 B5 73 09 9A 4F 5A
 EE A7 42 54 45 8F B0 F5 9F 46 3B EF 70 80 3D 60
 2A C9 47 4F 8E E2 F7 14 A2 BA 22 1B 5A 9D 91 65
 DA 4D C2 31 E6 6D 77 75 F7 E1 5D FC AF 6D BA 73
 D7 E1 D0 2F 80 34 14 77 59 78 54 1E 4D E0 96 CB
 DB 02 9D F7 5A 3C D9 D9 66 9D B0 8C CB 15 76 17
 2F CA 92 F2 A1 3B 23 5F 68 B4 55 F1 20 41 65 66
 4F 8B 74 66 46 45 E8 D6 C7 CF DB F2 84 69 60 61
 FB 9B 16 48 B8 B7 A9 59 3A 42 47 E0 8D BC E5 7F
 FE 04 D3 51 30 0C 6B 46 30 0E A2 91 44 3C 74 2A
 4F F0 FE 30 19 D1 9C A6 45 73 54 6E 4D AB E7 E8
 6B 5A 4E 69 CC 74 1A 90 2D 3F 16 5D BE A2 03 D8
 6C A7 A1 86 01 9C 81 57 D3 65 67 08 6B 03 47 78
 2D 65 17 B9 B4 7D 33 D3 0E CC 85 01 8B 17 77 E8
 CD B1 32 CC B1 84 E7 BB 78 42 93 C5 69 3C 73 A0
 65 98 B2 29 2A 8C 18 B2 86 D1 F5 04 BE 99 5B 0D
 9E C1 64 94 99 58 0B CB B2 0B 62 78 40 71 10 10
 CF 23 F7 84 94 7F 49 3C 92 F5 5A 9F 47 AF CF DF
 00 95 8E B0 EB 6F AF 2C 3C 32 9B 9C 8F 23 36 22
 47 A8 B8 B7 A4 68 CD 72 58 54 91 27 7A 2D 2C 0B
 11 C6 FE 16 02 63 E4 39 4A 88 57 BF 75 BD 17 03
 A4 77 B5 28 D8 41 3C 1A D3 6F E7 C0 4B 22 60 6F
 3F EA A0 CF DD 26 3E 11 77 26 C3 22 1A 9F F1 64
 26 99 09 33 3F AD 87 E1 0D E6 EE 13 06 1B 90 D9
 F1 0B CD 16 C6 A7 3B 65 CF 3D 42 65 2F 77 E7 AB
 FC 32 AE F7 33 2E 44 4C 58 34 C4 B6 4D CD 59 ED
 1A A9 3F D5 E4 65 CC 46 03 28 E9 98 D5 70 8F 79
 37 03 E2 58 2B C3 6D 12 E0 6B 7A E0 46 10 93 9D
 C5 AB BF 0D 41 94 C5 CC 0E 90 85 7F 8D 69 63 26
 D9 B9 12 90 01 62 01 8D A7 9A 63 68 E6 74 AE 02
 D7 F0 0C 20 10 A5 22 95 B2 5A 00 44 DB AA 20 0D
 E0 A7 B1 31 81 53 A3 EE FD 9A B2 84 60 D9 22 87
 B3 71 63 42 BB 3F 0C 60 BC CA CF 1B 4B B0 A0 D7
 BC 2A 43 46 20 DD A5 41 3D 4F D5 06 8E 26 AD 5F
 77 5D 57 7F BD F1 C0 04 43 2A 49 E7 60 20 10 16
 96 3B B3 A6 C0 87 11 4A D7 EC DE 32 02 3C 38 31
 E9 60 60 AD 97 55 29 7D 58 EA 38 0D C5 55 39 A5
 4B E3 A7 61 6F C9 E9 D4 E2 7F 63 5C EC 85 C3 0F
 A9 F1 A9 B9 C7 E4 30 1E 55 7D 18 EB 3D BE 0E 7A
 3E 94 30 48 21 3E F4 7D D6 9C 03 A3 DC AF C8 7C
 CE C2 8A D9 AE ED F8 AE 6A EE 9E A5 92 EE 6E 41
 CE 17 E5 B5 66 37 A7 F0 7A 04 E0 2F C4 24 90 6F
 61 3E EC AF 7C A0 3B 70 16 BF B5 9F 7F 15 85 A4
 9A 99 E8 8D 01 A6 C7 F9 E4 B5 A2 7A 7C 05 96 11
 A0 AC EE 9B 05 7D 0F 03 5D 0B D2 89 F8 08 C5 CA
 DD 2F 9F 63 E5 4E C2 F6 8F D9 06 20 FE 0E 40 8E
 F2 C1 67 F7 3B C5 E3 89 20 FB 51 BB 34 50 1F 36
 99 D8 EA 06 5C A0 1D 46 0E 3A 48 1A 80 7F 1D 8F
 96 B2 05 8D 6F 87 B1 97 5D EC 90 44 0C 61 A1 CA
 D4 DA 0B 1F 5A F0 11 53 1E 72 3D 07 FD D8 6F 66
 9B 9F 30 8C 47 E8 B7 04 DC 30 F7 68 F4 EB 68 E3
 FF C1 28 C9 93 A4 19 E8 B0 0E B0 8D 04 82 3E 0D
 0F 94 C2 0C 28 FF 94 6D 91 AA 80 01 A8 2D 70 50
 12 90 6A FD E2 EC 5E 9C 35 3E F0 F8 13 87 82 68
 54 02 84 A4 C8 2E 4E 82 FD FC A1 A3 29 65 67 88
 3E 27 2D 11 09 76 BF AC D6 5B C5 1A 7F BD 68 37
 F4 A0 75 31 4C 58 9D 53 29 C2 AF CC E5 75 95 6C
 97 2F 25 B3 69 3C 2B 36 A8 EB 0C AD 15 1B 1E F8
 95 86 02 43 A7 12 4A 52 49 5A 52 11 A0 23 9C 4D
 31 4C 0B 97 09 BA 89 E6 E3 FA 57 69 DD DE 6A 78
 95 DE B9 79 24 ED D6 32 DC 52 D4 E1 67 02 2E 63
 A1 51 25 72 EF 07 B6 17 78 46 18 28 C4 F5 EC 68
 D8 78 8F DA E5 CE F8 A9 CC BE 89 3E D0 FA D8 95
 A6 C2 CB BB 1B 09 55 3B CE F6 09 F9 C4 2D 7E A6
 82 EF B0 F3 35 88 95 FD 63 9A E2 78 9B CC 85 DE
 39 B5 D0 5C 4D CB 00 0D 8F 8D CC AC A4 F9 01 3C
 91 FC 17 49 BD 42 8D 62 6F 3D 99 B0 B4 BB A2 64
 44 94 E5 41 49 FD EA C7 74 05 4C 40 CF BE AB 60
 D7 CA 34 25 D6 62 BA C6 FA C1 44 E1 5C 83 A0 D6
 06 B0 D4 F4 25 AE 5A 29 35 B3 3E C5 1E 3F 67 3C
 C7 83 46 A3 07 D6 94 CF 8D E1 C1 C6 92 17 A6 86
 A5 35 AF CB A1 3C EE 2A 42 D9 C3 81 09 13 64 57
 33 DD 68 F1 1E FB 83 2A 31 9B AF DC EC 0A 39 22
 2E 2E 0F B2 98 5A 63 E4 BA 6E A6 89 5E 3F E4 36
 70 2D A8 2E C5 75 88 5F 12 39 14 FE BF 91 A5 F7
 EF 14 AA 92 8F 7C 2F 08 3C FD BB 4D 1A 72 55 C6
 78 BA 0B AA B0 EB 0C 99 E5 26 62 B5 1C 7D A6 96
 63 5D C6 1F BF EC 07 DF 39 1A DD 74 6F E0 51 2A
 77 0A 0E B4 2F 1A AB 19 1B 51 78 BD 42 6B 5A 0B
 78 C6 CD 2C ED 5D 9D F9 B8 F1 3E 6D 39 9C D8 C8
 67 9E A5 0D 7E 1F 13 42 29 C5 B4 8E 36 DA F3 59
 A6 3D 1A 8D 41 8E 5C 8A 61 9A 7C C4 77 85 B0 E5
 FF DE E5 C3 97 D3 8D A6 AF 58 1D 26 DF 6E 83 61
 69 A4 7A AA 02 96 75 FB CE 02 E5 A9 E9 E9 CC E2
 BE F3 E7 28 E0 32 26 E8 3C A9 DD 70 0B 41 FC 15
 14 98 54 F0 59 FE 49 19 03 64 C2 B9 8E BB AE 07
 28 D5 78 D3 BB 28 3B 71 79 AD 8A 7D 39 D8 D6 EB
 EB 32 C8 5B 08 ED 48 1F B3 52 DF 5C F2 85 9D DA
 9D 4C B7 FD D2 C9 72 58 1D D9 F4 F0 CA 4D 05 BA
 C2 7D B8 32 6D 1A 37 98 03 55 0A C0 BC DF A3 BB
 C5 EB 1D 8F 9F 85 F9 B4 4C 1E 2E 29 61 9E 54 41
 0F AE BC 6C E7 64 28 64 C4 8B FF 87 F1 1E E1 11
 1C CC C4 A9 1F 31 53 D9 FA F0 AD ED EE 07 F6 E0
 DD 44 4E 46 6A 1A 6D 67 A1 1D 74 0A 02 9E 2B 97
 4D 66 85 E3 FF 06 7F AA ED 24 18 77 E7 92 C1 71
 CB E6 13 CE 0E 56 65 C5 D1 CE 7F 02 63 0E A4 82
 26 FB 86 DE FD 47 11 F9 38 7D CF 6C 55 C0 91 58
 93 48 3E B7 E9 23 40 45 BE 19 98 28 DD 71 06 14
 D7 C8 67 47 58 47 74 72 08 FA DA 6A 49 C1 DA 91
 5A 47 28 8D 46 D6 F4 5E 87 1F 5D 19 E6 F7 FC D4
 C6 C0 A2 D4 3C 23 F7 F5 B8 75 3F CB 4E 33 AA 6C
 C9 E9 A3 F3 0A 27 CD 6E EE 2D EA B2 84 47 52 2E
 B3 5D EC 2D DC D6 A2 BC F7 F3 5D 1A 86 8C 2E 64
 3E 85 C5 20 8E 7C 82 0E 75 36 FC 78 4B F4 25 60
 AA 40 D0 BD CF A9 57 8D 93 5C 11 AA 25 5F D7 98
 48 D4 A0 73 B9 BE CB 44 23 18 7C 4D 8C 37 4B 53
 CD F6 07 A5 3F DC 3D 17 EF 6D 80 DF F6 95 D6 9A
 AA 84 A8 A6 AD BC 6E FB E1 DC 5C 6E 28 84 8D 71
 0D D5 5B 9D 19 53 47 4F 83 A4 FA 44 60 35 9B 2A
 04 1D 59 AE B7 BF 80 66 D3 B2 E7 96 82 28 F3 B3
 DE 05 EF 9B 19 2A 75 DB 82 6E 56 07 2A 88 C1 30
 41 B1 7D 7A 6E B9 80 1C EC EB 11 BE 16 5C ED 09
 8F AB B2 77 CF 83 32 46 C5 B0 8D 75 9F F1 2B D1
 59 42 BE 29 30 EF 72 8E 12 84 FE 1F 0B DE 82 95
 1F 1D A4 36 29 1B F1 E9 62 81 7F 0D BC 52 5F DC
 03 84 F3 1B AA EA C2 93 6B 7B FE DB 0C A8 DF 3E
 E9 E1 F8 A8 C1 7B 4E 7C 75 ED 3F 47 76 74 91 3B
 37 10 78 62 AC B5 EA B9 9A D7 D6 57 1E 63 28 3A
 BC AD 80 14 27 EA 22 63 79 4B 20 62 47 CD 53 57
 5F 9B 73 B1 FD BC E5 5B 5E EF 32 1F 87 C2 22 EB
 63 F8 91 E6 0B 59 85 42 61 9B 8E 61 ED 7A 81 C7
 1C 4C 24 F1 23 FE 8F F4 09 D4 01 AF 15 DF 22 AB
 1D 5C F8 31 41 4C 66 C4 20 3C 4D 09 12 3F 9C A9
 A3 D0 3F 0B AA 2F DF A4 A6 C4 B0 74 91 4B F0 D6
 2E 4A 53 A2 7E 37 F2 06 B6 DE 70 36 00 46 83 A7
 00 BF 92 6F A5 E3 5E AB 63 72 6F 28 9D DA 95 8D
 20 56 7E 66 C1 9D 26 5A 50 B9 85 27 D7 E5 9A 90
 52 61 80 9C 35 5C 0A 78 6E 77 5F B5 BD B7 D6 F4
 26 9A 0E 05 41 42 5C 67 C0 D5 CB 4E 52 4C A9 BF
 E5 CA A3 B9 19 03 6C 4C 36 9B 80 88 43 60 08 A3
 4F 41 56 67 11 41 2E B6 DD 45 E3 A7 3A D2 F0 25
 6A E3 77 EB 33 5C ED 5C 16 84 41 55 A3 C7 FD 0A
 D5 F1 FA FF 29 A9 5B DD E2 9B 9C 78 75 46 23 8E
 9D 7C D9 B7 44 19 18 3F 42 CC 67 EB A0 6F 78 A5
 C7 F5 3D B7 5E BD 96 8D 4E 96 C1 B4 F8 E0 EE 20
 39 B4 70 3D 32 5E 65 0C E6 93 AD D6 05 7E E2 CB
 4A 25 B8 D2 9D 85 34 4E 1F E8 94 FE ED E7 D0 A4
 73 92 32 ED 5C C7 FA EB 78 24 C8 B2 A5 4D BE 80
 77 97 10 95 F3 78 D8 8F 5A 08 B9 46 57 A1 BD 52
 0D 8E FC 6C B9 08 3E 93 59 BD 79 F2 2A BA E5 48
 3A FD AE CC 6B 54 B0 59 71 D2 F2 53 F7 A7 F1 30
 5F 1C 7B B0 A9 E4 8B EF FF 63 40 87 B0 15 3B E5
 81 53 B6 E2 97 D9 5D AA B8 1E 30 38 CD 9D 17 E9
 04 76 4B D2 AA D4 2F FE 3E 9A F7 BD CB 13 6C 87
 D1 59 CC B3 82 E5 B2 69 B7 67 A2 71 6C 0E D2 4F
 9E 2E DE EB AD B7 00 4F C2 DA 46 DE 94 60 74 27
 12 EA 17 54 6B C1 B3 CA 0F 66 AE 5C DE 20 FB 57
 D5 A1 F4 C5 40 CD 59 DF 73 08 EE 58 E1 B2 82 56
 E0 0C C3 A1 4A 29 1B 73 F3 02 52 D0 B9 F5 5B 26
 D7 6F D2 88 FB D2 D8 EC 54 59 3E 64 25 0D 69 B6
 9B 3D D2 23 76 24 12 43 3A 27 5F 81 08 55 49 D8
 8F 42 51 AD EC 7A A5 F0 97 F1 94 B7 26 2B 5F 6B
 1F F3 39 52 79 80 3D AC 30 1F 8E 58 5B 00 E5 00
 CD AC 1E 39 95 2B 3C 57 6F 96 32 AC 1A 89 6C 29
 A6 22 04 E9 21 2B 71 30 AB 2C F7 65 14 C6 07 6F
 98 3B CF 81 77 8B E2 DE 6A 62 34 2A BB 50 08 0B
 C7 1E 7E 26 F0 DB D8 CD 87 97 45 9F 6E 7A 02 F7
 FC 5F 29 88 0C 06 A2 45 6A 65 08 89 13 9B AD 92
 7E 75 BE E4 04 B6 17 B3 0D FB 2A 94 5F 0B 50 17
 95 CC 65 72 8B 19 E6 BD 90 92 ED 11 CE B0 6F 8D
 40 BA 0D 1E 7C 69 48 9B EE 30 28 8A 8C 2A 52 DE
 22 96 D0 F4 0A 8E 2E F8 92 D9 02 4C 83 19 A7 C0
 99 62 32 47 BF 9F 00 B2 F2 F8 D1 0D 29 93 97 88
 4C 7D 59 F7 13 BC 85 06 9E D3 34 1C B8 BC ED 7A
 2D C2 AE 8C 78 56 CC 8F 77 4F 4E 2B B5 CF 22 31
 17 81 3B D7 6A 32 29 6E F0 06 04 50 67 D9 23 07
 BB 66 D3 21 D8 D0 73 6C 28 7C 33 3B 2B BE 10 94
 DE 81 95 17 62 24 44 2F F6 1C E6 5F B4 85 CD 89
 1E 49 FE 2D A7 89 FA 3C 6D 07 B7 AD 85 FE 3A 54
 DE 34 71 A5 DC 75 D5 1B A0 59 3B 8F 16 D5 0E 4A
 3A E7 40 E1 59 2A 87 D1 E6 8A C6 9C 05 17 E2 CA
 2B 7A 2C 0C 13 CC 4B 34 08 5F 95 30 C6 0A 0B BD
 86 04 E6 77 78 A9 97 43 20 24 C5 5C 3C AC DD A8
 2A 5A 47 0E C5 12 E0 F5 F4 ED 5B CF 6F DC 86 24
 F2 06 17 12 55 91 D0 C8 88 CC 49 90 7F EA ED 34
 AC FD 48 FC EF 97 24 8E D9 D7 81 A2 48 55 D7 AA
 CC DF 75 36 5A A4 2D 5E 7A 7F E8 58 26 06 9B B3
 E3 52 D3 E3 C5 42 DD 43 F8 B0 F3 FC 16 BE 8F 7E
 97 7A 6C 2B BC 61 8D 4F 61 38 58 77 E6 99 F7 BF
 67 04 3A 3A E3 50 E7 36 00 F7 F5 CA 38 66 2A CB
 2E 2E F1 9E AF 57 35 22 AA 8B 96 14 D7 B8 92 75
 53 C2 10 02 B8 E6 8F 74 31 A3 20 0E 08 E2 A5 F2
 68 D7 44 54 4E 7F 3A 18 16 66 CF 82 7B 9A C0 54
 11 F9 39 2F E0 EB E5 6D 93 BA F9 51 60 89 4D 1A
 83 47 20 D2 BD BE 64 06 B7 11 A1 4C B2 73 CD 77
 49 6B 08 C3 62 B7 A3 A5 9D 89 C5 32 2A 74 02 98
 D4 1E 64 DA 72 7F 8A 31 B6 2B 12 E1 7E 78 D7 15
 D4 09 29 F6 44 63 34 A1 F9 E5 4D FD E4 8C C4 F4
 4E 1F E4 9A 50 10 C3 BF DD 1A 09 B4 6C 92 80 E6
 C6 F1 61 EA DF 26 6B D1 3B 4C 6A DC 0D A7 0D 72
 D7 FC EA 12 E4 EB 7C 46 6A 6B 36 4C D0 BC B3 4A
 39 04 0C 17 6F 2D 75 BE 7A 1F 5D 6F 56 91 71 EC
 A1 A3 B3 55 CD C5 CA 18 01 22 33 0A E7 3E B5 EF
 A1 B8 DE 05 80 11 CA AB 8D B7 90 69 4E 0E DC CE
 5A AB EA FE 4B 54 B8 4D 45 96 20 0D 13 C5 0A AE
 B6 71 4C 4B 4C DD 61 9B C4 02 56 A3 7F 01 C2 E0
 6C D5 42 86 6B 15 98 AD 08 53 2B 23 9C 06 39 F0
 0C 77 A9 F0 2E 24 E6 4B D0 30 78 6C 06 83 54 48
 68 C6 8C CE 7D CC 96 0C 9C EE D8 98 E9 B5 BC 10
 07 97 80 CA DB AB 60 E7 E1 01 14 0A AD 34 98 9F
 11 88 5F 9E 2A 76 64 2A 59 89 97 85 AF 57 18 2B
 E1 15 6D B9 E2 9F 1A 87 02 5F 99 BC 0F F8 1A FA
 69 80 BE 54 53 93 E9 4B C5 42 0F 4A B9 6B 92 A1
 72 68 01 48 5D 43 61 25 B9 9D CC 00 D9 7E 87 7C
 A6 A1 D1 BB E3 32 4E 9C 47 0B C4 07 8C 73 B9 B3
 14 44 3B C7 DC 89 29 A6 94 9B A3 B0 D5 12 53 DA
 C8 A8 73 CA 0A C0 1A EF 5F D6 0F A5 D8 0D D5 BC
 87 6D 2F 1D E4 4D D0 57 66 4B B4 28 02 31 78 B6
 89 B2 97 9E 74 78 12 96 6E 34 B0 E6 1C 90 6B 2B
 22 3B 24 E7 82 26 90 71 A4 D7 F2 E7 FF 8B 2F DE
 CC 43 13 47 FE DA EE EA 77 7C CD 0A 26 9F 15 CA
 E9 C2 D7 1C 5F 61 A5 0E 38 45 66 A2 D1 51 5D 5B
 1D B8 D6 C1 1C 69 03 93 C1 C5 E0 C3 B8 6B AA 19
 17 94 D3 73 34 B6 B1 1C 0A E5 AB 13 81 DB D2 35
 47 EA EA AA 22 3F B1 F3 54 B6 D8 95 BC 2B 27 0A
 55 F9 71 3A 8A 61 73 0C 8C E3 9A C9 B8 54 A3 0C
 18 B7 B4 1A 34 00 60 8B 4F 43 BC 9D 42 AE 04 CC
 3B 49 AE 16 DC 94 69 CD 0A E6 CE 92 F8 8B 6C E6
 7A 81 0F 31 3B AB 80 E4 84 57 31 6C 99 05 EC C4
 C3 0D BD 1C F7 95 9D 73 B8 3E 46 8F A2 42 2C FC
 1F 16 C6 FF 2E 34 92 DE 1E 75 7A 63 6A 7C 24 40
 88 0C BC A3 C8 3B 8C 39 2E 9B 7E 54 D2 A3 11 12
 E2 9C C2 E3 8C 55 65 15 40 FD 9B 55 47 51 42 90
 D4 5D 40 A5 F4 30 57 EB 2E 69 A2 57 6C BC 7E 68
 15 57 59 7A 45 6D 13 38 61 4C A4 A3 1D 87 9E 11
 DE 74 39 6B 2B 49 B1 2C C7 F7 93 A5 B6 6B B6 58
 DB 2B 62 97 90 C7 F0 FB F0 2B 1A 2C 1C 8E 8A BD
 29 26 EF D0 82 BD D2 50 62 0F 90 66 1A 69 D9 8E
 00 F3 AF 11 F2 37 64 79 91 0C 15 B5 7E FA 51 4D
 64 66 42 77 0E FA D1 D7 5E D1 05 46 75 DB E2 C4
 E8 A5 3E 81 A1 FC 71 1B A6 37 70 14 A8 75 EC 87
 36 AC 2A 65 B7 63 8E 5F 81 42 D9 A6 34 AE E7 B2
 58 54 CD 49 BF 16 00 F8 E9 90 71 C6 DA 77 F4 84
 55 F6 76 73 AB 24 10 73 FA E2 28 8F FE E3 90 1B
 91 CB 78 74 49 16 91 76 A7 88 D2 E8 81 2C 01 D2
 E2 38 EF 10 1E 4B 69 B4 35 1E 01 CC 1C 51 6E DE
 70 13 8A FD 5D F0 C1 D6 9B 14 F3 42 9D F7 CA F2
 2A 73 96 8B 71 B9 F9 10 F7 40 F3 E0 D4 28 36 6A
 09 D0 E2 B0 93 D1 B2 F9 46 7B 94 25 E3 9D 5A EF
 EF 80 DD 1D 43 48 22 1E 4C F3 5D 5F 6F 5A F3 FB
 F3 23 D2 22 4C 9C 86 D7 EC E5 2B 48 A5 72 5D 07
 E4 0D F1 F2 83 66 54 71 03 40 6A EC C7 64 6E 1C
 82 D5 D9 A4 26 7B 40 B8 21 AA 86 63 A7 C7 44 62
 62 A6 5F EE 10 95 97 14 5D 3E 64 67 4B 78 0E BE
 6A 61 9E F1 3A 8D BA 81 09 11 F8 2C 36 08 DB B1
 18 B5 A6 C7 D7 9D 11 92 EE 83 9D BB 97 0E 8B 8C
 C2 58 18 73 5B DC F1 F2 EC 78 38 9F F8 93 A9 96
 9A 92 3C 72 03 B6 66 4C 2D A3 03 70 40 4A E4 9A
 01 D7 D2 7F 8B 24 85 99 CE E2 AD 7B CB FC 77 9C
 23 F8 9D EA 31 97 D7 47 04 15 38 2F 83 A0 65 2B
 57 B1 9A 66 14 96 11 2E B8 01 1A 36 EF 10 91 51
 82 30 BB C0 58 BD 19 EF 61 75 DA 4B AE 30 15 83
 80 08 D7 84 9A 0A 0B 45 28 99 56 4B DC A6 E5 91
 BC AB 26 24 62 93 4E 6A C8 A8 9A 58 1B 28 3B CF
 E8 6C DC 2D 2D 6C 9D D4 9E 85 B4 CE 14 8D 6A 10
 9B 65 04 72 D7 82 AA 6F FC 7A 2E DA AA 72 82 DC
 22 E6 BF 04 F8 5F 1C F8 9E 34 1C 69 EE 63 94 FB
 4D F5 95 BE 75 1B D8 3D 04 79 6E CE 93 03 32 F2
 B2 D0 A9 D2 5F C7 9A 69 ED 26 EC 42 EF EA 38 B9
 79 BC 22 80 5D E0 01 CF C1 67 19 DD AD E4 4A F3
 9F 87 A5 8B AF E0 D5 D9 68 84 89 8C 0A 78 73 69
 7D 48 EB FD FC 85 16 FB 36 8A 3A 8C 9F 63 AF C3
 86 AF B4 10 2B 7C 3A 2F 30 AC 7A D2 32 F2 A5 2F
 CB 89 B1 C7 16 2D 0F 73 95 90 B8 DC 60 5F 0E 32
 04 9E 8F DF FC ED 5E C9 DF 94 C1 04 DC 85 23 C1
 E8 B3 F2 D6 92 AE 10 DE 8B 32 5E A7 CD FD 6F 08
 8A 21 4E D8 21 92 F8 01 E5 05 B1 4F A0 FA 70 76
 BD 6C 9F 87 C7 D0 F9 80 18 92 83 05 B3 F9 00 EA
 A2 AC 97 74 3E CE C3 C2 3D 77 81 19 3D 19 56 03
 20 10 0F 30 91 9E 11 68 8C 01 F3 42 B9 6D 72 D5
 80 00 6A 5D 8D AF CD 9F 6B 01 A4 E4 88 DD CE 32
 2A BB 66 A8 A1 42 A3 26 C0 83 BD EC 20 76 2F FF
 04 97 7C 6E 4E 7B C9 28 69 0B E3 FB 8F F5 AA CB
 BA D3 09 AD B9 8F 85 1C FA A8 3E 6C 31 6B 6F DA
 D3 B0 AB 91 A4 1A BF D8 8A F1 50 C0 8C 3C E2 83
 CA 1B 0B 7A E0 2A D6 1D 6C 7C 44 D3 FC AA 49 12
 FF 30 67 45 44 26 8B 4B F5 34 24 64 8E 75 9F BF
 37 4F 61 89 D3 47 39 8D 92 EF 41 44 1C 3A EA BD
 21 A6 4B 01 1D 20 F5 7F 6E 69 C6 0F B8 5E BA EB
 44 55 95 50 30 CF DB F8 35 70 7A E5 51 D7 A0 18
 1F 9D 82 B2 BF 53 1E 51 43 BE E5 67 12 A7 B7 8B
 7E D5 9C E8 18 E6 DB 0C A8 C9 25 7D 5C A4 FC 23
 39 F5 36 1E 66 32 DB 73 00 A8 31 4C EB 8E 8B FC
 31 2A F1 D4 6E 5A 98 F9 D8 8F F0 B8 4B 44 67 94
 4D 3C F0 AB 44 FC 95 7E E6 5F B4 5D D4 F3 64 3C
 C6 E4 36 B8 AB 9A 2C 51 20 81 EA 6E 00 D6 EB B0
 E3 30 90 27 1C 10 2A 28 16 5A D2 9D 24 F4 9A 96
 01 4E ED ED 72 81 06 2B 70 D6 AA 30 FC 88 8D A0
 8F DE A6 5C 5A A0 B6 78 D0 78 7A D5 1B ED 5B 9F
 0F 91 F0 EE DE 8C 52 7D E8 2D AE BC AB C7 7F EE
 0C 7D DF 36 46 40 9C B8 74 8A DD 11 16 7B 6F 0C
 C7 73 DB F9 27 31 83 1D 20 D4 0C 5F 8C 1E A7 2F
 60 54 96 F5 9D D7 95 E0 C2 AC 08 A9 69 81 1D 36
 BF 14 82 02 2E AF FD 3B DC 6D 0C 13 ED CA B6 E1
 91 4E 86 7F 0C 43 C7 E7 1A CA 69 62 71 94 92 27
 DD 79 AD 6A 9F 68 21 FD 73 29 73 8C 57 CE 5F 6A
 26 D7 F5 47 C2 0E 1C 16 DC 6C FF 89 55 C1 20 1A
 6A 55 AB 91 4B 4B 3C 81 86 6E E0 16 01 55 38 E2
 07 FE 25 0F AE 2E A3 E9 E6 1D 26 46 A3 CF 4C 16
 54 F4 C6 FE C7 8A 1C 1A CB 3C 7C 93 70 8C 35 37
 84 EA 7B 9F DA A7 42 D2 13 B8 26 5D 7D 46 B6 A0
 BB DE AC 19 43 0E D8 F1 69 B3 A8 52 C3 CD BE 50
 6E 67 FE 89 E9 BA 96 47 6C FF 86 F0 4B 6C 60 42
 4D B6 8B CC 4C 3B 7B CE CD 0B 4C DB 8B 1C A4 89
 71 36 9C B2 D1 8D C0 1A 05 F5 56 84 EC AE B5 8D
 B1 57 E4 F3 0E D0 57 C6 B4 BB E4 80 BF 17 85 70
 18 AB 48 3D 7D 51 58 13 89 45 30 A1 81 AA A5 DE
 E1 8B 9F 8F C5 2E AD BF 3A E1 A7 87 E6 03 1D 23
 7B 07 BA FE AD 29 F1 DD B2 E5 BB 35 B7 CD 45 C4
 1D D6 08 6E 55 3A B2 47 CE FA 8A B0 FA 0A 08 4A
 34 26 B5 98 99 D9 66 4D 3C EF BB 86 00 9E 4D FC
 22 5B 6C FE 4C 93 B0 9E EE ED 14 00 EA 26 D1 25
 B5 EA 00 F6 09 6F 3F E3 93 D5 58 9F DF 74 AA D0
 C3 5B 47 1E 57 76 44 23 71 06 82 54 15 6A B5 50
 3E BC 37 04 2B D7 56 B5 1A B9 45 14 99 95 64 5B
 2B 63 AC F5 AF 38 0C 75 70 93 F1 6A 74 30 AB 58
 FC 81 09 6C C1 3C EC A6 2C 70 7E 09 00 8F 3F 34
 8D 63 85 FD D5 F7 C0 39 77 E0 51 F7 A6 EA 1E 5E
 17 6A FD D1 5D C1 99 F8 DD 52 54 8E B6 F2 C5 9A
 B3 1E 7B 68 CC 06 13 DB 22 CB 8E EC 2D F5 2C 8D
 25 76 83 DE 24 90 7F F9 FE BB C4 06 2E F7 C4 AE
 F0 CA 59 3B CA 7C 07 BA BB 51 96 8C 7D 90 FB 17
 50 10 D4 28 F9 1F 64 72 7C C6 90 D0 93 EE 71 7C
 8A E7 43 EF FA C6 B6 33 97 F6 3B 3B F0 3A AD F1
 1E 37 D7 64 58 ED 42 84 50 28 29 1C 83 0A 12 3D
 20 2E 82 49 C7 E5 76 E6 D2 F3 A1 5B 09 18 15 5D
 54 83 B5 09 3F 29 70 BC 72 50 FF 18 35 A7 BC DE
 E9 59 36 9A 81 89 BE 81 BD 17 73 CF D1 83 EC 4E
 A8 19 34 A2 88 D0 44 29 82 E4 F0 1B 74 84 11 CA
 21 6C 2C 3C 41 92 00 08 0E F0 43 D2 B0 76 3A 2F
 4E C7 8C A8 63 DF 05 FB 47 B5 22 4D BA 6D 00 78
 BE 25 A5 B4 82 A4 04 69 89 4B 5A 6B D8 3C AD A8
 09 A5 4E 50 B3 31 B0 3D 57 D8 73 A1 5E EE CF 22
 B2 E2 C7 18 27 33 46 A7 FC C1 8D E2 BA 07 7A B8
 24 14 8E 78 39 74 DE 29 93 3E DE B3 6E FA F7 C9
 EE 14 4B 8E 6F F1 12 1B 6B 01 DD C6 47 6A 7F C1
 D4 9F D4 1B 4B 49 50 AE 67 70 AB C0 1E 19 43 1C
 23 DB 28 DF 06 46 5C E1 40 F4 A4 E9 4E 05 9A 3D
 30 CF 01 83 CF 5B EC F4 E9 A0 F6 E3 29 DA 7C 9A
 CE D9 28 46 E8 96 7A 1A D9 5B 18 43 A5 F4 4C BF
 1F A5 F3 DE D0 49 3A 80 AF 69 84 D6 1E 08 C0 43
 87 87 37 DB FB 0A BA 68 49 AF 4A 68 E9 B5 43 BA
 B6 6A 49 DF 96 49 86 65 D3 DD 5D F4 A9 71 A6 6B
 4D 22 CC C9 83 B3 6B 62 5D B8 01 A0 8B 69 F6 0C
 26 C1 DE B0 86 B2 82 C2 93 92 C1 CA E9 67 D6 EB
 45 16 A5 FC A2 AA CD 4A 08 A7 A1 FC FB E8 57 C2
 A0 B5 AA 0F 78 2F AD A9 2D DF 41 D9 F1 00 8F 99
 4A 92 FA DC DF 9D 77 E0 08 97 DF FE F4 8E 7F E3
 92 35 61 D4 2D 00 7D CF A4 87 7C CB 20 08 3C EA
 F8 C4 04 79 72 07 9C 7E 99 B4 BB 33 6F 1B EF FA
 2D C0 35 B5 29 8A E0 CC E7 B3 7E 39 32 79 53 20
 68 09 41 37 09 0F BB AE 39 F0 35 67 95 70 3F CE
 F4 05 3F 32 5D 03 29 50 60 EC 32 F7 C4 5F CE 2A
 D5 A7 8A E2 20 35 18 14 27 BD 15 FC 82 71 EC DF
 93 43 CB 94 48 98 A5 84 1D C1 31 60 79 58 30 08
 A3 E8 CA 63 D8 6D 60 DA 5C 5F 5B E0 C3 9F 5B DA
 3E F6 89 CD A7 6B 41 00 62 58 8E 0F 93 62 81 39
 4A 34 02 B6 CA E8 A5 25 AE DB 77 4E 0A 17 66 54
 4D 1E 0C F6 77 F2 DD 2E ED 72 8C 95 CD BE 82 36
 C0 97 46 1D C9 98 5A 5A 2E 1D 69 77 10 0C 19 1B
 9C 5C 06 41 EC D9 2D F6 42 16 CB 6C C6 BC 6D 01
 58 3E 79 0F 99 65 F4 59 B0 F2 77 3B 57 59 90 9B
 B7 7C 03 10 1F E1 C7 E1 A8 D7 56 F7 A9 58 96 F7
 D7 FD 34 C0 AE 24 31 B5 7C EE 37 7D 0C 2A 4D B0
 DC 2B 2D 45 78 EB 5F C4 E6 19 C0 3F 8A 9F 6E 92
 93 11 E1 2B 18 79 71 1F 66 BC B2 80 61 C0 31 C5
 06 50 1F 09 6C BF 59 82 48 E9 3E 14 CA 6A 62 2B
 43 0E 78 B9 5C D0 0A 2D 71 6C EB 77 5E 6F E5 5C
 BD D8 81 53 E8 AE BA 37 98 C7 0E C6 F1 2C 51 87
 6E 0B 0C F4 0C 5B 1D 75 00 4C 42 A7 3D E0 F2 12
 06 90 A1 F1 51 CB 1A 7F C5 69 EE D8 34 5A C1 5E
 9A 42 0D 9B EF 76 06 FE B2 50 EB B5 79 C4 D7 35
 E6 59 6D BC D4 AB E5 2F 6B 52 8E 72 74 51 E1 88
 93 44 36 29 E4 C3 99 9A 0E F9 94 96 38 36 69 36
 7B 8B 83 88 75 64 48 59 87 DC 5B 84 C3 B0 3D 11
 64 41 32 D8 45 C6 67 3F E6 AC F7 A4 70 29 0C FB
 5E D1 EC 5D 83 84 19 AE DB 85 48 5C 2C 8F 34 2C
 AB 8F 6E 35 55 1F FB 57 44 2B 88 E0 63 11 02 4A
 EE 54 BC DC 93 09 12 8C B2 30 8F C1 11 67 8F 36
 E5 06 D9 BC 54 B3 9C 83 2E A6 08 66 C7 F3 96 1E
 7C A0 1E 17 34 5A 79 89 C2 2C D4 FE 76 73 8A 0A
 FD 38 4F 87 C0 16 35 56 76 9B A4 15 9E BC E4 88
 A6 5E 8D 5A E3 80 39 70 A8 EC 45 5B 10 BF 82 FF
 81 49 AB AE 21 A2 FC 3D AA 06 1C 82 46 DF 3C 12
 65 E3 E1 1D BB 8F 3D 6F 1C F6 C4 8B 57 67 C4 43
 F9 87 12 51 2A 15 39 58 D3 37 30 48 7F D1 03 57
 03 23 B0 7D 70 28 28 50 15 47 9B 21 D5 29 27 FC
 89 D7 8E 25 1A 4B B4 9A 06 13 78 89 41 52 C5 E8
 5E 9B 83 75 9B 08 EF 9B 30 05 86 81 C6 52 8E E9
 F0 57 50 B1 15 48 FD B6 FE 36 85 9A 91 E3 B8 55
 ED 41 52 78 AD 16 57 8F 32 A1 D9 51 FC B5 2B 85
 44 E5 6D 6A 1B FC 3B 02 FD A0 52 84 37 7B 4B 52
 B8 C1 43 40 07 33 F1 0B 62 9C C4 F7 B0 5F 00 5C
 B9 FB 4B 83 42 E5 44 1D BA A0 24 24 F9 4C 8F D2
 D8 1A F7 80 1C FD B4 8C 66 07 EE 28 36 C3 33 93
 88 1C 8C 6C 32 54 DE 33 50 F6 8B FE F1 F0 B5 5D
 BB 2F 97 15 98 BE D1 32 86 F5 81 C6 E1 75 20 E1
 62 3C F2 1A 1B 27 E7 3B 9A 1F 94 43 3E E9 9D 84
 E0 D4 3F DC B5 50 CF 23 6A E3 63 BD AB 5D C0 E8
 B4 33 90 20 EC 76 AB 7B 4B 36 EF 9A FD A8 1C E2
 49 A7 96 55 A5 82 55 C7 BD B3 8C 2D 84 87 F6 8D
 30 75 C9 3A 77 97 D6 44 AD 7B 37 A3 8E B9 59 E6
 14 1C 03 F4 F1 46 95 A1 0F B1 2F CC FE 09 4F 40
 1A 69 E6 7D BC 69 BE 78 5C 21 49 C1 18 D9 C6 DE
 31 DC AA 35 81 91 E6 D9 D0 B4 C8 4C D6 35 35 D0
 B9 7A 89 51 DB B5 01 A6 93 2E DA EF D7 FC 15 BD
 B6 39 26 D8 86 12 C0 9A 28 4C F3 6A 6B 40 48 28
 60 39 E6 AC 57 73 98 51 B9 B0 DA BC 86 20 FE 49
 57 82 03 4F 77 6B 09 8A 64 06 C0 0C 2D BA A9 A0
 E0 D3 A8 12 6C 4E 45 E3 35 2E 7D 33 1F 1A 98 8D
 A5 F2 3B DF E2 CA A8 D4 88 38 96 18 3D 08 6B 77
 DF AC 4E C2 C3 14 AC 2E 64 76 96 B8 18 5C CC 24
 9F 40 5C 77 8F 1B 67 0A DB CF 31 27 AE E9 DC B7
 28 B7 C8 12 52 18 8D 33 19 8E 1A 9E 6E DC F3 3D
 D3 CA 49 42 4E A8 2C 6C 99 BE D0 26 4F 4C 9C 34
 92 09 45 D4 4E EC 8F 04 04 7A 54 1F FE A2 82 BB
 A7 D7 B6 BE 6B 5C BD 02 50 62 80 E9 AB E5 20 9C
 08 7D 6B 41 7F D5 33 AA 1F A6 DB 4A 47 63 58 7E
 30 E1 96 25 E4 C9 4C 3B F9 26 10 6D F5 71 A9 32
 C8 79 7E 51 F0 81 07 DF D5 33 93 FA 2A 78 37 95
 A7 96 B8 C1 CF 8A 22 69 0C FE 49 3D 91 EF 75 DC
 87 3F D2 70 9D D6 30 65 3E C8 D7 DE BE 99 DA 50
 D2 BA DC 4E 69 35 2C 21 9B 4C 4B 31 12 7D 7B CB
 FA F4 73 AC 36 C4 76 E1 15 FA 83 4A 5B 06 E9 6C
 A8 55 F8 E9 D0 59 E7 33 C6 91 88 13 60 8A FB 74
 46 EC 5F 03 81 EB CB D2 05 16 E7 84 60 94 73 69
 F8 13 C4 53 B0 71 80 B0 97 93 AD 83 F7 21 D2 83
 2B 38 FC DF 77 62 78 24 68 A4 E7 36 CB 6F 91 B7
 FB 83 F2 C9 B5 5A D8 C5 16 C4 CE D8 15 30 06 C7
 F4 32 BC CF A6 0A BF 68 59 9B 08 01 5B EA F2 76
 AB 43 D0 35 63 DB AF E0 6F 05 08 C8 EF EF C8 C7
 29 33 89 D1 6C 6F B6 7E B7 33 2D 10 CB 89 AF CA
 FA 95 44 B4 C7 81 9E AA 3B 44 1D 23 22 F7 B5 8F
 86 25 50 9A 56 F3 78 C8 54 6A BF 00 2F FA 4B 7C
 B1 E0 D7 6E 94 24 F4 AA 6B E3 32 A2 05 42 FE E6
 5C 16 0C D9 D7 C7 A2 09 90 43 93 B8 76 E8 E8 CE
 85 EB 73 E6 94 25 1B 83 18 18 88 1B F9 D4 49 7A
 EE FA 4D B0 91 F2 E4 93 EF 0F B2 C7 BE 3A DE 8C
 7F E4 90 09 41 49 86 CE 3C E7 04 FF 87 2A 6B 3A
 04 6C 24 58 35 31 3B E7 66 AF 0A EA 46 B3 39 45
 B1 B0 60 0C 3B A7 F0 48 16 AA 05 3D B0 72 16 FB
 93 27 4E A7 62 2D AE A9 55 B3 3A E9 A5 BD 90 06
 B0 FE 58 98 C4 2C 1E EA 96 AC 68 89 A8 D8 B3 7F
 13 AA 30 C8 5D 17 AD 5B 80 E2 FB F4 F1 EA BE 60
 9F F5 F3 16 90 D8 A8 80 EC 4F E7 1F 42 64 4A 47
 47 19 72 0B 1F BE 5A 9E 1B 62 E0 AD FB 2B D0 67
 BF 82 98 A9 9A A3 97 21 99 BB B0 E1 32 CA 29 8A
 F9 22 78 9E D8 E3 65 95 ED 03 70 57 BA 80 EE 6E
 3E 1F C9 32 DF 03 43 46 40 18 DE C4 10 08 3D 3C
 DB BB 5B 55 3B AF 2E 3D D8 6D 3A E4 AA 69 57 9A
 4C 5A AA 6E 0A 2D 81 D1 61 E3 EF 45 C3 BA 94 76
 3B 26 27 0B 72 4F FC 16 6B 17 06 94 5F 28 A9 42
 D5 3E 26 14 FB BE 34 F2 DF 9C 44 DD A5 BE E0 74
 E9 74 CA 69 0D B0 4D 0F A8 40 23 79 DA D7 9F 63
 3C F7 9D 7C 03 8B 63 EC EF CD 42 DA DF 5F 56 9C
 A4 47 A4 1D 76 1B 0C 35 25 25 E5 24 17 17 3E 72
 DD 0C 83 D0 56 DA BE 11 56 29 F1 8F 06 81 7B F5
 03 B3 25 FE 81 A6 86 14 EE F6 EE E1 46 97 43 B2
 B5 FE D2 37 62 6E 7B 81 C9 B4 66 8F 77 57 91 84
 82 9C E6 31 D6 D6 1B 10 ED 4B 27 A5 D4 F0 4C A0
 85 2C 3F FC B9 73 07 56 04 4D 5A 57 5E 54 2C E5
 CE D6 0B BA F8 8C 64 20 82 C0 61 B3 FC 22 23 83
 BB 89 01 29 D3 E0 A5 C3 30 A0 10 96 B6 C1 99 76
 55 29 3A 29 F5 4B B7 69 1C B2 7A 59 D3 57 DE A9
 35 11 6C 99 07 B8 91 9B AE 94 7E 4B 58 45 80 05
 11 E9 3B 99 1B F3 66 56 4C 15 64 6D 20 A6 30 EF
 A3 92 7B 58 D5 F8 51 DA 7B D6 43 92 11 B5 B5 A8
 EF 2E 41 90 D6 4D 11 28 18 93 6A F6 FD F4 4A F5
 47 A6 2F 0B 06 DA C3 46 5C FC 18 84 53 0A 6A 86
 24 39 52 D2 1B 51 13 A9 9A 9A C9 37 05 A3 B8 36
 77 28 D7 2E 51 BE 1E C2 B2 CB 75 2D 03 D4 0B 4E
 23 68 8D DA D8 68 B9 CC 43 13 07 BC 58 AF A0 72
 0E F3 18 CF 75 83 3F 4F 0B F4 E7 18 6E CF C6 15
 42 E2 D3 6A CD 68 E4 FE 9D 71 D0 FB 7C 41 BF 2C
 AB F3 9C 5B 25 23 66 50 BF 62 14 27 1B B5 BB 25
 3A 0C 66 12 6C 97 E1 F8 A1 D6 57 36 A6 AD 17 31
 3D F7 14 DB BF B3 90 0F 8C CB 9A 42 DD E8 6C 28
 A5 0A FD 38 FC 79 F0 6E 2A 5A B1 55 6B EE 90 81
 61 92 5A ED 32 8A 10 2D 5B 61 92 6F 50 47 EF 09
 F5 09 98 9F D1 44 96 EF BE 6C 02 99 D9 41 6E 05
 EB 5A F0 B3 FC 7F 0F 63 C4 2E 37 1A FC D9 1E E4
 54 A0 1C A7 B0 39 81 B0 F9 04 1D 2A 43 D5 D9 4A
 36 2A B5 44 27 B7 D5 D3 9E E7 4B 87 87 48 9B BB
 F9 A0 B9 C2 C2 6A D4 78 93 F6 5B EB ED 25 47 F8
 FF A8 E1 CF E0 FE B6 2C B5 37 6A D4 6D 89 4B EE
 25 FD C1 06 EE 0F D6 44 D8 BD A3 9B 3E 5B 13 F0
 81 D5 5B A3 98 E0 2A 0A 6E 6B 69 4F 51 C0 57 23
 1B 6B 0B 0C A9 DC 47 00 ED 7F D0 C5 D2 99 1B E6
 95 1D C3 E1 F7 CE AE AB BC E3 EB 4C 27 72 F2 97
 54 05 18 40 FB AC 8E 5B D9 2A C8 0A DF 97 CC 64
 C9 07 40 AE A3 1F F0 03 D9 3A A8 53 FA 14 30 51
 58 6D 4E 18 23 FE E2 A0 AA F8 76 51 C9 24 64 49
 01 0F C6 5B 77 48 44 7E 81 3E 8E 45 E5 FE 9F 8C
 9B 3D 0E C7 FA 32 85 CE 9D 87 A4 20 DE ED 93 DF
 6D 64 A8 4B 53 03 20 72 C9 D9 15 38 A9 83 86 F0
 F7 1E D2 47 FB B7 D9 5B EE 29 CA C7 A5 79 B9 4E
 FD C9 39 52 32 BE 61 09 74 78 E2 E4 D9 4C 4C 9E
 A3 22 51 9D AD 57 46 6F F7 AB FF A0 D9 F1 0B 4D
 D7 4B A0 CF 7B 84 35 A0 F9 40 07 4C 4D CF 8D B1
 61 1D 6E 1E 00 84 2B 87 22 3A 76 DC 82 E0 78 E4
 B5 EB 51 AE F5 94 1B A6 F8 4B 92 8F 4B 4D 8A D2
 23 BD 65 87 E5 82 B4 AE 23 BB 74 91 93 C5 72 0F
 9F 6B D7 3D 77 99 D5 BD 75 9E EE 49 5F FF D7 7F
 0B E3 ED 5D CC 7D C5 06 CF AB E7 EC 4D 7A F8 DF
 7F 83 53 E5 B9 0A C3 8D A4 02 FE 7A 22 90 D2 ED
 AC 12 FF 45 D5 D4 1A 2A 83 2D A9 E3 47 DB E4 64
 B8 DC 0C 64 0B 24 B7 B4 58 90 7A 1F E9 6B A6 3C
 82 6B AB A5 02 AB 59 AC 20 91 30 FE FA 9F 5C C3
 93 38 C3 8B FD 3F 84 40 DC BD 9A BD 4A A3 03 5A
 6B 79 AF F0 39 72 1D 57 60 A6 E3 FD 25 7C B0 1D
 54 A0 70 EB 0A EC 02 DF 53 BA DC 9D 41 24 DF D3
 C1 A1 83 F2 FE 78 61 6D 05 46 F9 C9 59 77 29 95
 81 13 A8 DB 28 46 C0 F0 DA 80 C7 7A 6E CD 63 80
 CA 2D 6B 0F 9B 14 4D 09 07 2D F1 6A 71 35 FA 3A
 81 B2 DA CA D2 75 AC E8 45 90 EC 53 F9 30 DD F9
 87 D8 0D A3 7A 1C 4B 5E 81 DD DC 63 CC 67 B5 A6
 60 26 7A 48 E8 A4 40 57 CD 6A 2D 88 EC 9C 72 76
 5E 1F E2 23 4D F2 74 C1 68 82 05 CD 2F EB B1 4D
 D9 3D AC 81 33 E9 74 B5 4D 3B 5B 70 00 76 83 F3
 E3 EC 12 DF 70 00 94 7F EC 4E 6E 9C 3B 47 74 F2
 12 59 5B 8B E6 E4 7D 0D F6 3D 7F E0 2B 16 F8 B1
 5A E7 70 60 6D AA 28 8A F2 32 70 19 50 C7 D5 16
 3C 3D 5A 93 1D 6B 47 06 75 D2 98 0F 96 F6 1C 80
 95 D5 3F 32 7B 6D C1 F3 F1 FA A3 2A 3E 6C 62 4D
 EB 59 EE 3E FE 63 31 53 57 5D 1F 01 BF E8 47 13
 CC 66 23 A6 F5 BF 1F 4C 1C 44 0D 36 EB 1E 89 CE
 5E E6 41 0F 77 A3 4C 51 70 A7 7F 4C 64 46 AD 3F
 1A 23 39 D7 6F 2F 7E 5D 22 7C 30 40 05 2B 40 FC
 FC AF 7C BD 15 D4 AD 02 3D 00 D5 7C 0C ED CB 66
 4F 80 08 25 1F 5F BE 45 60 CF 8F C9 97 5B 50 BD
 00 12 9F 2D 3B 4C F5 00 9B 1B FA 93 83 FD B7 EE
 BE 15 AD 26 03 82 07 A6 AC D1 3B BA BD 07 BD 6A
 8B 30 51 36 1C 03 79 E7 12 71 74 9C 6C 63 0E 7A
 57 9D 9C DE 67 2C F5 D5 52 7A BB 6E 76 A6 21 64
 BC D5 5C AD D5 DE 56 B9 C7 80 1B F7 92 DA 0E EC
 0B 6D 01 82 1F 4D 09 9D C5 66 D3 B7 7B 79 CC AD
 DB 0B 04 BE C0 52 40 BA 59 0A 05 B3 6A 77 B8 9F
 AB 73 3B BF 5D 0B C1 A6 F3 3C 64 06 F0 98 67 57
 4B 1C CE 07 79 87 1F 2A 36 00 70 A9 A0 72 26 8C
 45 8F 71 0F 91 0D 5E 63 4E 5C F2 9C 55 CF C4 C1
 5B 67 78 26 B8 B2 BE 5D 2C 11 3F 36 1B 6E 7F 73
 C4 C0 1B 13 E0 5C DE 79 3A 11 38 FD 26 C3 3F 56
 E5 0B 0D 93 BD 56 AE AC 1F BA 8A 9E 78 E5 FA F1
 12 B3 D0 4B 9D 23 AD 7E 28 D4 04 B7 A5 BA BE 5F
 90 8C C3 5B 6A 10 6D 92 71 70 18 65 F2 FB 15 B6
 66 AF BB 63 60 DA C5 26 F3 89 E1 C6 EB 92 A4 AF
 09 D1 31 0B AD 20 ED A4 D8 A1 04 55 F9 61 98 1C
 58 55 9C B3 80 2D F3 5D 1A 25 D7 84 8E C6 52 43
 9C 79 E5 87 F3 12 42 F5 4F 9C 12 DA BE DB 1D AF
 6E 23 9C EA 7D 47 FB 75 79 0D 3F 7A 33 A5 A0 AE
 B7 37 58 94 E3 E5 EC D6 92 F3 0F F7 4C 66 C1 CE
 B4 D9 55 F9 7C D5 43 D4 0B 8E 07 CE E2 14 40 89
 69 F0 66 4E F0 EB 7F 06 2C FA 81 26 F6 DF 82 14
 76 22 5B F3 C4 0A 98 50 90 0C FA 09 E5 5D 89 A7
 A8 00 57 48 34 56 0A DB 7B E1 0C 05 7C 6F 93 5B
 A3 1E EF A3 A8 56 A6 56 01 BB 32 FE 52 AE A8 59
 C2 5E 51 86 F0 19 55 B7 1C 64 89 4E B2 C2 96 84
 D5 19 52 E6 0D 00 75 E9 72 30 D2 4E 77 AD 33 8A
 AF 6D 3C 2C A7 13 C9 9B 17 C8 62 A6 54 D9 43 96
 92 D8 2C D5 C2 86 DB C8 15 D1 73 47 B6 E8 D0 31
 28 AE 0B 60 2B 7F 2B 5B BB AA B7 AF 03 2E 24 FF
 DD 72 4C B4 93 57 99 BF 4D BC 24 0B DB E1 C7 94
 F4 A7 B4 0E 7B 25 FF 50 49 1A DD BE F5 35 C1 75
 51 2A 7A CD F6 93 AA 3A 19 72 6C C1 DA 88 8B 6D
 92 77 E5 D9 A0 95 48 63 04 0F 51 E8 9D 60 B5 B1
 24 B0 CE 77 B9 84 21 E9 56 1B 12 78 EB 6B 9B 0D
 5C F2 FB 23 67 30 79 76 6B 20 BF AC 93 41 64 3C
 55 FA 83 8D 61 08 C3 EC D2 FD C3 10 69 3B 5D 10
 F7 E6 6C 54 14 9D 9F 74 B0 35 9F 5A D8 DF 5C 70
 BF 0B A3 DF AA F1 54 09 33 AE 1D EF 8E 0E 82 4F
 21 91 CC 10 85 30 87 F1 1E 45 42 31 13 D8 07 78
 7D 82 AD C5 6E 41 3B C7 9D 37 6B 5E B4 B5 BA AF
 66 86 EC 7C 7B 42 DD 2C 09 AA 9E 9B 38 06 8B 63
 4A CC AA 57 5F 47 E8 0B AA 26 96 C3 2F 80 83 65
 42 73 77 EA 7A 95 32 6F 1B C8 A3 2E 96 44 24 D0
 74 6A 3B 2C E4 57 19 5E AA 77 EE D2 7B 97 17 AF
 EF C1 0D 4F 59 46 48 8C C2 50 69 F4 E1 38 9E 6C
 80 90 AD E4 66 5C EF 9A 3A 33 D8 AA 85 30 99 D7
 19 8A DB C5 31 5A BC C3 7F 32 06 2A 5E 08 7C BF
 E2 19 4F 52 34 4E 7D 04 22 1F 03 F5 EE 0E 95 97
 0F 9A E9 F1 44 2C D2 6E 3E CF 11 92 FA AE 00 21
 EF 7A E0 15 81 C8 FB 90 F9 2D 81 D9 CC F1 65 B5
 57 20 A2 F5 49 B4 5A 96 BA A6 36 2A 6C F0 21 37
 FE 7E 9B 27 82 E0 BF E7 A0 A4 D7 9C 3B E1 A4 85
 79 E9 9F 88 58 0B D1 AD 7E C5 ED C6 0B 1B A2 9D
 4D 2A FC 52 E7 92 4C B7 51 42 FE EF 0E 2E 5A A4
 82 1B BD 16 03 0D 79 31 73 D8 37 1D D4 FA 03 B8
 FD CB B9 3F 4E B7 C8 0E 3B 71 B3 12 7A 98 81 10
 02 4B 24 63 5D EC C3 DB 54 1F D1 BC 7A EF 04 9E
 EC C5 CD E6 39 6D 6C 53 5D 34 D5 5E 27 6F C3 CE
 BF 02 35 F5 27 BC 32 2C 87 49 C6 72 E1 50 6D DC
 AC D0 F1 CB 2A 53 3D 9F ED 4B 49 85 F8 92 39 0F
 28 AE E7 23 33 EF 9B 3A A2 78 5E C8 C4 D7 03 60
 B7 24 6D 0B 58 00 0E D8 E3 83 2F 93 7C D8 3C 42
 0E DF 64 06 35 74 0B 2E FB EE 59 0C 4F 04 B6 3D
 DE 86 14 CD BC 51 00 31 BF 3D 53 12 B9 BE 78 5C
 5B 11 A2 4F 64 7D 11 0F 6F 94 A4 B0 B0 4F FE DD
 8D ED 45 D9 36 F5 37 0B 23 39 D8 40 B1 0B F3 1A
 51 42 56 C0 9E 6E 75 F0 7F 4B A8 85 9B 11 F3 4E
 3D 52 39 FB C1 A7 68 CA 85 DC CB 9A 72 53 70 F4
 20 93 F3 B5 47 EB 36 2F 38 E0 EE F1 3F 8B 49 E3
 F2 1C 83 AD 41 E9 D4 EE 2A 42 59 92 D9 6D 71 2F
 1D 99 BB 12 BD B4 90 85 BC 22 F8 A6 BE 03 7F 5D
 FC BA 04 F5 CF D1 3F C9 7A 13 73 D6 D1 4B 23 44
 44 81 05 9B 86 91 F4 FF 35 9E F1 A1 37 12 CC 76
 21 20 06 A2 A2 7C 98 64 A5 8E 38 09 27 2A F5 58
 8D E7 58 AA 2D 4D FB 3C 47 FE 9E F0 E7 8D 57 F5
 BF 1A 9F 8F 1C C9 79 77 E3 24 CA 4F 98 88 C3 DF
 F2 93 9D 6D 87 C2 8D AC 7F 52 06 9D E7 42 86 B5
 81 76 22 8A CB 75 2F 50 E1 4E C4 08 A5 12 B8 34
 03 EA F7 D0 6E 94 93 9F FE 0E 6F 2F 8B E6 2D 2E
 FF E3 DE AE 7E 5A 91 38 CE B4 3D 13 72 E0 61 FB
 B5 54 50 BC 5D 54 98 DF 49 B2 65 E1 EB FA A6 38
 9D B8 03 73 CA 22 32 49 62 17 4B 24 CD 27 CA 01
 4B 52 71 AD C9 C6 F0 66 A8 D6 9E EF CD 46 8C 7A
 CD 2B 69 5A 84 D2 62 CD 6C F8 A0 F1 B1 3E 6B E3
 FC A6 62 56 15 73 E1 3A 99 88 68 F9 D9 CA 18 82
 23 CD 62 6E D6 51 C5 86 78 1D C6 D6 72 18 61 63
 E0 8B 7B D5 4B 1A 87 13 A6 EB 30 40 32 3A 5F 1F
 AB BB EE 20 56 E6 57 BC F5 4E 90 F7 AD 7E 0A D6
 FF C9 D7 3A 76 F1 DE 25 36 5D 41 65 A8 DA E5 25
 48 50 77 49 AF F4 9A CC 7B 92 CA 2B 04 70 E5 7E
 EF 90 4F FE EC 34 1A 9A 24 59 3D 57 2E 34 51 2A
 0A CE 92 71 9E 74 64 17 AB A4 EF 3B 05 88 6C 36
 C3 35 EA B3 62 36 74 5F 87 8D 5F 19 27 6F 64 48
 EC BA 02 12 D4 D9 17 A7 2B 31 7A EA 4C B0 50 E9
 A8 B7 74 77 7E 20 B6 27 F1 E3 ED 41 13 30 67 05
 86 96 99 89 44 86 31 99 D3 0F D3 EB 40 D1 E1 6E
 E5 30 98 0A 27 45 8A F4 1B B4 CA 96 93 53 C5 8F
 3D A1 8B DA 06 B7 A7 41 68 B8 E8 C8 2B 94 0E 4C
 D1 1F DD 7A C7 CD E2 2C 41 F7 81 D5 72 70 02 EB
 0C 3B 2D 3D 78 4F 8C FB 4B 78 A6 D9 70 C3 2B 28
 5A BB 6F BF 65 A9 27 B2 DA C9 CC 2D BF D6 32 5E
 C8 D9 26 91 23 D3 8D 80 19 C3 8C 06 97 D2 DD BA
 9B 19 CD C1 AB 26 6A F6 B0 A4 5B 1D D6 38 09 7A
 FC 21 A3 04 28 DB B7 35 13 BB 65 D6 65 E6 AC D3
 B7 B4 DA 4A 3D FA BF 21 49 2F B4 1A 4F D5 86 80
 47 D7 9A 61 5C 5C 00 8E E8 AC DA 72 68 20 D8 0C
 D5 56 2E 5C B7 F2 BA 31 85 C2 1C D0 7B FD 5F C3
 12 C9 41 3F 9F 76 8F 88 64 11 69 17 F3 BF 7F FD
 3C FF 20 E6 E0 07 41 AB DF A5 97 F0 9E 4C B8 FF
 DB 3E A8 B0 0B D4 A4 E2 CC 57 D1 44 0C 78 B7 CC
 CF F0 53 BA 73 CE F6 D9 86 7C B0 3F FA 18 A2 5C
 3E D8 36 F7 F6 D5 E1 62 DA 28 73 59 EE 18 83 07
 D0 9C CF 71 51 C4 3B 2D 84 01 60 68 52 B1 B8 5F
 2B F7 9E FC E7 57 A7 8C 64 F5 D0 3A 80 3E CD 6B
 54 AB F0 8D C4 E2 F5 A4 8F FC 0F 5E 94 31 5A 0D
 DD 1D 7F 10 1A DE 37 A7 C7 88 04 AE EB A3 18 F5
 C8 38 73 92 EA F8 B3 D9 40 8B 2C 0F 88 8A AD 7B
 C1 7C DD 30 CA CC D7 09 9F 2A C7 0C 98 E5 63 2A
 89 1B A7 50 44 14 CE E6 BF 87 9F D0 45 3C 2A 71
 E5 DA 62 06 06 B3 B2 3E 6A 3C BA B9 9C 5A 38 B5
 D0 45 7B 72 55 28 64 72 E8 55 5D B2 D2 23 1D 3E
 49 E3 0F 18 FB DE 99 86 B2 5A FA 39 88 B0 7A E0
 E8 3B 35 75 C5 B8 86 EA 9D 72 03 02 15 B1 F9 8C
 0E 00 73 AD 4E 57 23 69 6D A6 7E 0D 72 BE A8 6C
 95 F9 4A CD C7 94 98 38 52 AD D8 E9 CB 21 A9 EB
 D5 0C A1 7E 05 D8 7B B8 36 E4 DC F9 D5 DB E4 C8
 EF 59 D7 CA 92 4D FE BB 1C 3B CB 13 66 79 FB 4B
 98 5D 48 7E 9E 02 62 AE AC DF 99 13 93 79 50 07
 13 3F 89 3E 2F 43 42 A4 A6 DF 66 92 BD 96 F8 D5
 31 A1 14 56 35 65 35 5B 2F 5A E7 D6 A6 53 E0 0C
 C6 AC 9C 5E 9D 7F 3C 88 51 9B AD D7 41 6B ED 64
 4A D2 4F B9 5E A4 5A DF 04 34 9C AE 31 D4 FC 85
 C1 95 98 76 11 5C 10 63 02 4D 27 0B A5 41 B6 D8
 20 35 5E 02 3D 8D 49 C3 95 48 8A 6C C1 7B 07 B3
 14 95 2C 05 65 90 16 B0 39 9A 61 7F 8B 5D 53 CA
 53 8A FC D3 49 F3 53 B4 DF DE 68 39 12 90 8A F6
 A1 41 F7 3B 54 26 33 C5 AD 14 F7 CA 46 07 B3 FB
 53 25 E3 81 A4 8B 7F 43 39 75 DE 38 21 AF B8 EC
 CE 5E F8 B8 9A E3 C5 B5 91 11 E5 D4 22 7D DD 4A
 92 78 AB 5D A0 4F 4E B1 A7 1A 69 78 DE 05 AF DB
 D3 B4 A3 69 3C 49 EE 5A 9F 61 87 34 CC 5E 08 C8
 ED 59 84 E7 4C FD 5C 51 6D 0B AB B9 B0 2C 0F 15
 C0 96 4A 87 2E 5A 89 F6 E0 84 68 7B 40 21 DD 97
 0E 0A 36 68 FF EC AD EB 1A 27 2C CC 57 95 7B 39
 C0 6A AA CF 50 E6 87 24 FA FB C3 26 83 2E 28 B4
 13 05 39 FF B9 D3 29 C1 76 17 70 2D 0A 34 85 30
 50 EC FC 38 94 8E 9A 21 D2 BA 13 34 C3 57 49 BD
 68 42 13 17 13 0B 8B 81 B0 9F 71 24 E0 AE D7 D6
 FA 33 E4 98 62 2B 5B D6 9E B3 03 E8 2F A8 2B 4E
 A3 F1 2B FE A9 2C 95 C1 2A 04 50 25 BD 4E 8D 2A
 57 31 8C E8 CB 73 FF D6 74 C9 EB 97 60 39 14 7B
 27 FB 1B FC CF C8 BA E0 2B 70 20 D1 D9 2A 25 DE
 70 B0 EA 16 B7 9A 5C EC BB F1 54 9E 79 CE 0E 8F
 BF A5 EC 17 14 01 C6 E4 82 B5 75 3F 13 F2 1C 37
 C6 FE D4 D4 71 63 8A 1C E7 BC C5 52 FC 28 BD C0
 AC 01 A6 46 45 1B C2 69 50 D4 3E B4 0C 1F 14 2F
 F4 9C 5F D4 52 D8 CC F6 5B 09 22 B4 06 A9 EA 7A
 56 DA C7 E1 AB 8B 82 81 14 E5 6D 1F 44 04 80 D8
 5A 4C D1 05 1E 2D 67 4E 57 E1 4E 6C A5 F7 F7 4F
 14 FB 54 89 DD 05 8A C2 74 39 C2 71 3F 6B 31 16
 02 AB 2E 51 E8 53 80 C8 4B C9 72 40 D3 04 C9 61
 9A 29 91 5E 17 66 E9 7A 74 91 36 C2 94 51 A3 A6
 39 BF 18 C9 DE 96 0C B9 CB 87 F5 44 BE 07 5A 0F
 A3 8F F7 D9 30 F8 90 0A BF 0F 79 39 56 C4 59 CD
 9D 80 04 6F DC 79 AC 13 40 8B B4 44 3C 05 49 0E
 8A 50 F0 F0 F3 57 93 4F 81 77 36 64 70 4D 3C 84
 01 31 3E AF 4B E7 AE E8 E1 4B 5F 5C FB BE E3 70
 6F 28 52 56 81 38 A9 7D 7E 46 4E AB 55 99 8B AF
 B4 6E B2 10 17 41 AD D6 1C 60 4D 30 3F 34 0F 4D
 BD 6B 4F A3 47 93 9E A7 09 BB 40 B5 CD 0D E2 0E
 A9 45 7A 6D 4B C1 B0 F6 A5 18 42 96 48 17 54 6D
 4A D6 88 B8 92 55 CE E8 03 B8 14 54 D7 BC 76 C6
 64 AC 53 F5 B5 14 EC 37 92 53 21 96 68 D5 38 A3
 0E 8E 31 16 AE 17 0A 11 94 55 52 14 3C 3D 76 01
 BB 0F 1A 2D 5E EA CC 61 1E 7B B6 A5 EF 96 6F 30
 93 1B CC 3F CC 76 10 4A 50 CC 1B AD 27 04 CD 3F
 4C 86 E9 99 1A 2C D9 96 C8 92 9E C6 C7 8E C9 BC
 68 6A CD F3 AE 21 86 16 09 56 3F 3B 41 3D 77 CE
 24 00 C4 33 14 EB 3E 0C 39 A6 60 4C 76 7E 1D 70
 2E F3 D0 AE 72 27 5A 03 F7 C2 02 B6 2C 32 B8 06
 41 C1 1E 8B 31 DD CB EE 1A E9 DF BF BA 59 5C 4F
 13 B4 EF 7C 34 EB 5C 29 E8 BD 52 46 99 56 13 59
 A8 02 47 2D E9 3D CC 41 BA 86 CA 7F 62 A3 9E 27
 30 3C 05 E7 7C AF 70 A1 9B 68 0D 48 96 61 D9 0C
 CA 53 1C 35 56 A1 73 3E A6 88 40 F9 86 F0 1A 2F
 D0 67 4D DD CE F7 50 6F CA 90 A7 38 0A 96 15 3B
 48 C1 74 1B D3 2E 39 44 E2 F8 6A 41 70 56 06 1C
 56 6F 12 03 7E 44 13 58 8C 48 0E 87 E9 23 EE 28
 5A 39 78 D0 28 D5 EC 9B F7 4B A9 5B A3 21 FB 37
 ED 2B F6 D7 C2 D5 4B 9B 1A CF 7F 23 B2 99 CA 49
 40 8D 6D 5E 14 9C F8 96 07 AC 4E B3 14 13 9B FE
 7C 86 20 E4 52 72 9B 44 FB 60 A7 37 0F 26 C6 95
 D1 5F 7F 15 C7 C4 9E B8 93 35 3C B6 28 A4 B4 A4
 CF 13 45 49 22 C3 97 7E 81 C3 5D 36 AE 98 CF F2
 54 16 86 75 90 5E 29 E6 6B E3 77 74 99 83 CC A6
 DD F4 DF 54 3B 83 5B 0F 80 C7 07 6D 05 5B 8B 2D
 E6 F8 FD 68 68 AB 5E A6 A8 84 EC 48 0E B2 48 7B
 62 B7 95 F1 FB B7 44 C9 7A 85 03 D7 88 D0 D8 86
 D8 5C 9D 30 05 EA 01 85 39 96 FF 6A 58 9F 4D 93
 45 F5 23 C2 D7 57 55 13 29 C9 22 5A ED 00 08 9C
 9E 13 18 D5 DA AA 15 86 CB 50 34 E6 23 54 36 38
 72 7E EE 14 AB 01 5A 75 65 8D E4 14 59 9E CA BC
 D2 69 EA 7B B3 4F D0 01 47 8D 1B 5F 10 FD 68 41
 4D D1 7F FF 11 A2 F7 80 08 E8 A8 A0 09 A6 91 1B
 B6 A7 ED ED 82 AB 75 C2 34 75 6D EE 92 9E AB 61
 B2 10 57 10 3A EF 24 0B EA 75 70 1E D4 21 8D 01
 31 2F 0F 2E 36 B6 21 DF D2 FA 0C 2C 41 BC 27 5F
 91 22 7B 1C 10 35 07 69 44 EB 1D AE FB 98 95 B5
 75 0B 03 74 F4 D8 86 AF 12 6A 44 6C 9F 4B E0 08
 DE 28 06 E3 14 A6 76 38 65 8F 2C 70 13 FD 05 50
 DC 12 16 DA 61 63 AA 42 04 83 E2 F3 2C FD AE 40
 3D C9 D1 51 98 5B 27 EF 2A 77 9F 99 AC 41 B5 D9
 2C 6C A0 2C 98 62 B9 8A 07 8B FC E6 67 94 90 4D
 DF 2E AD 29 2D 1D 37 67 A4 20 F3 F3 6A A9 37 DF
 9A 9B 87 08 AA 3A A8 12 DE 0F 22 69 C3 A0 73 29
 12 F4 6A 74 87 73 C6 98 75 4D C7 6B 0D FE E5 FE
 A0 50 0D 29 B3 3E AB 44 16 4E F7 26 20 AB 6D 91
 A5 51 31 D5 90 23 5C 43 84 10 BB A5 A1 0B 15 44
 F1 F6 18 A3 47 1D E4 E0 AF 6C E6 96 9B DD B4 73
 00 F3 58 82 82 49 70 88 36 3C 57 36 5F B6 11 3E
 AF 55 1A DD B2 40 7F 08 22 33 95 5A A3 B2 3E AF
 EF BB FD D1 21 A1 A8 B5 FE F3 0D 7E 13 E1 0F 67
 E5 DB 3B 41 68 D0 95 92 A6 1A 5D 05 C6 A1 C1 88
 A5 EE E4 54 50 3E 87 66 83 7E AC A4 E9 54 5A 2E
 AA BC 2E AE 1B 08 B5 9B EF 85 BE C5 43 EE EC BE
 F6 F5 77 9A 33 6E 84 68 4D 54 AE 34 19 2B E8 97
 9E 17 C4 DA 2C 39 D1 C2 A5 86 16 99 0B BA A5 3D
 88 0F 91 86 40 72 40 09 86 DC 5E FD 24 D2 66 C2
 8B 60 26 BF 76 D1 2D A3 93 C2 F3 AC E8 DB 6F 13
 18 6F 0B 6F 34 D6 CF F3 9B 09 77 38 C3 2E C4 24
 F7 FC 2C C1 07 28 DA 61 B0 E6 2D 87 FA 66 22 30
 18 49 C0 F6 E8 4B 99 8A BA E4 36 58 D2 3C 6C 98
 A3 12 03 FF D1 F1 E6 8C 45 1B EA 01 9D 51 93 61
 E2 C3 D5 92 F7 85 94 3F B7 67 2D B1 A9 6F F3 05
 2D 2E 53 89 61 AC B5 2E 00 8D 55 ED DF CE 6F 88
 91 F5 9A CD 68 D8 24 49 D8 70 35 FD 81 58 C5 28
 A0 FC 7A F7 74 B7 26 6F 76 2D 3A 83 90 45 7C 0F
 02 9F F1 A6 A3 5C 6A CD E6 DF 71 BB CC 5F 70 4F
 94 50 38 22 03 51 5C C4 D8 F2 F9 AF 22 B3 65 B7
 97 9E DD 69 99 01 B4 16 D1 47 27 FF FC 32 A4 A6
 02 DB 47 CF 0F 70 F7 1F 13 83 66 73 4F D9 1F CF
 BD 21 3E A2 F5 E9 72 5F B2 69 34 BD D0 32 BB 69
 C2 85 0D 3C 5D 61 16 5C D3 44 6C F4 31 8F 0C FF
 C9 A2 18 D1 5F A3 11 CB 61 39 69 A1 D1 DA 8C 46
 D4 CF E6 4B C5 D3 36 C6 78 62 11 B1 49 D2 3C EB
 A8 00 44 4E D8 33 56 CC FD 54 AD E2 37 19 68 50
 C0 AF 1B 75 00 CD B8 EE AD 34 58 1C B7 C0 30 F3
 65 6C D3 0A C4 6E 8A 5A 0A 34 36 8E 25 C9 BA 1C
 B9 60 AC 9A CE 9C F4 84 A8 EC 26 1C 83 D0 9A 44
 73 F6 59 DF 98 CD B7 D7 FD 54 5A 8F 32 69 54 E9
 16 FA C5 EB 16 65 D2 D3 06 A9 8F 8A D4 B9 72 AC
 E8 C0 91 45 83 47 D0 A1 6D 9A 35 9D 60 5E FC 42
 D5 DF EC 8F 72 DD 2E A8 3B F2 47 F5 BC E8 7C 0F
 3C 7D 60 59 51 8B 7E 5D D9 14 84 13 46 D2 95 C5
 50 20 EE 2E 07 80 11 D4 A3 3C 18 DC B8 E1 4E DC
 9A 7B 4B 59 D9 39 3E 09 9F 0D D9 BA 76 6E 81 8B
 48 6B 11 CD 9F 76 44 86 43 26 8E 9C 40 9E 29 5C
 88 F0 E8 F0 95 A6 D5 6A 05 EF 89 8A 55 AB 55 A5
 4A 60 18 F9 E6 C5 FF 8D E7 D3 F5 53 05 53 6B 20
 78 A4 82 67 C0 56 8B 11 D8 2C 32 52 DA FE C9 E7
 E6 93 D0 3D 4E B9 1A 85 AD 94 F0 2D 93 A6 FE 4F
 98 C6 15 4A D1 EE AB D1 5E 3A 99 B0 28 03 F6 79
 73 28 E2 7A 0F 6F 63 4E AE 7B 97 DF FB 8F 09 F5
 1D C1 B7 85 35 68 78 94 DC 16 E3 D9 60 29 6F EE
 D4 1B 1F 3D CF 3D B4 48 87 F4 82 E6 89 38 29 49
 0A FA 6C 61 66 F3 11 C6 AD 45 A2 30 9E 04 66 B1
 10 4A C1 37 CC 9B 42 CE 2F 25 29 64 3F 67 FD 79
 1D C3 FE C6 F1 60 C1 D6 A7 84 93 12 01 6C 71 8C
 73 8B F0 D4 9A C3 F5 53 B3 6F 78 C0 21 3A 8D EA
 20 BA 36 79 00 2E B2 B6 B3 A0 F3 2E 60 97 E8 7C
 36 0E 39 41 F7 84 C4 06 C8 CF 23 21 BC 92 1D 17
 B7 D7 72 3F E5 80 6D A3 CB DB 82 B6 6D F3 9D 8B
 E0 A5 55 54 30 E5 62 08 A5 EB 94 72 67 7B C1 6B
 02 50 21 6A 84 7F 59 A9 5A 8F EA 5B 81 5B AC 6E
 11 D8 F5 AE 28 D3 C1 BB C1 0E 45 B0 DF 2B 9A F7
 EA E5 E1 C6 8F 20 DE B5 A8 D8 03 0D 33 B3 85 5D
 CF 3A C9 23 B2 7F BB 97 BD 26 AB AF C4 DF 91 73
 98 0C B4 9D D3 2E 61 AD 2F 30 D4 A7 D6 3D 24 40
 6D 28 3F 6F F1 5E FF 36 7D 18 F1 8B 2D 1C FD F3
 9C 71 C3 58 DE F1 87 AD 32 23 AA 94 C4 CE 44 A9
 83 4D A5 83 42 5A FC A1 52 3E 11 EE 7F F7 9A BD
 3A 08 03 97 76 4F 11 0E DC 3B 7B CB F7 4D 96 5F
 79 BB 24 3D 26 39 ED CA 2B 0B F0 B2 CA 90 3F 5E
 51 63 06 4D 29 BE 6D E6 BE 1B 6F EA 99 3A FF 50
 5E D8 53 4D B9 6D 0A 69 DA 64 33 15 B7 33 09 20
 66 19 89 A8 69 44 04 65 99 2A D4 BE CC C5 57 9F
 83 5F 02 9B 6E F7 29 E1 90 B9 61 65 85 6C C3 FC
 35 C7 6A 37 E2 B4 D6 F9 6A C2 9D 9F 66 09 82 CE
 47 EA AF 8C 63 38 32 E2 E9 13 06 1B 43 DA FB 0E
 C8 BE FA E5 1C AE 92 FB B7 FF 80 AE D6 8C F5 EB
 AC 93 95 AE 68 BE 7B 28 50 A4 57 D4 CE 98 89 A6
 D2 3D F8 2C 3C FF 9C 53 79 F7 71 6B 9B 06 E8 79
 F4 0E AC 5A 0B 7B 02 BD 87 8D 76 C8 0E 89 FB 07
 8D 08 DB 5C B4 76 45 A1 C4 B2 08 9B 2B 5D FD 7B
 A7 74 CD 6F 57 19 42 6C BA 87 0E 4D 27 7C 3C 4E
 B4 3C E9 4F CB 3A 5F AB 28 E8 06 50 F2 A6 4C A5
 F0 B3 94 DC AD 9C 81 16 05 E0 F7 A7 1E F8 82 43
 A2 68 71 57 60 FD 50 12 A9 6A 64 DA 4D 52 A6 CD
 0A 63 4E 9A 19 94 3C A1 8F 62 AF 18 B8 68 0A 89
 65 F9 C1 87 9B 57 26 25 68 6A 8F C4 FB E3 74 05
 81 0D 2A 99 C4 3F 0C 5C 32 37 4A 64 D8 C1 6D 3D
 B3 A7 D2 DB 38 FA 15 92 DD B5 FD 77 BE 02 D0 33
 A4 F0 55 BD D5 04 B0 F5 FB A5 EC FC C1 91 F9 F5
 7C 23 F9 15 43 54 D5 F5 06 A6 24 AA 92 F6 6F 37
 DB 35 A8 66 F8 05 18 DF B6 B8 84 76 79 DD 69 34
 25 81 93 68 87 D2 3B CA 36 BA 2F 1D 7D FF A5 1A
 F4 2C 8E 7D C9 1A 65 C7 CF CD E7 64 F2 C1 31 CE
 FD 59 93 3B 53 98 B5 AD F3 02 47 95 6A B9 6F 83
 91 4C 91 A5 02 E9 81 0B 4F 63 55 A2 29 5E FF F4
 F4 8D 01 16 13 93 FD 7D 19 AE 23 5C 1F E4 F7 86
 B2 8C 31 77 D5 30 C3 E9 26 81 AB CB DB BB 12 16
 77 3E 84 86 8C 6E 0F 04 F4 3C BB 3C 23 A5 E9 6E
 74 CE DB 4B C5 D6 E6 19 CD E1 2F 43 9F 1C B1 45
 04 8A 5F C7 A3 4C 73 5A E1 72 4B 8E 4E F0 BA A1
 19 8A CF E0 9A 22 8E A6 D3 6A F4 0E 17 74 32 4A
 2C 35 01 CB A2 36 57 43 89 99 A1 9A AC 73 8B 68
 B3 3C 54 BE 19 5B 39 2F C9 70 DC 9C BE D1 36 65
 59 45 07 C7 D1 BC 50 FB F0 81 5D 6F 1D 04 B0 BD
 70 8F 4E 8A 9F 00 E7 06 CA 4F 65 9D EF 81 35 DA
 C8 F5 BC 36 93 19 E2 35 C0 36 E4 42 37 EC B0 AC
 3A CE 80 09 0B 2E C5 EE A0 DF DB 7C 2A E7 92 06
 3F 7A 39 E1 5A 2B A5 84 07 D9 55 D7 72 65 32 18
 4D 52 4C FD 19 56 7E F9 49 A6 F7 FA 34 98 8D 7B
 94 26 39 EB FA 1E B9 AB E3 2F F8 1B 0B 2D E1 46
 65 09 FC C9 30 70 DE 53 74 12 FB B6 24 7E E6 A2
 E1 3F 82 01 EC A2 CB 0D 4A 04 23 9A 22 14 A8 75
 41 5B 55 B1 60 DA 5E 9C 48 77 83 4E C2 7D 46 D4
 9B 5A 83 4E 31 99 D2 BB 68 AF 6E 59 8A FD D8 87
 79 99 8E C7 0E C9 EE B6 5F 81 02 BA B1 08 49 3E
 4E E4 A9 E3 90 A0 57 78 E9 27 A5 AE E1 5A B2 24
 AE CA 95 88 CC B4 52 EF AD 53 61 10 D1 04 C8 0E
 73 7E B6 41 94 C9 75 20 AA EE 00 1B 62 56 8E 75
 29 C3 BC 73 DD 91 25 0A 05 66 33 9C C3 CB 8F DB
 E7 61 96 97 27 BD 05 9D 8E 2E 91 89 38 05 1E 73
 60 45 75 3A 80 EA B8 CA 38 DA 9C 07 ED C5 73 F7
 2B 4B DF C5 54 A9 81 9C E4 24 C8 EF 6B A9 BD 1E
 FC 45 10 7C 16 04 4E 21 F1 A4 BB AF AC 51 6C 1D
 C9 9C B1 1D 52 7C E6 5A 9D BD D1 7C 71 C3 66 19
 08 44 E1 90 1E 9E E5 98 EF 7F 86 89 85 A7 05 49
 DB A5 48 35 CC AD 33 0E 3E 41 E9 E4 E5 C0 B9 22
 2E 60 9F 9D 0F C1 A2 F1 35 9B 27 63 02 CB D6 DD
 E8 AF 80 BD 71 1A 39 39 77 A3 A4 1F 3D B4 56 16
 4A 3E 46 8D C1 68 8C E3 73 2D C5 1D 77 05 F2 D2
 DA E4 05 6B E7 B7 BE 6A CB 6F 0E 5C 49 1C F6 E4
 B6 08 F9 4A AB 22 9F 6A B7 31 3A 40 29 28 42 52
 3E 9C 87 B7 1B E9 41 E0 FE 16 45 E9 ED 63 DD 4E
 71 58 E7 F0 2E A9 AD 6C C1 30 54 E7 9E FE 91 5E
 2F 7E 6B 18 89 9D DD AB A8 54 16 F8 CE 89 AA 74
 B3 53 F2 E5 1B 2D 10 4A 6C B2 5C D9 D2 83 2E 8C
 C6 2E B9 26 5E DC 7D 2F 7A 7C 85 1E 96 68 C2 91
 8D EB FE 23 55 C9 7B BA 2A 07 29 F7 21 37 B3 39
 53 13 BA 79 3F 7F 5D D0 59 F9 1E 56 46 14 A1 0E
 D7 EC 82 2B 37 66 F7 BC 90 63 18 62 AC 22 CE A0
 1B 3F 2F 00 1A 06 07 DC 6C B6 89 D4 98 A0 8A 4A
 13 8D A8 02 93 DB 47 FF CA 8D 27 8B 5E B1 1B 50
 D7 F8 0D 7D 4C F0 C1 E3 66 BA 7A E0 9B 95 07 17
 F0 F9 C1 02 CC B5 B3 12 F0 A3 FB 6B 7B A4 3E 8D
 16 7F 75 4D 23 BE 51 2A 08 2E 34 B9 00 B8 49 63
 20 A4 77 DE 37 D9 6F E6 17 C8 19 F8 B4 10 28 62
 02 E3 6C 12 2E 78 E2 E3 80 6B E7 57 F3 99 66 E5
 25 B9 0B A5 70 9C D4 6D 1C 5E 10 B6 40 E8 36 3E
 F6 85 99 8F 99 BC E4 EA 0F BC B3 2B 95 E7 CD 20
 84 4B B8 81 A4 4D 57 2A 34 42 CE 17 85 BA 45 42
 B5 51 DB 6E 4C 1E 80 FB 26 FE 85 81 CA F7 10 C1
 DF 2F 2C 7A A5 F6 8D 30 01 C7 24 F6 7F 1E 22 32
 CE D0 F6 FB C3 36 F5 45 51 17 B1 CD 5E 43 28 A9
 99 BF 48 DB 6B A6 38 94 85 EE 73 77 DA 9B A6 06
 BA CA AC 02 EF D2 C2 CA 1C F8 56 1C 3D 5A 54 5A
 E4 7C 55 C8 FD EA D2 3E 14 55 E8 C9 E2 85 30 D8
 18 B1 B9 B2 CA EE 43 C5 D1 14 88 E6 A0 B1 99 61
 61 1D 67 02 DD DC EA 33 2E 83 B1 94 34 68 E6 FE
 CE 39 D1 46 AF 5D 6D 88 A4 CB 9B 20 5A 4B 20 15
 E1 58 89 49 1A 07 9A 9C 4E 33 30 5E 99 5B 93 70
 B7 B1 70 41 BE 5F 35 8B E2 3C 62 37 70 68 9E CA
 16 55 6F AE E4 C5 9F 5A 63 42 07 F0 0F 84 05 F6
 33 C0 DB 4B 2F 67 3E 03 0F 8B 2D ED E0 2F 69 DE
 82 39 A5 7F 44 1C 22 59 D8 37 1B A5 C3 4B C7 9B
 58 81 3F 44 79 14 F7 42 C5 59 51 5A 6A 55 48 83
 15 76 25 48 1E B0 8C D0 07 2C 61 00 70 F9 49 74
 80 F7 EB C1 66 30 3C DC 72 F2 FB 37 89 42 DD 56
 EF 1E DC 3B AD 05 24 3C 44 E4 18 DC B7 6A 7A 42
 20 91 4C 1E 15 36 4B 92 17 ED 67 34 32 90 A6 EF
 ED 9B E7 5A 8B 9C 67 0D 92 D6 23 8D 08 A4 A5 F1
 73 0C 38 BD 6A BC D3 A1 69 9E 52 A9 82 CA B5 D8
 4C 57 18 AC 0C A1 06 ED D5 FD E2 1A 7D 36 C9 93
 F0 17 26 82 67 EE 7E 89 A5 D0 E0 D0 63 AF 6F 3D
 21 BA 74 4B B1 E2 94 49 0E 26 44 88 DA 43 5C 9D
 C3 43 F7 22 6E 16 A5 5C 28 B6 A5 6E B4 C2 41 88
 50 DF 90 4C 9A 5D 36 C6 6D DC EF F8 2E 5F C5 B7
 E7 4D 64 06 21 16 62 71 F2 F4 C7 F0 05 6B 0B E8
 AC 93 9B F6 22 F9 7C EE 03 3A CE 1A CA 7E E4 C5
 16 D9 D0 39 75 A4 34 8D 0E B3 D9 D1 3B 51 E2 BE
 F5 5B 85 1E 1D 48 7D 3A A8 44 1F 82 D7 43 67 FB
 9C 01 AE 63 74 AB 5A DF 6B C0 63 86 D3 BD 86 9D
 0A DC 37 DD 9C 9A E8 29 27 C7 8B D0 0B BA 08 ED
 AC 14 07 A1 B4 85 D0 DB 94 22 0E 72 9C B6 5B 24
 B3 90 78 85 DE 00 53 14 21 2E 86 99 03 F4 D3 10
 D6 8A D7 6C 73 F1 EA 5B 6E 22 9D 59 67 10 8E 51
 A7 21 1E B8 3B 91 34 53 F3 7C A1 F3 B8 90 D6 D5
 FE 27 E8 91 5E 07 17 E5 89 48 5B 40 4F 02 DB 1C
 0F C1 70 F5 7B 11 FA 4E 46 81 26 3A 51 93 63 7F
 38 A2 D4 B9 60 1D 61 04 64 79 2B FA 84 96 D1 2A
 20 76 C8 BA EA 75 27 2F B5 EC B3 6B F1 EC 48 D0
 0F 35 39 C2 03 06 14 65 40 09 6A FB 4D 5F F7 D7
 02 84 4A 1F C7 96 35 B1 76 E9 00 9B B5 DF CB 0B
 32 67 7A 09 72 0B 9C 66 A9 3A 8F 60 B8 31 11 94
 63 6A 09 24 43 01 BF 50 00 9D 31 09 26 80 01 94
 B3 32 C6 35 42 DD AC 49 DE D3 A8 AD 10 D0 74 47
 30 07 4A FA C4 A4 2C B2 12 B1 13 E7 7A 7A 0C A5
 0B 1D 45 D8 C6 DD 43 08 67 3A E3 8C CE FA 5A EB
 29 8F 92 2E 72 99 F9 37 5D E2 92 8B 8B 54 43 30
 B5 38 56 97 CD F0 94 1F 10 B0 8D 34 71 37 22 94
 81 78 20 04 D0 9B 6A D4 DA A9 45 BD 23 F5 70 51
 D9 F8 26 6D D9 A1 F6 22 D3 0C DA F6 D0 F6 19 07
 41 9A 3B 7A D3 85 67 5A 26 67 22 3A C2 D9 99 81
 E0 85 27 CC 0A 89 26 98 B8 28 F1 06 B8 F5 BE A0
 50 22 27 E1 27 07 36 10 A2 3C 68 58 09 4D CF 4E
 46 6B DC 31 64 74 80 A0 B1 C8 4C D8 54 CD D1 20
 BE 05 6B C0 E3 0D 32 22 3F E2 F7 5D F6 75 C9 DA
 22 13 27 F9 48 5E 3E 3B 70 86 3A C6 3E FF 1A 44
 68 80 C2 35 2C 89 1C 7F 2E 28 CA 3D 5F D0 DB E8
 A6 4B 27 70 94 12 12 A0 E9 B4 CB C2 DB BF 87 21
 CB 7F 66 8A 5C 51 39 90 0E 41 4E B7 4F 28 F8 6A
 EF 7D 1F 17 A8 F5 8D 5F F0 BC 6E E9 7D E2 1B C4
 15 37 0A FE EA 61 3C 14 B0 7B F2 16 1E 6C 61 1C
 F7 03 DB 5B A0 22 76 20 19 CB D3 11 F8 66 8A CE
 99 90 DB BB 49 D9 62 CE B1 3A 4C 85 F3 80 F0 C2
 87 00 CB A3 9E 10 2A 30 2A 8E 8E C9 AB F5 96 7B
 37 10 BE AB 8C 3B 54 87 A7 7E 6C B1 72 CB B8 96
 08 C5 C4 71 0F 39 7D 66 AC 9D C1 87 EF 70 5E B0
 CF 81 4F 6B 47 64 83 73 D2 42 0C 96 85 E9 94 6F
 DF F5 1D A3 30 6D F0 4A 49 F6 AF 30 FC AD F0 D4
 DF C3 4D 1F 88 D7 2B 0C 22 69 70 17 51 C0 1A 5F
 17 E2 3B BE 4E BE F7 4F 34 FD 4D 8A A7 40 B3 70
 93 4B 1A 2B 24 32 A5 AC CA 6A E5 89 C8 B4 3E 16
 EA 64 E4 FF DB 38 AA 4B 13 F5 8D 9A EE 74 89 97
 B3 33 13 94 5F 7C D0 16 38 EF 4A 0E D8 33 43 4A
 99 4A DA C9 03 45 B7 53 58 C5 E6 B8 DC C9 BD 90
 DA 03 1F 88 D4 E7 1F B4 1B 4D E1 23 57 46 F6 D3
 16 43 20 C3 D5 3F 74 76 90 F2 98 EB 89 4E 0A 18
 A4 D9 AE 60 88 28 5D B9 BF 7C 96 0A D8 84 6D 68
 2C 32 38 4C 03 6A 01 DD AC 1C D0 18 67 17 73 79
 62 EA C2 58 6B B1 EF C3 02 15 97 6F 86 41 67 15
 42 D4 B0 EB CC A5 49 07 EF 86 FD 05 36 F7 D0 77
 1D 27 EF 14 95 19 04 1E 13 F3 B5 D5 56 50 89 BB
 6E C8 CF FE 92 D4 81 7C AF 29 44 76 03 E6 AB CE
 20 13 3B 55 C7 82 AF CA C1 40 57 2B 3A E3 2C E2
 C1 92 D3 7A 4A E1 A2 D0 27 E8 52 9D 20 AF BF A0
 78 CD 2F BD 95 4B 5D B0 0F 40 68 B9 FB 62 EA 86
 73 CA 1F 08 DB C9 9B BA 35 2C F3 AA 6E 99 28 30
 AC 87 5E DB 1D 03 19 47 95 AB 9D 5C DA D1 BA 31
 2C 6B DB BE 9D ED 35 DD 75 BA BE BB FF 22 1C 14
 5B 60 4F FF 67 00 BB C0 3D EE B1 A5 70 A4 5C 2C
 92 ED 99 1F 9F 71 C0 01 01 6A 2A 45 CE 21 BD 9F
 83 75 3B BC F3 BB A7 DA F6 AF 5E 1A 6E D5 70 8B
 3E E9 97 8A A4 E3 F8 41 65 E1 D7 06 71 D0 79 87
 9A 3C 78 CE CE 4C AB D2 57 E1 03 1C 75 1C E4 1C
 74 65 F9 59 7D BE 8E 4B B9 19 51 7F 0E F9 3C F1
 90 5F CB 3D 28 84 65 C1 B4 78 CC 7B 02 DC 5A 06
 4E 33 AE 02 B9 F4 67 0C A2 5A 3E B2 80 CD 18 FD
 49 92 59 FD A0 61 F7 A9 35 0B 4F F1 45 0C 6E 47
 2D 55 1D 08 C4 C1 EF 62 9F 51 7C D8 F8 81 66 B8
 1A BE 1F 46 53 64 B7 60 C9 5C 4E 4F EB 20 2D 6C
 1E 88 7A 40 18 CD CB 05 B7 63 6D 0F 8A D4 86 5C
 FE 56 80 12 71 89 4F 13 4A 24 3B 47 3F CE AC A4
 DD 0A B9 AA 54 13 E2 EA A0 AE 0E 65 81 A8 DB E2
 17 A8 A7 1F 47 CE 2A 0B C4 8A 40 6D 43 31 EE 20
 C4 B0 6F 37 4A 49 E4 20 43 CC 6E 4B C1 F8 07 57
 19 99 FF 61 03 FB A6 FD 60 84 DB 3C 77 C7 06 AF
 30 AD 8D D7 8C 7B 0E EF 99 B7 39 B3 D3 15 77 3F
 13 AB 08 18 F2 66 03 97 18 0D 64 B0 80 FE 15 D8
 4E 48 23 74 24 16 CB 94 B1 F8 EA 95 B6 9C A1 69
 23 79 E5 6A 4F 1E AB 80 F2 06 BE B9 EE D6 FB DF
 25 A3 29 30 D1 94 09 91 CE 57 9D 0B E2 57 6F 1E
 19 C8 CF 71 A0 7B A7 E8 66 57 FF 54 70 4D D2 80
 9A 07 50 C1 44 8D 05 17 AB 7E DC F9 58 21 AC 0F
 F2 CD CE 4A B2 5A 29 55 0D 10 E2 CC 38 A6 15 F3
 9F D6 5D AF D8 D3 59 9E 79 48 41 FB 2E 54 20 1A
 B8 5E 78 0A 4E 18 D0 EC 5E 72 ED 3E 68 5C 56 73
 2C 9B 89 88 3A D1 D9 F3 00 AA 8D 0B BC 5F 73 82
 86 DB 1E FA F9 75 97 F6 16 54 5B FF CA D1 DA 6B
 86 F6 35 F4 03 37 C3 53 89 15 7B 17 29 F4 52 DA
 79 64 70 94 BA 47 83 7B 0F AC 22 C8 46 90 96 A9
 47 B1 F1 F2 AC 1D C5 1D 89 E9 0C C4 CC D4 AB 24
 EA 26 7E 81 5E 1E 1F 52 ED 9B E2 F4 77 80 EA B9
 90 25 50 C2 0B CD 6A FD E7 59 02 29 51 4A 95 CF
 93 37 EC 77 A1 A2 C2 A9 0F 54 47 88 CC 81 38 E3
 3E 03 E9 1F 7B 5C 34 AD AC CA 32 02 C5 97 AE 58
 D3 1D A7 1E 59 17 40 2F 65 9E E7 1B AD 4B DE F7
 53 C5 A0 25 EF EE 8E 91 B3 51 E2 00 DC 55 12 96
 F3 3D 41 9F A1 64 67 56 F0 B9 03 6B 31 9A 34 8B
 30 A6 AF 2C 77 06 E5 F2 18 00 84 01 EF 5A E5 70
 CB 81 AD 62 FD 9F 1F F4 4D 44 0A D3 DB B5 BE 44
 5F 6D EC BC A1 2C 58 DD 5E 61 0C 2A DF EE 70 7B
 3A B7 B6 E5 17 48 7F 4B E2 B0 90 17 98 DA F7 FA
 DB 88 37 40 33 A0 95 03 6F 46 24 EB 57 C3 1A 70
 51 C5 03 9E 10 48 A7 D1 E6 41 A5 C4 73 77 67 64
 8B 2D 6D CF 31 79 57 08 04 EB 09 1E 8C 96 82 6A
 BC 0D 5F AA B3 E5 BF 49 62 44 E6 6D E5 C3 B3 32
 DC 6B BE 3D E0 0D 08 41 C3 AD 08 7E F6 8D D6 9B
 23 DB 8F C4 FE 56 05 AE D1 7D E0 72 D4 95 B6 60
 5C 15 4C EB E5 ED 31 AD 09 A2 FA EF 96 DC 03 A0
 F0 AE 1F 1E C4 52 A5 86 E4 68 8B FB B8 97 BA 30
 7B 9F 6F 82 68 25 E8 A8 8A E6 CD 07 22 3E 39 96
 58 38 D3 6A 41 1E 5E A4 A0 F9 5C 08 83 7E 14 2F
 1C EA 43 3C 7A DE 8F A3 4B 7F 3E 04 FB AC D7 40
 49 B4 16 C1 A4 3E AA D0 F7 CD 05 16 9D D1 8B 89
 2A D5 33 64 39 D7 21 A3 01 01 68 B8 1B 3F 28 E5
 04 73 F1 A2 BF D9 46 3A 64 F6 A3 45 41 07 99 C0
 1E 57 D5 25 7F 1A BC 24 20 A9 55 CC 22 25 90 07
 9D 5E D1 AE 47 C0 DF 6D 67 71 19 DB AD 2D CC CB
 F4 89 78 B3 7B 2E 0F CA B1 E4 DB AC 91 F9 F1 7E
 73 DC A2 06 EF CD 67 E1 5F 89 90 14 96 EF ED 7E
 D1 8C BE 16 F1 DA E1 E6 EB 10 21 9D 9A BA C7 75
 20 50 48 74 33 91 4C D9 86 AF 8B 18 9A 51 4C A8
 A2 E7 DB 45 DE 74 E5 88 80 99 E2 C7 64 EC 42 09
 6A 67 95 FE 9F CF EB 34 0A 75 21 1E 5F 46 13 D6
 3D 33 BA D5 EE EA F8 10 BC EF 73 D1 09 78 73 A5
 6D 88 C8 EA 3A 12 40 C9 07 40 9A 5B FA 69 55 82
 94 9E 09 E5 8B E9 E4 9C B7 C3 79 C8 81 36 CC 96
 C5 DD 7F 60 19 48 1D 95 A3 42 BB 0E 31 C5 54 05
 4A 63 68 7A B2 1F 56 2B C7 C6 C1 5D E5 43 54 AF
 57 A9 E9 36 28 B0 1E F0 48 91 65 FA 7C 05 7D 4F
 BA 8F FE 83 B0 79 90 D9 A8 ED 57 7E 18 0F FD 1C
 C8 DB 81 54 21 8B 54 DF 42 A9 B0 62 45 05 55 22
 73 CD 72 CC A6 29 9B 70 E4 1D EF 14 10 55 99 C6
 74 14 8E 6D 18 4C 6A 97 69 0B 6F D9 D6 75 78 59
 95 D0 D0 8E C2 10 6F 41 04 BB B8 D7 F0 89 65 7D
 D7 33 DA 38 E2 32 5C 38 34 D0 3C D6 23 0D B2 41
 CB 15 A9 DE D5 EF 76 B1 5B A2 AA E9 A8 95 98 95
 B0 E3 27 2B D5 7C 91 A8 CB E9 0C A0 D2 A1 62 A8
 BD 5A B7 4A 8D 9F BD E9 A9 B3 9B 52 DE 7A 79 5A
 EA 0D F5 71 E6 F8 FC C1 43 0B FE D2 C6 44 35 EA
 8B D4 FD 19 DD 2A 53 7D BB B5 DE 86 90 2F 7A 52
 E5 E4 A7 95 B4 D4 4E 2F DC 8F 65 1E 10 F1 E4 38
 6C 7A 90 8E 63 CC 06 E6 D0 81 27 75 BA 15 E0 D3
 AF 20 DD 66 22 8A 9D A7 16 46 B2 96 B1 56 F2 12
 00 49 05 53 5B 4F 8A 2C 4C B2 CC 04 9C 56 89 48
 93 2C C1 72 B3 A0 1D 2F 95 EA 83 5C 20 F1 AF 6D
 EB 6E F7 55 2E F8 C5 AC EF FA C3 91 18 3E 2F 95
 A3 F2 C9 57 BC CE F2 2E FE 92 39 4E A1 3C EC 09
 BD 11 81 7B 01 A8 DC A7 55 95 F2 64 40 F7 3B 85
 24 DA E5 E0 BD 19 21 02 97 46 2A 4B D9 09 29 0F
 61 19 90 72 25 09 FC F4 DD 7F A7 FB 2E 45 7D 0D
 FD 69 43 09 AF 30 1C DE 06 69 4D A2 C0 BB EC 7E
 D3 A9 C6 EE 9E 88 64 15 13 95 F3 1B E5 F1 72 01
 5C 3A 45 4D 36 2B 7A BE 41 6B A5 F4 6F 22 BA 2F
 0D A4 80 3A 1E EF 68 3A D1 0D 18 56 AC 8F F8 85
 4F 37 A9 13 9D BF 40 31 B3 AE F7 8D 15 97 E0 C3
 CF 0F 0E 5A 97 9F FE 09 68 B7 B5 E0 BE 63 35 C2
 52 E1 0C 35 32 F2 1B 4C 58 F2 FC 25 EC 61 F5 B2
 B5 83 9D 65 FA 6F 39 13 68 5F 11 0B 97 C5 7C 73
 6E 76 E5 33 9F 10 E8 C8 62 37 1B AB D2 EC 11 5D
 72 6C 4E 0B 13 DE 26 CE 4F A5 B0 87 E6 52 68 D1
 BC 52 B5 27 E6 29 F5 31 87 73 FC DE 9C 5F 2E 58
 1E C3 39 96 E5 2B F6 34 65 B0 BD 4F 61 C3 5C A6
 4D FB 06 FE 67 AB 9A A8 6E 6C 6F 94 84 79 F6 97
 79 55 CF 30 C9 9C F2 DE AA DB F9 F7 9F E9 91 D4
 11 71 8D C5 55 3C 59 8A 2A 52 63 51 3A 29 3A 68
 8E 9D 18 9C 92 A8 0B 5A 3E EE 4E E3 70 71 D2 6B
 CB 8F 24 73 ED 60 19 6E AE 4E F2 42 A4 A9 B0 BC
 90 E1 0E 68 DF B0 24 6A 89 FC 64 C4 0F 40 9A 3A
 BE 4C 5D 2A A9 73 61 68 26 9A CF EA 3B BE D9 91
 1C 05 22 6D F3 F3 E8 8B CC 7C D0 71 30 79 B4 7C
 3F 2A 59 93 4D CB 62 B9 FC 19 0E D2 4A 2B 2A B6
 67 F7 CF C0 39 68 60 6A 1F 97 7C F9 42 67 14 2A
 7F BD B4 B3 5D 29 5F EA 90 53 70 94 DC DC B6 25
 D2 A5 3E 21 92 FD 8C F5 E2 4F 09 39 28 00 C2 01
 8D BB 88 A7 F3 BC 15 98 C2 F7 E0 91 5E 2B 81 1F
 2F 80 83 E9 C9 06 44 5F CD 03 83 20 15 1C 3A A1
 53 36 F1 D1 5A 66 99 95 A4 54 EF AF C3 21 DD 63
 3E B3 19 DC D1 6F ED B8 2F 05 A3 8C 32 97 7D 47
 33 96 41 47 D7 86 E5 4E 61 EB 34 F8 31 35 91 0C
 6C B7 65 4B 0A 47 D5 22 D5 B5 43 27 F5 81 FB DC
 32 2E 0E 33 2F 70 8A 47 06 49 67 7C 73 80 EA FA
 11 DB 6A D4 AA 9E F7 5E 43 0B 26 C1 F0 94 E0 AA
 E4 C1 E4 EA 9E 8F B1 FD CE E5 89 8D EF 0D 5A 9C
 A8 D2 BF 0A 45 E2 F9 87 88 75 40 E2 5E A8 60 65
 07 CC 78 0C DE E7 85 66 EE 8D A3 C1 D4 EE 9D 61
 0E D3 07 7D 79 DA 1D 73 B7 20 09 61 59 DC 04 DD
 8D 57 71 B9 6A 96 0E 82 93 81 E6 92 F1 A1 B7 9B
 04 76 97 25 1A 5D 02 02 C0 02 56 81 CA 2B 75 8E
 0F 4D 56 AA EC 9F E5 D7 2F 9E 1A 17 9A E0 DB 24
 05 27 E4 B4 E9 09 1E 25 AA 6A B1 12 92 11 9A 46
 73 4E CC 55 54 C0 07 4A EA 95 28 3D C6 0E 9F 0C
 9B 6F 7D ED B1 72 AC 72 8D 63 57 81 6B 97 9F DD
 5E 58 FE 93 0D 77 4C 87 8C 84 83 4B D8 BF C8 B6
 21 79 05 79 59 2A 15 EB B9 F6 BF 40 10 76 42 8C
 81 FF 75 1E C2 7E F8 04 7A C5 16 95 0D 0D E4 19
 BB 36 CA 53 5D B2 9C C4 7C F7 24 74 A8 07 0E 78
 4A 72 E1 2C 58 EF 50 A4 6C CC 10 D6 84 E8 1A E8
 F2 9E 3C FB E1 88 D5 D1 94 2C 8A 78 FF 6A AA F4
 BB 2B CB 30 D3 87 7A 00 32 C3 BE CD 32 C5 E7 C6
 42 F2 D9 65 91 43 33 94 0B 19 92 E6 07 07 F2 39
 0B 7F E1 01 95 F0 77 D5 B5 DF D4 6C 7D 65 07 46
 3B F4 4B 30 08 49 4E DF 94 55 BE FA 31 40 E6 ED
 BB C7 05 9C FB CA E5 74 70 E2 14 A5 E6 52 22 E4
 55 AD F1 C5 AB CE 9F FD 6B B7 17 4C C4 1C CB ED
 1F E9 D8 1B 93 0D 9E 44 D8 E5 C1 D5 B1 45 34 9B
 35 7D F3 C9 81 EB C0 08 33 2C 12 D7 D5 E8 6D E5
 BB D8 03 07 9B 7C 58 BC 6B B8 EC E5 C7 30 57 17
 72 B1 16 20 41 53 78 9B 0B 4B EF 50 0B 39 8B 3A
 79 65 84 5B 2A 3D C4 29 35 1C 27 4A CB 81 3F 91
 DB 07 E5 30 52 6C 69 10 32 77 50 30 B3 DB 0E 97
 17 03 AC 26 F5 5A 4B BE 3A 90 AB E2 39 5C 48 63
 6D 31 D6 FB E0 67 C4 55 1C 5F 0C 89 46 F1 14 B4
 96 E6 75 62 22 67 02 27 6E BC 69 62 C3 74 94 72
 C5 6E 44 D9 D9 A7 7C 42 E4 40 69 F3 39 BE E1 E3
 3C 61 D1 07 0A 9D 4E 08 95 CD 7D EA EF FC AD C1
 CE B5 D7 54 95 1D 15 FA A4 56 B0 44 B5 1A 0C 2B
 33 C3 70 DA 62 D1 5A 96 CA FA 58 BB F0 56 DD E4
 38 BA 75 77 C8 21 B5 C9 C4 F7 45 20 7A F5 6A 56
 A5 7D 14 51 67 25 F9 12 42 A8 99 85 C3 4D 21 5C
 23 D7 18 AF 05 A1 0D 9F D1 3F D7 6B B1 17 23 53
 F1 02 E3 A0 7E D7 D6 E4 6B 01 DB 3F 92 CF CE CD
 B6 5E 5B 76 29 E6 22 4A 9A DC 92 18 B6 37 2F 6E
 89 84 80 D3 B7 5B FD 8A 95 EA 8C D5 98 12 22 4C
 0C E4 CA 0D CC BB C8 81 2D 77 51 1B 6C D3 99 00
 D4 61 2F 6A 5C 40 7F 99 A0 6B BA 5D EF AA 7F A9
 39 4F 67 63 61 C0 47 31 FE BE EB 60 00 97 4F B7
 92 22 92 54 EA 7A A8 7C 38 8F 91 F2 7C 5A 7D 47
 BA 2D 83 98 D9 18 C7 6C 40 65 D0 A1 67 C3 4D 8C
 13 A6 90 12 24 A5 70 73 F6 A1 01 1F B5 7B B4 B4
 2D 06 84 6E 13 B3 EB 2D 50 10 F1 E4 AE 4C 5B A4
 58 C4 02 0A C5 26 84 F8 94 BB F2 3D EF E0 8F 34
 7A AE F7 B0 6B 01 8B 29 6C 9A DA AC EA 30 CC C2
 DE 9C BF C9 B5 09 92 49 49 67 C8 96 4F D6 F9 71
 A9 F3 1F 22 73 90 C1 CD 63 54 20 42 78 8A 77 CB
 F8 BB 48 79 5D 37 86 3C 0E 92 82 01 A8 59 FD 00
 1E 6B 9F 69 EE BA 74 80 F6 33 DB DC 5B 38 A8 CE
 CE 06 52 0E 67 4B A2 25 89 52 15 13 B2 89 41 B2
 13 D5 0C 2D 81 17 F9 9A CA C3 40 47 F0 6A 5C 19
 E8 4D 11 9B 4E 46 50 F7 CF 2C 71 A4 ED F5 B4 AA
 FC 95 C7 23 5D F2 38 98 F5 D5 03 D0 7E BF 09 BF
 B7 CF F2 6E E4 2A 61 80 C0 4B FA B8 8F 5F 3C C6
 78 37 79 25 1D 84 08 7D 2B EE E9 F0 80 CA 94 D8
 61 67 9D ED 86 55 65 5C 66 C4 F7 92 07 80 F6 51
 72 16 AF 5D 21 40 5E 37 10 7E CD 93 E5 A9 0C B3
 88 F6 E3 71 4B 6A 95 09 66 B7 67 2F 26 D7 D5 DF
 F1 FD 79 CB BF 31 2A 42 25 A4 9F 23 11 9B 86 B9
 2A 86 56 DA 38 4E A3 34 08 AB B4 A0 2D A1 E1 58
 F7 29 6D 6D 95 C0 E2 27 D2 64 8B 53 6F 9E ED E9
 13 86 0C E8 E6 43 48 9F BD FC 4B F9 08 AC CA 62
 CB 80 34 B5 E9 90 7F 08 1E 79 F1 02 F4 15 B5 CC
 C6 FF A8 AF B0 B9 74 6A 13 B6 D0 87 D0 D8 A5 AB
 88 87 6B 85 ED 7B D3 60 63 F0 C0 94 1B 5C F7 59
 98 98 B4 F6 04 A0 9D D1 6F AE D2 53 DF CA F3 F4
 FA C7 71 D8 FB E1 05 F2 AB 2D F7 46 03 D9 82 94
 08 64 EB 2A 59 FC 43 86 33 A1 74 E9 C1 CD 5A C2
 1F 19 93 9A 09 3B AF 02 66 B2 7A DB 4A 6E AB 4B
 B3 E0 C2 3C 79 6C 14 A6 F1 78 22 5D AA CC 91 E2
 BA 59 9A FA AC 21 89 EF 89 13 E5 39 5B DF BD FB
 8B 0A C2 B6 CF 2E C4 2C 5B 81 93 30 D5 95 2F E5
 A7 5D 09 CF 84 E7 68 03 A7 D8 67 2D 6D 05 62 DE
 45 48 90 D6 C0 93 B1 03 59 71 6F FB 9D F9 A3 6C
 45 1A E2 EC A6 F6 C9 19 21 80 E3 67 C2 A9 D3 1A
 DD A5 45 2D 5A 7D 78 71 A5 C6 19 D5 F4 22 EB AE
 D3 DB 0B 68 CD 75 7B 46 C3 93 8D AF 35 20 25 49
 C2 DB 61 B6 80 14 17 0A B4 B1 86 C1 35 01 06 91
 10 42 CF 46 D4 CD B2 22 F7 AE 50 D1 5A 19 CA 57
 46 E0 69 97 87 81 71 1D 20 DC E9 C1 3A B2 AA AF
 9D AD 62 75 CD 1D EA B9 1B 7F 6B 6B 62 DE ED 72
 2C 1C CA AD 17 32 2C 41 DF CE 96 D5 96 F9 08 6E
 E8 32 52 7B 6B C4 42 68 AE AA C2 DF C2 96 F3 5F
 F7 74 95 70 23 3E 22 07 85 07 89 14 BA 11 2C BB
 19 9B 25 99 CF 22 8F 9E 94 DB ED 76 1C D8 9C 32
 A3 0A B2 B9 FB C0 CF FD 0C 09 E5 AA 86 4C 05 CB
 14 B2 82 5A 0A C9 C3 A6 F5 29 29 9A 4E 9C 82 98
 AD 2B 9E EE 8F F6 CC 57 D9 53 62 7C 85 F7 96 14
 B1 C1 A9 2D 1F 20 77 B2 91 6F F1 4A FB 00 A1 AF
 DB 49 3D 18 5A F7 E4 96 56 ED 89 C7 93 1B 34 29
 E3 D3 0B 9D 7A B8 F8 05 EC 9B 9C 65 35 CB 3E 02
 ED 04 E9 30 71 C9 E4 44 E3 D2 B4 A1 78 9D 05 C0
 41 EB 86 BC 88 8C 08 90 37 30 52 67 2C 73 10 3F
 7B F2 FE C5 46 1C 90 59 AE 6B B4 F6 3F 06 A7 F4
 50 2C 7E 0A 87 C0 26 09 D8 78 C6 F9 0F A3 0F 05
 DE C8 D2 2B 52 98 E6 AB 51 DE 27 75 20 F1 D6 FD
 F0 53 AF FB B9 5D F6 B7 C2 70 FA 07 3A 61 C2 7F
 03 B7 50 D1 57 29 A8 AF 0B 19 AF A7 D6 75 78 31
 19 F6 76 A8 64 0B 58 73 D4 6D 05 E4 F6 DA 11 B4
 B1 C4 BB EB EB D2 19 56 AE 9C F3 6F 64 F0 DB E8
 AE A9 1A 0B 9B 69 89 BA A4 75 A9 EC 04 DC 73 BB
 29 4F 15 9D 7D E1 10 28 BD 95 48 12 4E 84 DF 70
 F0 D7 BA 71 CF 86 43 77 C2 E0 41 02 D7 B6 DE 2B
 29 43 CD 0A 49 EB AD AE 88 13 C5 9E 63 CA A8 79
 C6 B4 D3 E3 02 8D 21 B9 7F 28 D5 88 4D 12 37 1E
 C3 00 3B 31 06 6C B8 DA 5C B3 22 4D 3C 5F 11 F5
 EA 0A EF 42 0F 42 86 71 2A 29 6A DE F0 EC D1 3C
 3E 52 56 93 CB E2 68 A5 B1 C8 41 32 8B 10 C7 92
 ED 9F E4 BB 84 08 04 2B 84 0B 1C B1 0B 42 A8 8E
 A2 3E 6F F4 5E B7 D4 94 04 31 4B 5F CA B5 AC 37
 30 4E F6 27 73 55 C3 93 F3 E5 00 11 25 4A C0 FC
 34 C7 0B 61 AC 7F E5 0C B1 A9 24 95 70 E9 C2 BB
 CF 31 4D E8 B2 9C 1F D5 8E 2A 94 0B 50 51 03 57
 4F B2 BD 5A AD 57 DF FD 78 7C 57 B1 CF 59 AB 38
 01 2E 54 E5 4D 7B 24 C0 79 2D B7 13 0F CF DD 94
 18 5C 00 41 88 04 DA AB 07 BB 20 D6 81 57 A7 11
 DC B4 9A 24 50 99 13 6C 6C 78 F5 7F C9 98 07 F9
 C5 AF 94 6E BF E8 DB 6F 11 68 67 8C 77 47 C3 44
 7F 05 81 81 35 75 9A 45 74 D8 F7 2A B9 D4 E0 50
 7B AA 90 F3 A7 30 4A C0 F8 C6 45 3C D8 EB 8A F9
 03 FD 09 3A A7 86 21 D4 C3 FD 29 8A 70 81 8C 48
 9D F7 3B 17 44 07 43 5A A5 A8 FE FE 7A CC 25 97
 0E 0B EB C7 D2 D7 99 FD 57 21 CA 27 9F F1 CC 22
 0D 18 C0 2D 7F DF FF C1 FE 59 23 1C F4 73 D9 52
 86 14 AC 6A 03 84 2B 03 FE 21 23 F2 6B 9F 79 D5
 D6 64 73 FA DB F3 53 05 E0 5C 78 4A AB 7F C3 58
 91 A6 98 F6 A9 D9 E4 2B F9 1E 5D 53 E4 7A 2A 2E
 F7 6F 03 8A F9 EF 68 8C A3 5C 89 63 73 46 AC D0
 DE 66 EA 76 AD 32 1A 6C ED 21 34 EF 78 BC 8E 50
 00 71 4B 93 50 36 9B BC 81 18 23 59 0C 79 81 12
 4F F1 EB 91 79 8E 39 38 03 55 7D A8 29 47 BD 89
 D1 EE 88 0D 58 DD CD F4 76 3C 6B 1D 9C 6F 09 15
 5F F4 64 D4 3B 63 06 59 B5 0C 27 41 4A 35 CF 33
 AF 09 BF 1C 3F 93 A3 3D 22 05 08 A1 ED 77 BC 38
 98 27 DD E6 6B E6 91 18 21 07 3E AA 5B 11 EA 97
 29 A0 5D 73 50 A3 C2 2B B9 99 64 7E 6B 86 89 3C
 AB 24 07 35 AC 07 C6 13 C2 E8 FE DE 90 0E 16 CF
 E6 29 D3 66 8C DF EE 7D 1E AB 5F 55 B8 72 9B EC
 93 42 8A 8B 86 BD 31 24 A0 4D 5F D1 1F 2F E1 C8
 88 A5 8A BD 24 0A B5 B4 C5 0C 08 9C 46 F0 20 08
 51 03 4B FF 64 80 45 FD C0 E2 BE 2B 13 FB EC 41
 7C 08 72 5B 2A 54 E4 0F 75 B8 F8 93 CC 5C 17 A6
 C1 0F 50 6C A2 D9 AA EB 1F AB 64 59 E9 64 25 01
 9E D4 5D C9 47 4D 6C 1F 72 EB E8 18 E1 30 F1 90
 FE 63 74 43 09 DC D2 A5 F6 17 B1 7D F6 E8 00 7F
 02 F9 04 74 E9 80 7F B8 9F C5 8E F3 3E EC C8 71
 2E F9 03 47 20 BE 93 2C AE 7B AF 23 6D 9A EF BA
 29 CF FD 8D DD D5 68 33 6B 66 56 1C 94 D3 B9 59
 AC ED 4B 98 FF 2B E4 74 0D 3E C3 5B ED 7F CC C3
 7A FC BD C7 33 9C D5 DE 47 E8 0E 55 EF 93 9E E4
 7C 05 4D E4 39 77 30 6F 8B 3C BB 89 40 72 E6 5A
 58 F1 AE 67 98 8B C7 D5 88 BC 20 D8 0C FA 6D E7
 5D 64 CD 0E F6 74 77 1D D8 D2 A1 10 BA BB 8E ED
 8A B2 2B 1A B0 9A 16 CC CB 6D 82 CE B4 B3 67 AA
 84 8E E2 70 F8 DA E7 6C 55 67 71 6A 61 D5 61 F4
 66 CF F8 A4 E3 B0 0F 5D C6 37 0F FE 42 56 B0 0E
 F8 D6 03 5D 2D C0 D5 FC 72 7A 8A 57 1A 53 FF AF
 AB A2 F6 64 F4 9B FF E3 C5 FE ED 25 9D 15 F2 1B
 3D 4F 15 7E 88 3A 88 4C 84 04 38 46 72 71 E2 74
 5C 0C E0 D4 E7 6E 06 51 0F E2 13 DD 89 5C 6B BE
 6E 3C B6 29 28 A8 F3 A1 6A CF DC AA C3 A6 2A 52
 C2 FA E0 B7 EA 37 18 E6 7C 4C 40 E7 20 47 71 18
 E0 33 16 5D 6B FC 85 19 0C D5 40 9D 2E F4 95 88
 AD F6 C6 E3 22 74 08 BC D7 40 E0 99 8D C5 1D FC
 35 97 56 30 AA 18 4B 7E F7 E4 A4 04 E2 C8 01 5F
 3F 2C CD B1 AC 6C EB C9 22 13 DA 67 5D A2 F5 20
 55 C9 6D F8 39 8B 16 FF 88 EF 88 B4 7B A2 0A 9E
 9A 4A 51 20 37 A2 AC A2 F0 3F DE 27 1D 28 12 2F
 0F E5 06 F5 42 CB 35 A0 3C 77 62 A5 E9 38 3D EB
 ED 1A 5A 74 55 0A CC 18 3E C7 68 57 D0 CC 38 80
 35 84 37 64 8F E1 7E 31 04 1B EE AF BD A6 AB 3D
 A5 67 9B 0E 01 40 B1 AC F4 AD 1B 01 BE 9B CC 17
 20 92 82 BC 97 1E A5 22 97 D2 8D 65 80 D7 64 56
 49 D4 CE 81 CB 38 5C AF 5E 3B 77 B2 EF 45 A2 3C
 3C 80 49 1B D0 9B CB 69 81 23 4C EF 5E 5F BE 03
 BC DE 14 CF 17 21 2A 5B 37 F5 B2 C0 28 29 7C CB
 00 27 16 A6 7E 09 31 99 F4 F9 06 CC 58 CF E9 D0
 A1 6A 06 8B 94 1B FB E4 B8 2F CD FA 58 DE 42 9C
 50 7E FD 57 F4 2B FA 5B 89 B7 4D 24 09 48 03 10
 62 04 F4 00 A8 66 3F F1 7B 3C 5E AA 78 7A DE 69
 C5 BC EE 41 9C CC 7E 30 69 58 15 1A 02 50 34 26
 1B 21 60 ED 38 19 43 15 38 AE 83 C4 24 FF 3F 70
 58 66 25 2B F1 E5 BA 9E 9E 8B 93 F9 A8 E7 0B B7
 71 2E 6C DC 30 43 81 85 49 EE 0C A4 B2 70 AE 96
 40 65 BC 1E FE 9D 36 6E 8C 63 75 36 3A CA 1E 88
 7B F9 3C 94 FC 97 CD F7 EC AD EB 0A E1 DA 94 FB
 1B DB 4E B3 B0 66 44 20 8D 07 8C D9 85 C4 92 7A
 AB 17 D4 36 36 98 AD 86 ED 9F F8 63 0A 75 17 EC
 AC E0 BC 37 D2 49 F0 6F E3 4E 5B 0E 6B 27 DE AD
 C3 9E B9 84 A9 69 BA 0F 68 40 AA 06 72 37 C8 37
 95 C5 B5 E4 2C EB 3E 5E 53 EC 62 38 53 E2 5A 64
 10 B1 95 A5 56 53 24 D8 C1 B8 1C 38 73 DC D3 4B
 BC 8A AF 70 80 A9 DF A6 DB C6 E6 AE C7 EB 94 FD
 5C 48 94 06 9E FF DC C1 C8 E8 B2 05 FE 07 94 2E
 12 26 DF 18 50 99 0C 90 47 D4 A6 38 32 5A 4D F5
 F0 F2 54 7C 91 0D 13 5A CF 43 E5 79 A7 EE ED 05
 B6 10 56 FD B2 48 EC 6C 76 27 D8 1F 12 03 83 E6
 A5 C5 80 D0 81 21 A5 EA 46 06 D9 CA DC DF 48 A8
 6C 76 2B 9A 34 09 95 C5 EC 3F 74 B6 03 F4 07 32
 BD 34 88 AF C8 A2 38 E6 C9 89 8D 6B 49 B3 81 EB
 84 59 1E ED 08 27 F2 79 C7 A6 C5 53 B0 4D 3D 53
 3D DF 56 D0 A0 DB 5F AE 21 0D EB 32 48 FD EC 79
 2B 0E E2 DE 2F E3 D9 F1 3D 51 EE BD A1 FA 23 D4
 DE 13 A0 30 F8 13 A3 8F 68 E4 4A CC DD 9B A6 AB
 C3 61 DF 48 ED 6D 12 25 5A 0C 80 7C 90 8B F2 57
 F2 9A 5E 36 15 39 6A 6D A3 F1 85 24 22 7E C4 31
 B4 11 B3 8B C7 1C 2C 8A CA A6 B9 D0 0D 5C CD 22
 96 C9 8E CA F6 0A A5 C3 A9 A7 B2 DE CA 98 C9 0C
 20 2D A4 9A 1A 44 6C 84 C4 EA 6E 8D 57 55 3F AB
 88 93 48 DC B1 24 D7 19 E0 9B 20 1C 21 01 C5 B8
 FA 23 C1 AE A0 48 92 CC 11 D6 B9 D9 A1 DB AE 77
 3F ED EF 8B 5A FC 6D 9D 19 07 EB 86 AE 1C 10 C7
 62 3B D1 39 B5 4E A5 DB 1C D8 6D 0C 84 9A 44 D3
 B0 8C 76 56 E5 8F 78 8E 2D 65 8F 92 9D B5 41 C9
 C0 1A FE F9 6F A6 7B CA 14 AE 76 95 95 37 5F 0D
 2D 72 DB CF 4D 22 DD 6A D5 C5 BC E4 7C 69 A4 F7
 C1 3D 94 12 2A D3 58 74 98 5A 58 BD B4 C3 C1 93
 8B 92 2F 58 00 C6 99 DB E7 A0 2F 3E 67 BD A7 3B
 E2 B8 5D 61 F5 3A 42 A7 70 D8 5A 32 C3 24 1A 2D
 D7 29 92 CD 1F 99 3F 45 DF AC D8 AA 5A 21 62 C7
 AF DD 3C 02 5D C7 90 55 32 63 9D D1 C7 F3 C2 83
 6B EF 69 DE EE EC 39 E9 4B 78 F2 1E 13 5F 11 94
 7A A9 B2 4D B0 D4 70 AE 7E 6B D6 6D 18 30 5E 81
 20 DE E3 3A F5 D0 FC D2 BC 46 ED FA 02 95 14 CD
 59 4C B5 48 96 74 47 AE 18 E4 72 48 E7 7A 26 C6
 AE A2 B0 CE 49 1F 06 7A 70 5C 82 B5 E4 BA 1B 10
 17 82 EB 50 C0 49 6E 10 C8 2D EE 89 99 3B 4E B8
 B7 DB 3C A6 83 FA 55 FF C5 33 28 84 62 1A D8 3A
 BE C2 D2 B0 1B 1D 65 C9 C5 CF 3C C0 2F 95 33 DF
 5D 1B 7E EB AE 34 67 49 98 5E 84 C9 10 7A 9B AF
 AF 2B 43 07 D3 6B 28 49 D4 43 BE F4 A1 55 6A 7B
 AF DA 8E F0 4B D6 E6 6F B4 C4 17 ED CB 24 E5 F1
 7A 1A C6 B6 FA BE E3 40 51 53 69 78 7E D4 C6 C9
 C3 48 C6 6C 18 80 A1 51 30 C2 38 E6 09 AE 29 16
 D7 72 A4 96 AF A3 AF B9 34 0B 8F 27 9C BF 9F 5E
 AF F8 E3 B5 10 88 89 72 B5 5E 08 EA 2A FE B3 95
 5F 22 FA 20 D6 8C 7E 47 31 A8 6E CE 6B B5 BE 4B
 0F BC A1 27 77 BA 38 D6 3D 0C 5B FD 84 42 9A 21
 96 97 32 FC 44 DE FD C7 C6 B4 24 51 59 30 FA AE
 BC E2 68 83 86 BA 68 63 51 A6 A2 C8 1F 2E AC A5
 AD 83 13 2A 84 4A 16 47 1C A4 82 C8 97 A7 9F 58
 6A CF 5C 78 4E A7 A0 00 72 18 B3 89 4F 03 C2 91
 FB 01 74 21 96 73 3C 3B 80 CF 75 3D 4E EB CC FA
 F0 C9 E7 D5 A9 A6 A6 ED BD 75 B7 35 F6 A3 C1 42
 26 E5 C5 0B 55 5F E1 B8 8A 8A 98 F6 8E 76 F9 DC
 BD 92 CE 5C F4 2C B1 A6 9E 8E BE AE 51 04 BE BD
 94 0B A4 9F 11 FA 20 8E 81 67 D8 6F 86 8B 76 39
 49 9C 14 5E AF D9 6B 4B 76 8B 91 54 B3 85 57 5F
 99 3F 7E C7 36 A4 B3 63 15 AE 30 97 F4 22 70 30
 32 B7 1C A3 68 78 0D 4A BA F8 48 66 4E CE 93 2D
 59 7B 2C C9 3E 3A E6 06 9E A8 36 F4 56 B2 9A 25
 6F DA BA 30 23 31 64 73 4F 93 65 61 18 FA BE 72
 78 20 21 F5 D2 8C 99 44 0C C3 6A 80 C8 F9 EE 1F
 D2 74 7C E8 EE 5C 55 BD DF 9F D8 97 63 25 60 41
 51 C8 EC 77 F8 46 80 05 39 D7 5D B7 E5 BA 67 07
 D6 32 0E 95 D3 0D 15 0B FE D6 CD 77 F5 03 C8 5D
 94 BD AA 32 7D A7 27 41 AA 14 53 3E 99 D5 16 AA
 52 BA 23 2C A6 13 DE 75 2B F1 7F E0 D4 3C 5D 1C
 6F 42 99 9C 1C 72 1E 67 4C B2 6E 0B 03 3E CB 9F
 2A AC A8 80 78 B9 B4 72 70 52 6C BC 4C 97 1D 52
 53 34 A5 97 FE 87 A4 79 DE 28 65 BA F5 67 A6 8C
 B3 17 E3 6A 2B 6D 66 7E C1 B3 81 16 E3 64 BA 82
 02 F3 92 50 48 97 E8 DC D3 4F 09 30 8B 48 DC 98
 88 31 A8 32 F0 38 F7 6E A0 71 90 46 62 3F 6F 22
 6B 4E E9 53 16 AA BD 7C 1A D1 74 BB 61 35 B5 71
 85 21 7E CE 42 29 E2 1A 1B 67 08 AC B5 EA 0D E9
 0F 25 96 4E DB E1 1C 1D 67 6E DE 4A BE 61 BF E3
 C8 4B BE 3B 62 F1 80 A8 24 70 F1 10 78 61 39 D1
 55 7C 93 AA 3F 97 43 70 65 7E FE 7C 0B 90 00 F8
 14 2E 53 7C 9B 41 87 18 0C 9C 65 5C 85 FC C6 C5
 6F 9E FC 45 C3 9C B0 9C 4B 6B C5 9C 0D 77 08 2C
 A9 1C D9 B7 BD 3B 71 AC 80 C2 46 04 EA 5E 5B 65
 E3 11 CA AB D0 CE 08 DB 2A 09 26 DB 9E 0A 6D 1A
 B3 ED 4E 66 CF ED A5 C3 18 50 82 EC 5F 8A BA 31
 6F 21 DC 89 12 4D 2C 4B FE 52 56 FD A4 10 6F 59
 9A 23 03 D9 94 8B 7B C0 C6 62 FD 5D 88 71 A7 E4
 C8 63 DF 42 74 F9 A7 F2 F9 45 AD F1 F9 2A FE 18
 9B 1D 02 48 E9 BE D5 99 2A C7 2B 3E 4C 72 3C D2
 EC 1D CB 36 C7 5E 94 61 72 46 C0 72 80 F6 2F B3
 7A 5B F0 EB B3 0F DF 7B F5 F2 F5 01 CB 22 05 48
 50 CB 8B DB 65 C3 FD 72 39 16 2F 56 3B E7 B2 DF
 AF 02 45 09 E5 AF AB FC 08 8B 14 7E 78 5A 4F D0
 D1 22 5E 3A 11 4F 25 50 4C 5F 0E 1E 94 9C B9 50
 CD CF B0 01 F0 67 CD 3B E5 3A 04 8D 60 89 6C 6F
 28 B7 43 9B B4 0A EC 38 E3 C2 8B 1A AE F0 74 03
 42 EA D4 A4 29 00 4B 12 7E 70 8D 86 38 25 85 F8
 FC 33 06 23 D5 70 63 91 3F 2D 10 EF BA 92 1C 42
 14 3E 31 20 2C C9 2E 79 C3 8B 97 28 4B 5F 30 D0
 FE 75 CB C6 16 8E 6A 36 EB 80 77 CB E1 1F F7 A8
 37 60 91 2D D8 90 60 4B DF 7F D0 B0 D1 7C 97 41
 5E 36 52 20 40 10 F7 AA 7D 4F F2 4A 5A EB 74 48
 F4 82 0E C3 BF A9 E8 72 AB 29 F0 22 01 4E 7A C6
 0B 73 E2 0B 2F D0 3E BC 28 9E C8 AC 5F B7 6D 2A
 8C F4 A5 FD D1 2E F1 84 47 B4 3C E8 03 F2 BF 47
 A8 D9 C3 3D BE 58 65 CC 1D FD DD CE 65 90 0A 84
 F0 D2 84 27 EC 01 8D EE AD 0C 42 63 C2 E3 E1 98
 1E E8 04 8B 5D 44 56 30 75 26 5E 95 34 F8 78 E9
 ED 32 F8 3F A2 2D 39 C1 C0 A5 73 89 68 FA 0E 24
 48 06 27 C0 F1 F2 7D E2 A7 7C 35 F1 7F D3 CA 7E
 99 0A E0 C2 41 DB 19 1D 0F 10 0B 7F 6E 1C 29 73
 8B FF 0F F2 07 41 42 DF 6A 53 D6 A1 8D 1B EB E5
 46 E3 DA D9 11 AF CF E4 BA 3A 7F AB 70 E5 E7 4A
 EB 8D 32 A2 6E 5F 9B C6 65 31 0E C0 BB AF 05 BB
 CC 00 B3 9F 2A 4D 56 67 66 0B 3C E5 E3 61 06 1E
 01 E6 7E 43 EA 55 EB 09 64 00 7B 40 1E 43 D2 D9
 DC BF 92 2D CC 70 23 24 6C 38 A5 EF F4 30 1D 92
 69 09 44 63 55 75 83 F0 88 F6 55 1F 61 61 4E 20
 9E 7E B6 E0 92 EA B0 DD C2 5B 24 96 60 8D 51 16
 29 EF E1 AB 55 50 24 4F 44 77 A9 B2 4C 6B 34 93
 F3 17 68 99 A6 1B F3 43 93 61 14 65 B9 D3 2B C5
 A7 60 60 3A EE 3A 97 F2 16 D2 16 DB 51 CF CB 3E
 58 E3 82 EF A3 AD 53 C0 3F 60 32 57 65 45 DB 8E
 8C 7C A1 B6 07 FF B4 D5 7A 9C 1C 7F 68 90 D6 E0
 78 66 8B 7F F7 5C 2A F8 D0 29 FB A7 68 DA 48 22
 D3 0E A2 45 EE D1 A6 1E D5 FB 9E FF 8D D4 2D CF
 C1 CF 36 C9 CF 57 DD 2A 0C 9F B5 7E F3 D8 BE F9
 35 BC A4 2F 3A 50 10 A1 20 CE 63 FE 3B 6C 6D B2
 00 D3 3B 9F 24 9B BE EE F8 91 45 30 0F A9 96 FC
 79 A1 4A 08 FF 16 02 84 3B 12 68 B4 9B 04 B8 73
 F2 FA E6 94 59 40 A1 C3 75 22 3A 79 C0 22 83 96
 CE A3 23 C7 8D 8F F1 4D EB 1A B4 2A FD 84 08 32
 B8 85 78 CF AD 16 4C F5 F9 D8 3B 32 A9 7F A5 FB
 B1 4B 33 C0 18 2E 1A 59 0F 5A E5 39 E7 B4 2C EC
 31 2D 49 25 22 8C 5B 5E 57 F2 65 68 2A CC 58 9A
 27 0F DF A9 84 3A C3 33 A2 3D A4 E8 B0 EF 08 82
 C7 30 78 C9 9B C0 F0 67 82 C9 C5 0A CF D5 B4 61
 BB 1C 3A F3 3C CB 87 EF 78 91 9E 44 18 B3 83 DD
 F8 63 38 75 A0 7D EF 02 02 2D 7B 87 FD DA 47 4D
 A6 1B 19 5B 31 92 A7 FA D6 15 FD 27 3B 7B 8F 8B
 E5 09 C5 38 AC 71 FF AC B4 B0 F3 E8 97 4A E2 FB
 6F E5 74 76 A3 47 3C 30 8E A2 78 58 21 33 33 D4
 F1 96 3E 74 CD 24 B3 B0 3D B3 28 6C B2 B4 45 D8
 E1 2B 3B D3 BD FC 23 37 67 74 6E 77 4F 55 EF A2
 1F 85 7B 15 46 75 8E 13 9A FC 74 30 CA 15 EF D3
 2F CC 4B 79 86 F0 3A B4 F6 CD 05 4E 92 81 16 7E
 CC 6C F9 AF C4 28 FB A6 92 A3 72 5F 10 CA B0 F9
 24 8C 44 9A 08 E4 BE 64 07 2E 9E 9E A6 DD CB 92
 D6 DB 47 1C C3 C3 9C 67 C2 A8 73 03 92 6A 38 5B
 93 04 68 F5 C5 34 01 3D EB 65 D1 B3 0C 1E 94 08
 EE BB 4F 9D D9 BB 7E 38 38 A1 76 BC 99 1D 8B 4C
 27 7E 30 26 81 5F 52 60 B7 D9 2E EE 4B F5 39 78
 08 8C F2 B1 45 2B 29 89 21 13 F4 3B 47 5B E7 32
 67 FB 11 D2 80 2B 8A 1F 5E C3 47 36 85 7D 88 85
 E2 FF F1 46 30 C3 7D 77 8C CA DB 6A E5 FF AD CC
 C2 51 27 DE 6E BA D4 77 34 EE 84 45 33 74 8B 63
 B6 81 DF 1C 07 F6 8D 41 EB F6 BE E5 76 4D 3E 69
 3E B3 E4 96 3D 66 A6 7F C3 A4 84 79 E7 1D EC 7A
 98 CA FD A5 4E 8A 2A 8E 61 E0 57 C4 2A F5 E5 11
 B9 7F 19 BD A1 E5 5A D7 02 E4 63 6F AF A9 01 AF
 1C A1 1A C6 C0 E3 78 87 08 E8 7F 9F A7 D4 E0 D6
 38 20 AD B2 37 DF B6 C6 A3 BF 1E 80 E5 43 77 46
 29 35 BF 39 2A 88 37 FD 91 9E 5C 9C EB 07 42 DB
 80 71 C3 BA 7F 76 CC C5 65 B9 1B AE EF 43 7C 8C
 5F F9 75 98 7B 94 12 96 E1 32 14 7B 21 F3 13 81
 7E 76 A3 E0 19 8D B9 B8 B3 94 85 5A DA 25 18 DE
 43 E5 A5 F2 CC 11 0C D3 81 93 69 04 69 A6 F7 2D
 0A F3 AD 8F E5 A0 98 73 B4 46 EE C4 35 9F 0D CB
 5C 47 87 2A 71 4C 14 76 61 1B BA 93 75 20 22 46
 77 40 9E 56 7C B1 7A 61 44 32 92 BB 39 F5 9B B3
 C0 C9 F7 F0 77 EB A5 B3 D1 90 38 47 27 2E 6A 0F
 A4 21 74 FA E6 E9 B8 80 A1 CD F4 C9 CB 7C F1 B6
 03 F7 21 E4 FF 05 82 26 9C 5B FA 1B 02 59 07 8D
 2E 4F 47 5D D3 BC 27 87 D5 00 9D 81 37 52 A4 FF
 F3 5A 35 E0 18 17 61 13 86 5F 0D 1E 52 FA BD BC
 7B 24 18 76 FC BE E4 CF 59 7D 26 AC FE F1 D3 0B
 54 78 78 8A 49 A6 47 5F BB C2 9F 1F EB 44 BA FC
 D9 2A 00 94 47 CA 58 BA 54 F6 8C 06 7C FC CD D5
 83 76 FC 9F 8D 33 7C 47 71 EE 5F 0B A7 6B 95 EB
 11 E3 F6 D5 17 AA 65 1F D3 08 B6 86 81 ED 7A BF
 D9 12 6C FD 8D 9F D9 D2 96 53 03 F9 AB E9 EE B4
 B5 B3 2D 30 06 D0 7C 72 08 88 F8 AB 44 FD E6 BC
 E9 2B DD B6 5B D6 9F 3E 54 7C CD A5 38 C0 8A 85
 E1 54 0F 0C BB 45 D4 1C AC 8F 65 8D 98 D3 EB 97
 94 EE A6 75 52 6C 69 BC 3B 4D 7E 5B E6 B4 2F 97
 6E 50 26 C3 A7 A4 30 A4 3D 5E 32 7D 2B 64 BD 0F
 1E 28 BB D7 5B 4C 4D 1D 1F 1F 96 89 E4 B8 2C 74
 6F 9C 80 B7 7F 2D 95 87 EC F3 3B 16 3C CE 91 23
 26 85 DA 0C 0A 1A 5C F0 AA 44 C1 34 92 8C BC 35
 8A F3 80 CD 46 9A 0F 89 71 A5 04 59 F8 BD 51 D8
 54 F1 A8 0E 0F 53 77 08 B1 DF CC A9 26 44 C0 34
 6E AA DB 34 E3 74 95 DC 53 79 41 9E 48 19 F1 CE
 E5 ED 94 59 9E 90 63 AF 96 72 4F E8 96 D1 28 29
 C3 B1 B9 D3 E6 31 48 C8 05 88 95 04 5A 5F 4C 6D
 67 69 C6 09 3B BB BD 19 10 CD C2 B2 12 3C A7 60
 05 14 E9 A4 81 DF 00 6C A0 F6 A3 04 EB BB 8F 10
 02 C4 08 8F 7B 62 2A 41 EB DA 2F 90 C5 FD EA B8
 58 CF E8 BC 35 9B 8E 71 39 57 42 BE BB 8B 09 59
 89 76 50 B8 CD AA 1C F3 43 47 3D 53 5B 69 2D D6
 42 F0 9B 34 9B 5F 6B 38 4D 95 BB 2A 7A 1F DE E5
 73 D0 E1 A8 0B A5 FE 66 38 33 D0 CE 85 7D F1 4E
 6D 7D 15 0B B5 24 92 77 78 B4 81 12 44 6D F1 F5
 21 BB 37 7A 29 22 6E 56 CF D4 6F B7 18 A4 E1 AC
 B4 FF 9B E3 3E D1 37 0E 38 39 D3 70 14 EE 6E C2
 87 E1 27 1E BB 13 35 74 60 7C 09 CA 74 4D 17 F3
 B2 00 0D 50 0F 96 7D 46 8F 38 72 DB 9C 38 CF E8
 64 00 F4 57 93 46 25 D5 73 48 05 AE 53 74 F9 98
 BC E2 F7 4F 0F 17 13 31 C1 91 E4 10 97 97 C9 D7
 54 00 6C D2 4A 04 E7 8D E2 99 59 6A 53 B1 5C 88
 F5 28 76 71 4A 9E 1A 5C A2 39 3A D4 2E 9B 90 DA
 B9 DD 1F 26 2B 77 05 97 9E 5C 70 44 C1 6A D4 89
 2A A0 14 92 B8 05 DC 41 66 40 0E 0A 47 56 1B 35
 AF F3 18 DD 4D 8A 02 F9 2D E2 40 6B D9 11 4C F4
 B3 28 98 08 83 EB AA 09 FF E7 8D EA D7 C6 C9 76
 BC 62 C6 58 57 3C 22 05 24 23 31 2C 61 34 D2 A1
 99 49 72 B5 95 A1 6C D8 FE 47 7C 68 B9 F6 26 2B
 9B C8 3A 90 D7 FB 13 19 C7 76 04 CA 42 43 9A 3B
 98 77 69 36 12 9E CA 86 D8 B6 2B D3 89 25 43 90
 6F 4F 41 2D 7A F2 D2 EC 88 41 FE FA 20 E7 4C 68
 31 FF 57 B2 1B 6E 4A E8 FC 5E 7D 4F 8C 49 F4 13
 9B 2C 98 4D 76 4C 74 E8 60 93 AF EE B0 19 14 A4
 75 8C 00 F3 2C 04 C8 D0 0F B1 F5 A9 13 A2 AB 8C
 26 3A 32 12 4D DA 59 66 41 E8 F8 02 5C 5D 34 C9
 BE 2C C9 76 B8 CA 47 67 19 4E 64 56 77 B2 38 35
 27 73 FD 88 F4 1A FA D4 D0 D6 7A 69 EF 5D 39 7A
 BB D3 2D 7B FF 07 44 74 8E FF 35 4A 6B 9B 4F 7D
 95 37 EB BF 84 7A F2 57 83 74 9E 7A 53 62 99 DA
 68 FA 9C AB E7 56 99 B6 D5 F5 15 9B 4D 5C 26 6B
 37 12 00 94 26 F5 97 AE 0A 89 16 92 50 86 8F 84
 3B B9 D9 4E C7 DC 96 18 FA A4 0C 57 24 CB E7 A3
 59 FB F4 F9 59 56 F6 B5 8E A1 6A 08 55 45 47 4F
 7B 00 1C 79 7F E5 40 81 F3 FA B5 43 E7 D5 41 1F
 09 46 AC 26 3B CD C7 B6 CC 79 99 16 2A 99 E1 10
 F6 3F EB 5C 51 D7 38 75 DF F9 CC 9E A9 A3 44 C3
 76 45 D7 26 BD 90 FC 1E B0 54 DB E5 F1 38 35 10
 7C 57 A3 A8 96 F5 6D F6 76 C4 81 DE F2 7D CF 7B
 7C 1B 7E 6B F1 18 49 8A 37 5F DA DD 56 1E 35 16
 81 21 12 14 15 65 46 20 84 CA 65 2A D9 76 E8 B3
 A5 29 8B 77 94 3E 8A 92 A9 BB D4 1B AB 68 65 6F
 72 90 91 3F B4 37 9B 43 37 1B E1 C3 BE 1B 75 D1
 1A 63 4F E5 2B 8D 90 AB 66 57 03 2E 06 EE 6A 26
 7F 46 15 C6 89 EB 74 A0 C9 5E 5B E3 E4 CA 48 35
 2B A0 D7 70 11 44 EB C1 3D 62 B4 DF BA 5C DB 91
 86 2F E1 5E 3B 5B D7 04 32 80 01 DC E0 25 C0 E9
 A1 57 04 83 33 8C 01 6E EB 04 56 F1 12 04 D8 18
 23 DC 53 F4 91 1C 5D 4F 19 F9 D1 29 D6 E2 CE EC
 4F 92 5F 0A D4 35 4A C5 A0 BA 4E 2F FE C8 DA 4B
 8B 75 FE 84 63 2F D6 5A E6 66 D6 6A 8E 95 62 2E
 49 F0 4D DB 61 38 DD 05 AA AF D9 AE 45 C7 A4 3D
 82 20 FE D4 43 E0 0D 97 81 4F 86 C5 6F B8 8F E4
 03 01 14 EA 5C 07 2B 9B F2 20 A2 09 D4 8F C2 9C
 9C 2A 0B 7D F7 7D C3 18 B6 98 D1 7A A7 1A C4 A7
 A9 7D AD 46 B1 E8 69 01 E9 ED CA C4 E0 A6 17 57
 50 AE CD A2 5B 52 18 B6 B9 6B 07 E0 05 49 9D EB
 0F 89 39 D6 F7 4D 27 5A 95 1E E0 4E 80 44 17 4F
 6D F1 BB CD B8 73 D3 01 88 1D 97 1F E2 C9 34 C4
 53 49 2E AE 7F 74 D7 E9 65 D2 50 7F 1B BC 4F 3B
 38 A3 C4 4D 1A EF E1 4A 5F 42 91 9C AF 22 C4 73
 61 4B CA F7 40 AA 2E 90 4E 36 23 6A 56 3C 93 58
 0C 8F 2A C1 AB C5 B6 69 7D B6 0D AE 9C 14 15 A8
 18 B1 46 14 AD EB C8 8B 5D D2 07 A7 66 26 78 17
 A2 C8 1D 94 F6 AB 89 A4 07 DF 0B F8 1C 2F FF EB
 76 19 A3 F5 12 64 2F ED 6D 2F 7F F3 D9 5B CA 84
 47 8C A8 D3 FC AD E5 FA 61 E7 95 E9 61 1E E7 6A
 9C 0D 54 69 B9 7C 9A 48 5E A1 77 CC D8 8F 86 37
 65 6A 0D 5B B6 CC D6 F1 02 11 91 0A 86 53 9A FC
 25 34 ED 3A 13 E7 D0 9A 1F F8 E5 59 3E 1A 99 0C
 83 26 D2 74 64 A5 C4 76 D6 21 1A 5D 31 50 BA 55
 52 73 49 14 15 A5 BF 84 CA 2C DF 02 08 11 1A 52
 92 38 B3 90 E7 34 47 8D E4 C9 99 14 D7 FA 39 1C
 57 08 E6 6A 24 F4 E0 3E 0C D3 69 3D 3D CB 63 0D
 51 3E DB 32 BC 82 E4 95 94 F0 25 A9 2B 4F 56 FE
 C0 21 82 92 F2 48 12 F4 8A A2 21 72 08 9B 6B 82
 79 1F 90 00 8B 1A B5 49 A8 DC 70 C6 C3 8E 56 12
 57 8F 8D 21 7A FD 85 9A 07 FA 5C 2F 36 72 60 24
 55 61 A4 17 2D 42 5C 99 D9 7F 35 A4 A5 9B BB B4
 57 ED BC 83 80 62 B4 36 9A 8F 9E 3E D2 ED D9 D7
 A5 BA 2C A9 8B 81 4F 49 AD 59 62 90 49 EF 48 D8
 31 B7 5D 5C 90 1D 2C DB 18 FF E4 FF DA FB F0 1E
 AA BB 06 45 C9 48 47 CC CD 64 00 FE ED 55 3B 43
 41 1D AB CB 04 9D F6 38 2C 24 6A E5 A5 A1 AA 43
 3F 62 C6 9C FF 40 F8 08 0B 2B 55 2B A2 BF 3F F2
 31 37 25 2F BF 1B 36 F2 79 08 00 F0 10 2C DF 5D
 3D 0B AC BD F4 BC 29 62 6D 74 78 0B 8E 74 98 8E
 01 FC 5E CD 5E 24 38 86 21 FE F2 41 3A 5A 8B 3C
 B6 7B DE 13 14 3A 5D 76 CC 30 D7 D8 99 D8 5C 25
 DF DE 51 8D AC A7 31 2F 05 26 DE 8A 49 0B B9 17
 A7 DF BB A9 48 D9 C4 96 0F B8 E1 A1 E0 8B 48 07
 3F 2E C6 4B 81 5B ED AB C6 95 65 27 74 CF 7B EB
 F3 6B 03 C3 28 DF 53 74 6B AD 54 FB EC B6 92 BD
 D5 1E CB 7B C3 50 F5 F8 28 C7 BD 65 5F DB CA 7E
 13 1B 47 11 F2 C6 ED 58 31 DC DC 42 28 1F 95 2D
 EA 1B 3C E9 CC 6E 8C D8 04 B3 55 65 D8 3D 73 8E
 85 E0 E4 4A 19 07 77 32 C8 A2 6A 06 F0 5E 2B 86
 6C 7D 9C 79 C7 C9 92 B7 DA BD 1E 98 DC B4 10 53
 2A 09 32 6F 45 3D C5 86 95 9E 9C F6 C0 1F BE 26
 78 D1 63 75 AC F2 08 B6 64 1B 86 28 E9 36 BA 5B
 40 BB A3 CE 06 91 47 0C 0F F9 E5 A5 8A 8C 9C B0
 9E D5 58 BB AC 8E 9C D9 57 44 21 60 E3 41 B9 71
 FC 1A B4 89 70 F7 54 52 45 3C FE 43 CD 79 D7 4B
 10 DD 53 7B 5C 4D 0A EA 16 37 8B 83 67 FC B6 37
 BC 6E E3 45 85 A2 B3 E1 CF 59 0E 85 7C B5 3C 6F
 DC 69 78 8A 01 4B B1 87 40 CF 39 70 DB 9D 8E 24
 C0 7D 7B D1 E9 01 A1 43 48 B1 91 96 66 F5 1C E6
 D7 AD E9 F4 79 BD 23 3F 4D FA FB 67 C8 A6 7B 64
 60 EE 69 78 A4 FC 08 D7 DC 39 92 0C 48 CC 2F D6
 1D 26 8A EF 27 30 80 1E 1E B2 D3 5E 4D E2 97 64
 6C 3C 3D C6 8A 59 A5 64 12 80 9E 67 FE 3F 37 E6
 B5 2F 2E FC 66 14 8B 8A BF EA 66 47 A0 D6 C2 8A
 47 E9 9D 3A A6 47 95 EA F7 53 55 B5 FD E0 AA 9A
 C7 C8 28 9E 93 36 A3 CF F5 01 B2 10 D8 AF 2A 7D
 56 A8 FD CD B2 78 A9 33 05 91 AF FB CE 5F 74 67
 0E FC BC D4 FC 1F B7 84 34 FA A3 E2 4D AB 05 84
 0E 3B 39 F4 30 F2 62 A5 55 93 5D BD 20 C6 7E C6
 08 1D 5B AB B7 93 64 89 D2 38 DB 26 D3 56 00 ED
 06 D8 FD 89 0B FC 18 FE A0 0A 81 81 64 3C 4E D5
 CA CA 41 5F F2 49 FF 59 85 C7 61 E0 68 15 0A 1A
 4B C4 09 B0 77 78 7A 6F 14 EC BF 4F D2 3A C5 59
 09 78 15 3C 80 63 0A 00 E9 5F 5B B4 6B 70 AB 9F
 F0 5C 82 DA DA 4E 19 75 12 AE 28 C7 7C 85 2B CA
 C0 5A 36 68 8A F6 70 EA BA BF A5 EC F5 B7 4E FB
 B5 19 B8 7E 54 78 30 1F 40 30 3E BB AE 15 11 99
 98 C2 0B 77 D6 3C F0 33 6B AA AE 72 FF 31 28 13
 E5 55 57 7D 59 5B E7 8F 3F E7 D6 BB FA CA 83 F7
 32 C0 11 08 42 A6 35 3E 15 A6 67 D8 08 BA 0D 0B
 BF 39 16 EE B5 50 0B E9 B1 B0 FF 39 F7 73 92 6F
 F3 D3 DE 4D BD 13 29 67 3E 7B 55 A9 11 44 EF E1
 F7 DF 24 FC 3D 3D 25 08 E5 D8 0D 21 EE 30 2B DC
 0D ED F1 FF 5E 28 55 70 BA 60 A1 4D 92 E2 04 EB
 67 E5 76 7A 17 02 0D 5B 30 47 BD FB 94 6B C4 37
 F1 81 DF FD D5 20 D8 00 E7 50 2E 32 93 38 02 AC
 A8 2A 62 23 C5 DC EC B4 DE 02 62 46 75 D4 9C E0
 BA 53 CA C3 C9 64 FF CD FA B7 00 10 8F B6 85 E5
 33 27 27 14 39 12 59 61 70 9B 57 44 71 E4 8E 4C
 1B EC F4 F5 33 DB A8 B1 31 A6 5D BC 84 C0 D5 40
 AC B0 E8 5E F8 61 68 84 01 5B C5 60 D5 3D 0C 06
 1E 33 88 9A 9B 87 66 87 ED 0C 44 C1 7B 63 98 05
 79 95 20 64 45 07 1E DB 29 D4 9B 74 B0 29 91 9A
 B8 87 D5 24 5F 34 DD 63 07 F2 CC 9F BC DF D4 C4
 01 84 F9 9F 62 36 F6 7C A3 BF D2 CB 96 A9 D0 F8
 0B ED E8 75 09 43 67 A8 F3 4C 42 D7 D5 35 81 F3
 FB F8 2D EE E2 D7 A9 81 F8 4F 6E 76 D7 C3 7D 2C
 E5 39 BF 11 3C F2 7F A3 61 25 94 17 20 90 41 D8
 82 34 7E E6 36 F5 B7 D1 56 FD B3 0F 8F D7 62 C1
 A9 C3 F5 D0 90 B5 6C B0 04 C4 B9 BD 36 B5 9B 79
 8B A5 EF 07 5F A0 19 63 82 EB 6E 32 E8 E9 C4 50
 0B 86 46 1D 91 CF 3A 64 BD 23 C4 01 54 B5 FD 04
 47 FD CA FD 4F 4A 90 E2 CD 58 14 60 EE 27 4E 4C
 A7 9B F2 2A 7D BB 1A 51 F9 E2 F8 EE 9F 39 AF D6
 AE 46 0E 61 5F 93 C4 3C 74 6E C6 10 B2 B1 CC 9D
 F5 93 63 74 BC 36 BA 9D D1 86 96 64 D6 15 A7 71
 46 88 61 7A 88 3E 76 2D EC 01 73 74 98 34 CA 36
 FB 3D 85 8B 73 94 C2 F4 A5 94 20 6E 74 CC F5 2B
 B4 BC B4 DB 0A C9 A9 70 B8 A7 CB CB 36 04 9C 73
 74 89 F7 CA FC 61 12 62 4D CD 1D 3F 45 E2 AE 3B
 DC 73 F5 27 DC BE FF 6E 33 33 0F 72 D4 0A 50 4C
 8F DA 29 48 F7 EC 17 10 EE 1A 91 30 44 76 8C F7
 48 FF D4 D4 A3 E7 10 61 11 A0 0C D0 4D 36 80 90
 21 3F 9E BF 53 6D 77 66 8E C2 6F 58 C0 99 DF E2
 D8 5B 31 8B 60 B6 BA BA 9D 69 AE E1 C2 04 75 DC
 50 14 42 74 A4 E4 3D 88 07 74 3F ED 55 07 FD 3B
 AF E9 BB 5B 50 42 41 15 E4 1E 3B BE 07 C2 6C 89
 5D 8C 54 FB F9 24 A9 AE 9B 2A 6C 20 59 6C 12 B4
 DA 33 C0 08 62 1D 7D 43 8E DA 1E 7B 33 42 96 AD
 4F A6 74 19 13 38 D7 41 45 1A A0 57 4F 48 42 D8
 A0 80 B0 2F 75 EC 9A FF 24 CC CE AA 5D 78 4D 71
 48 B8 84 16 75 8F 5D 4E 78 1A 4A 73 99 05 D1 AB
 6D 2F 94 C8 28 29 B5 44 33 6E B7 CE 21 04 2F 93
 ED 2B 5D DD 28 51 FA D6 3D 42 EC F1 AE 3F BB 25
 4B 17 53 20 91 4A 2D CF 5F 1C 62 3A 4B 7D D6 DE
 F0 13 16 0D 03 19 6C 30 CA 5A 27 D8 66 D2 91 59
 16 8B 6D 86 23 75 66 CF C5 E6 A5 69 11 36 A5 6C
 DC CD C1 F0 AB CC B3 E8 BE CA 9E 03 32 6B 94 0B
 07 D6 E7 73 32 CB 00 C7 46 BF 5D 0C E4 78 22 63
 14 7A 10 34 E2 3D 6F BA 26 B0 36 63 25 17 18 15
 1C 9A F7 8B 45 84 D0 06 96 17 B7 2A 8C 29 53 59
 2C 51 AF F6 DB EE 5C 74 6E 17 AF 74 94 DB 73 96
 27 18 32 24 BA 21 2B 15 F6 C2 6A 0A 2F D7 F5 16
 92 F3 3D 06 C6 A4 0C 9A 1D 3F 1E 8D E1 1F E5 14
 A8 DF D7 0D 4B 9C 9D 32 75 F5 52 87 4F 42 71 70
 05 56 E4 86 C4 34 07 ED A8 47 63 A6 74 E2 72 68
 45 4F F7 1D 08 FD 71 25 E2 DA 09 91 AD D2 C8 43
 8A E4 3A 10 2C A2 BA 24 AA 66 39 E6 32 09 E4 98
 EA A4 23 DD AF 32 DB 00 F3 B8 E9 7B 0A D6 23 C4
 51 BB 06 C6 46 7A 3F 59 46 65 A6 D5 12 24 32 70
 DF 85 CB CA 62 E7 CE EA 4C 6B DE 73 E9 A6 D2 B7
 AC DF 96 31 CA F3 34 F9 BE DF AD C0 FD 99 48 3E
 29 FF 6E E8 7A D2 25 A8 70 36 56 67 5D 55 D4 F2
 AD 6C C1 4E 2A 8C 83 E2 63 B5 35 4E 75 36 4E 31
 DB 2C BA 0E BC F2 C8 62 6C D9 71 7A 4F 0A 11 5F
 6C BA E6 B8 75 27 70 64 C4 E5 2D EE 1B D9 A0 40
 6D B3 0E 20 C4 B2 28 A2 23 E9 B2 49 2B C6 07 42
 63 99 7B 39 CA F2 3E FA 41 D9 E2 A6 22 B3 32 54
 47 78 78 A6 1A 3E DD 38 3A 19 48 DA F5 38 D0 D8
 30 FF 70 E7 D6 BA 3A 4F CA 74 57 C7 76 2A 75 22
 81 0F 63 E9 AA 1C 7E F7 98 D8 B8 A8 A6 4D CE 1C
 63 1D 65 46 2D 50 1A C7 2D C0 D8 A3 7C D9 E3 79
 C2 57 35 45 1F 66 A3 10 1A DD AD ED 9D B8 D5 23
 76 B7 96 12 3E 8C DA CA D3 BD 67 0D F7 BF D8 24
 8C DA 3B 2A 67 19 59 8E C9 0C 56 43 F1 C4 06 48
 B9 C7 33 04 EE 32 11 64 F5 89 73 64 A2 35 12 BB
 A5 AB 77 48 B7 B8 97 FB C9 75 E1 A2 31 02 85 B1
 11 CE E4 88 BE 1A 60 D9 BF 92 BC 6F 85 24 67 E6
 46 76 AA 6A 92 A9 AC D1 FB 75 17 6F 1C 38 33 9A
 E4 22 DE 77 A2 73 DE CF 4C 3A 47 A6 7A A4 D9 93
 FC 5D 28 54 36 90 F8 5D B7 8E 1F 9B 9D FB 60 E1
 F3 A0 E0 40 64 8F 27 F8 04 C8 8B EB 6D 30 38 4A
 AE F9 1F FD 82 7B E6 BC F3 D1 00 A4 68 DD A2 23
 4D 81 49 1F 9C 3F 9D 2C 9B 10 B1 34 C8 B8 5E E8
 FB 9B 09 6D 81 C2 F4 C2 25 85 79 AE 6F 90 48 BA
 21 C9 D4 26 C6 BC F1 11 42 8D 65 CB 8B C6 89 F0
 5B C2 B6 76 77 CE D6 44 55 13 F5 E3 88 5C 7D C5
 70 F4 61 88 5C DB 0E 15 07 52 03 FC 69 32 20 C7
 F5 21 10 AD 5A 11 DC F7 3A 29 1E C1 9A 05 BD E4
 82 10 7E 3E 16 5D 13 F5 A4 79 95 A8 23 27 E4 E5
 3D 35 19 F7 02 7C 36 1B AF C0 50 3B D1 A9 84 C9
 30 18 87 9D 47 21 92 F1 AC 98 97 2F 57 15 EE 5B
 C7 2F B4 C2 D9 B8 E9 28 EC E6 5C 11 A1 DB B5 FC
 0C A9 1C 81 B4 76 9B E3 53 63 A4 54 90 66 FE 3D
 46 20 37 88 80 D5 80 83 63 6B B1 38 E4 09 09 E8
 CC FA 06 C8 3A 69 24 1B 37 AE B1 40 75 2F D1 A8
 10 23 3D A1 3E 68 59 76 9C DF EF 53 29 DC BA 95
 59 6D 4B 6C D0 02 5B 05 12 84 3E 58 A1 A7 39 59
 1A 6D CA AC 40 48 97 6A 2A FF 02 15 C2 A4 07 5E
 87 CD F5 54 92 AB D4 2B DA 94 A7 59 45 BC 27 0A
 DA B3 69 09 51 B6 26 C7 B2 02 38 FC AD BB 62 73
 F2 1A 82 4B 71 B2 CF FB 2F 40 5D 91 C4 87 26 14
 48 A1 21 26 19 E6 00 12 6B 7A 7D B2 E8 3F 7B 01
 D1 A8 6F 66 5A 16 35 52 6B C7 6D BB 20 FC 70 94
 54 C9 AB BC 37 F0 A5 82 F0 74 01 2A 60 4B 9C E0
 0F 79 ED 1C C8 8E 38 B2 10 15 03 22 A2 40 62 FD
 3D C0 B4 2C 6B 99 C0 98 1E E3 00 05 00 89 A3 48
 AB 7C 03 2E 27 80 C9 E1 A8 8C 38 85 FC 33 15 BF
 AD 22 99 EE E9 39 AD EF 6F C0 6A 2A 73 66 95 AA
 8C 7C 14 6B 85 E3 87 49 87 81 28 69 24 57 70 20
 9A A0 88 EC C1 CF C0 8A D1 00 04 89 DB B4 06 F2
 56 CE 40 BA 66 88 7E 76 A6 A5 56 97 D8 59 CD 1B
 AE 74 93 9C 69 87 7B 6F A2 A6 AF BC EE 4E 38 A5
 E5 31 9E 03 0E F2 2D 9E 2F 49 67 F6 BD 03 C0 68
 17 AD 13 FA B7 1B 33 58 CA 06 07 4F 89 1E 90 D1
 3B 0B C4 6A 09 38 ED 85 52 1A EB B9 CB 28 84 32
 AB 13 0E B7 45 BF 9C 3A FF 55 8B 72 23 9C E6 7A
 9B 40 7D E1 50 7F 30 3F 2B 8E 68 DA 77 68 FD 16
 67 AA 52 6C D0 44 10 31 B2 23 01 87 62 28 68 36
 0F FA 87 7C 9B 85 86 33 2B D5 97 62 40 49 3C B3
 45 34 40 D9 EE 1D 74 86 14 F9 AE 71 09 A9 95 5D
 40 19 69 91 0F C4 D8 1F 22 9F 85 D0 B7 35 89 CE
 45 7E 98 D5 21 0C 72 DE 99 9F 01 E8 45 E2 41 C6
 4B 5C 4C EC B7 ED A5 CF 50 38 12 30 85 20 AC 4C
 21 71 7F D5 2E E7 A4 0C E6 2C 6D 50 27 98 91 0C
 DB 58 D9 75 5D 95 39 D5 59 52 7B C3 33 15 FA 1D
 47 8E 84 91 16 8E CD 48 1F 92 A3 58 6D 0C FC D7
 95 DE BD FB 65 8F DB 64 3D E8 AE F5 DE DA 11 75
 6C 78 D7 90 D1 43 B6 37 0E C5 28 69 9A 37 24 DC
 DB 1A 25 E6 F5 0B B6 71 A6 B9 EE 35 A1 F3 32 AC
 65 B6 38 BD BA C1 8C ED D6 D8 B6 7A 11 44 18 48
 9C A2 E5 F8 B6 7D 99 55 7A 87 46 37 19 AA 49 50
 98 02 3D BA D3 13 C7 AA F9 E5 5C E0 77 0B 7B E9
 A8 C7 CA F5 0B 82 5C 35 AB CC F7 AF F9 D6 1C 57
 3E FB 8D E3 26 68 85 1C F1 0D 8D 91 52 C2 24 61
 AD BA 57 6C A9 19 EE B3 53 FD 7B 3F 35 3D 7B 8A
 61 E0 93 52 E0 9A 2A 36 52 F4 24 40 77 26 FC 92
 BF B6 08 57 C1 F7 C0 07 2D 4B 5D F2 AB B8 05 12
 8C 34 AD 6C 96 4F 51 6F C4 C5 C4 24 64 88 05 3C
 27 8B 82 FD F1 80 58 7B C8 0E 32 BA 9A 66 C0 81
 68 67 69 6C 29 4A 74 5F A2 CD 70 DD 6D 9C 3D 25
 D4 BB E5 5D 51 55 E1 AB 7F FF AE A0 1B EC 10 F9
 C6 4C 45 20 59 C0 08 ED 77 A7 C2 45 40 99 AB DB
 CC 45 8C 2A DC E0 D6 71 13 00 05 90 AB 3F D7 2F
 E5 BE 26 9F A4 04 D2 E7 2C 18 5B 76 3B 9E 71 A4
 D7 E4 6E 31 CE E9 85 66 44 78 03 AA BC D6 7F 8A
 2D 4D 2D 1D 7B 68 5A 54 DD 03 66 62 CD E4 96 87
 C8 A8 39 05 2A 47 42 84 D5 58 7A 5A FA 8C EC F1
 22 FC 8A D8 6E 38 BB 04 98 9E 84 AE 27 E4 8E 5A
 07 65 83 55 BD 5D 01 3B 4E C3 3E 58 25 A8 54 22
 2F 38 FB 0B 23 40 1C B3 6B 1A C5 B9 35 93 9D A2
 89 D0 20 9A 16 6B B0 01 B7 4C B4 1B A6 7D AC BE
 40 C1 91 C6 7C 31 B9 54 62 C5 E1 B9 13 6E 0B 89
 A9 FA 81 58 92 32 98 EB 41 01 9E 4A 83 61 BE 92
 B5 65 30 1E 8B 6C EF C2 89 5C 2E E1 71 C3 37 1E
 34 A8 24 6C 41 B8 36 67 F8 B2 16 D7 FB 97 1A 4D
 AE 0B 69 2F 67 D6 23 7C 0C E9 17 12 78 98 21 49
 FF 39 9D 75 AA FB A8 56 B4 35 07 AD 23 EE 0A A1
 A7 25 81 AD 7A 8C CB 1C 1B 79 E8 75 72 B8 84 10
 14 86 88 13 70 F1 A2 01 F7 E4 DF 23 5B 24 70 CE
 97 8C C7 64 CB B2 3A AB 8C FE F0 11 1F B5 C5 BD
 C5 0C 1D 99 4D C5 B5 CE 65 EF 9B A1 8E 8E AA B9
 18 56 90 84 23 D0 32 37 36 14 D7 68 BA C0 4C 9F
 90 61 A4 17 A4 F7 C0 C6 8A 62 FB F9 05 6F 7A 84
 0F 34 69 2C 09 82 4D 84 6D 1E 3E A8 66 FA 6D F2
 BF 9D CF 7A 32 9A ED 01 7D CB 1E 11 0B 8D 8D 52
 97 7A C5 A9 F8 E2 56 F0 8F AA EE C0 91 A4 3C 5A
 B3 37 20 F6 EF 80 22 CC 7A 85 75 75 03 19 B3 B1
 3D 3F C9 25 91 26 D6 3F CE 05 F7 EF 35 7A E7 F8
 E2 23 99 E8 9A AD 24 18 12 C2 1B 59 1C 58 53 ED
 7C BE FB A5 4B 7E CB CB 40 CF 6A AA AD 91 8A C8
 F3 6F 93 49 10 3A F9 F4 F4 43 F0 7E F9 C7 B7 BA
 F2 28 60 21 1C 73 54 E5 61 A1 81 21 D4 9A AA 97
 52 75 19 E2 02 F7 1B C8 5B 03 33 B8 01 3B 8B B2
 10 3F 68 0D 75 A1 36 E7 06 C0 CB DF 4B 26 73 B9
 2A 94 63 99 44 81 1A C4 DB 8F 8E CD 91 E8 21 E4
 44 EA 9A 49 62 14 48 6D 8C 5E 20 59 B3 D5 49 F1
 0B 78 5A A4 50 C9 5E AA 7B 60 A2 42 3F 51 6E A0
 90 7F B8 07 27 9A D3 03 96 29 B1 C4 E5 67 00 C7
 24 08 6A 27 C4 61 C6 5F C5 91 1A A1 B9 00 2B 35
 9B 55 9A F9 84 C9 E8 2A E3 31 32 04 61 2C 73 39
 0E D6 51 DC 75 E0 A9 C7 81 19 9C 0E D4 73 13 98
 AB 4C 36 8C FA BE 31 53 07 30 A9 59 5F 37 37 4A
 FA 3D 75 59 72 CB C2 FB 26 84 5A 07 6A D1 7D D1
 54 5C 87 1D FC 48 0D B0 C4 DF 06 3A 5B 6E A7 37
 E8 96 B3 39 B9 03 A3 99 40 24 CC A3 AD 89 87 B1
 64 40 07 9C 19 EA 09 57 E0 64 44 50 FD 4C 26 C5
 28 C9 1B 4C E4 CF 51 E3 62 36 AF 6A C5 E7 26 3D
 94 2B 23 F2 C1 DB 75 25 3D 9F 22 49 7A 49 A3 C7
 4B 6A D9 AC 56 73 4E 43 94 C0 03 6D E0 B3 AF F2
 22 7B 7B A1 AB 4E 2F 0B 28 CB 98 6A CE F4 C9 84
 33 DA 94 33 30 6D 70 BE E0 96 0F 91 75 45 CE 2A
 7D F4 A4 24 41 61 B4 2C 47 67 1F 86 5B BB C3 2E
 53 BA C1 B8 6F 10 0A 9B E1 14 DC D1 3C CD C2 E8
 C9 07 73 BA 07 CA E6 15 15 F6 ED 39 EF BF 69 C2
 10 C5 F3 D5 82 24 11 20 DF 2A 61 1E 63 02 33 FE
 B1 D2 92 5A 81 80 2C C2 47 54 FD A5 07 B7 B5 88
 67 34 32 9B 43 85 24 32 8B FB 72 16 E1 AE 15 F0
 5B E4 FD 71 3D CE 67 E8 BB 97 BC 6A 06 1B 9C 7A
 8B 60 E6 D4 22 B5 F3 95 EF B2 A5 E1 84 CD 03 E9
 76 EF A4 0C 7E D8 5F 9F 3D 0C 76 88 EE 0C 4A 38
 2E AA 77 E8 BD 7B 70 A7 72 62 15 D4 25 81 7C 5E
 2B F1 FD 24 5C 1F E1 CA 31 9F 2A D8 37 E9 F8 D6
 80 14 1D FA 6D FE EA ED 87 B6 16 87 4A F4 50 49
 E6 A3 62 90 E4 5E B3 48 79 94 23 7C 50 64 7F 27
 BC A1 83 A1 84 22 23 50 60 31 9F 50 10 4D FC 76
 4D A2 0B 2D F4 37 89 66 16 A4 86 12 B6 F7 19 A6
 70 D4 ED 7F D2 E0 62 3E 99 B8 8F 76 39 46 90 2B
 6E 2F B0 A2 5B F1 64 1F 14 AC 4F 3F 3E 68 74 F9
 A3 DB 59 70 8E DD 2C A4 DA 0A AF 36 E2 9C B9 A8
 A8 58 24 5D 14 0F 1D 93 9C E8 FA BD 31 CA 47 9D
 68 F1 81 42 0F FE 2F C3 F5 C5 12 5F 26 0A CF 8B
 83 7E 36 08 0D F5 59 2C 7C 3E AF CD 31 67 8C 4D
 07 02 F1 85 F8 B8 2B 3D 65 C7 AF 2F 5B 23 DA C7
 BD 89 9E 2B 09 EB 12 83 36 56 F2 AF AB F5 FE D6
 09 05 88 F1 9D 67 0D AF 08 54 23 51 B2 22 A4 6C
 58 D7 23 F8 0B 7C D5 8D FC E9 9D A4 F5 1E 22 62
 11 A0 E6 9E 24 87 50 13 EA 4B BB 15 C3 01 B4 0A
 E6 6D D8 2C D0 43 EC 15 83 BD 37 1B FF 5D C1 26
 87 16 28 34 22 D5 10 76 A1 A8 79 FD CB 60 0C 24
 BC E2 D7 93 73 EB F5 E5 DE DE 2C 18 A7 72 D3 E3
 C3 51 F7 8C B2 25 3E 83 94 66 39 3E 0C 5F C5 FB
 43 3F 31 9F 37 50 16 10 92 3B 81 99 20 58 E9 AB
 55 78 C2 F5 E0 A6 FA AB 26 EF 7E C3 23 2B 56 90
 69 2E F8 2E 2D 67 3E D0 17 3D A5 54 E8 1D 7E B6
 33 F4 2B 25 B5 D6 65 59 71 C2 E6 BF BB 48 C5 02
 01 1D 3C AD 1C 63 DF 90 7D 28 8D B5 7A CC 52 71
 3D B6 53 2D 34 22 81 A7 50 54 ED 18 3C B9 1E B7
 98 CA A7 3E 0D 87 9A 31 A6 26 5A 84 2F 22 86 66
 AC 4B 22 33 6B 15 2D 48 8F 55 F6 12 06 73 76 0F
 BB D9 D9 D1 AA 10 5C 55 36 D2 1D F8 EF FA 68 4E
 F8 18 7E A2 FA C8 77 77 19 DF 8A 58 66 16 60 67
 A0 E6 8E F5 A2 63 6C 7D 0E 6F 55 93 24 7D C4 20
 C4 97 81 F3 6E A6 5B D9 2A 7F 21 FC AD 4A 51 E7
 A7 66 F7 05 E7 F2 4C E6 29 0C 59 1C 1E A5 20 EB
 01 02 96 AB 87 79 57 36 D7 2D 21 55 F4 C8 7A CF
 F5 10 32 7D EC 65 00 DC 5F D2 46 98 2F F1 F5 79
 92 C1 5F 91 14 7B 23 25 29 6C 96 92 B7 58 78 6D
 F0 C3 F4 89 BA 27 EE 75 4A 5D DA 94 38 FD 04 59
 26 06 1E B4 1D 4F 23 22 D2 F3 3A 75 77 D7 41 3A
 82 9E AC 3B 17 9B 91 C2 BC A8 85 7C 12 80 42 68
 EA F8 63 E6 CC 6D C8 09 D8 8F 2C 98 D4 66 60 31
 E1 FB 7C EA 86 0F 4D DC 46 C8 38 00 8D 4F BD 37
 03 A5 D7 24 67 E5 BB 92 46 E2 30 DA 67 EA 83 73
 6A 33 AB 77 47 B6 66 C5 FD A5 CB A0 55 E3 93 31
 3A 4F 4C 6E 35 7B 85 AD 73 01 76 8E 74 D4 14 26
 91 B0 C6 72 7F 2B 44 7C 0B 65 F2 EE F5 83 F1 17
 FC 19 95 5C 5B 01 2D 6C EF 44 C2 C2 15 5C 8E 49
 B4 7C F8 92 50 90 5E 7D CD 25 81 1F 4D 73 71 D5
 15 08 27 26 2A 27 BD 3F 2E 12 3E A0 C3 E9 63 8E
 99 F6 D4 49 E5 C7 C6 FA A1 EB 3C 62 F1 FF 21 DB
 29 38 1E 16 67 32 61 04 BD 11 C1 59 77 95 F9 FB
 61 D2 B2 CC C5 B1 63 4B 01 BB 18 1D 1B 02 90 44
 A0 E0 B6 01 7D 14 EC B9 E8 8C FC 6F CC C6 E3 16
 76 E7 3A 1D 01 AC 1B A3 3A 55 41 2B FC 8C 3D FA
 56 D6 8B 1E 9A 06 F5 EA DE 14 05 32 B3 21 EE C9
 92 61 7C 76 67 98 6D 6E 04 99 8B F7 61 43 5C F0
 8A 18 DA 40 B1 77 08 B8 35 12 82 9E DB 6A 83 5B
 A9 2E 2A 6B CD B4 08 F7 B6 9E B5 0C DB 0C 7B E2
 F9 5A 1F F9 C5 FB 1C 3C 9D F2 C1 EE EC B5 67 91
 08 13 EA B2 91 8F A2 D3 D6 B9 76 CE 67 03 6E 8F
 0B 65 B2 17 85 0B 42 3A 10 BA 56 44 A1 3A A9 6A
 99 54 86 C8 29 97 97 AD CA 5F 7C 13 F2 A1 17 86
 E0 D7 65 83 84 28 22 E3 A6 E5 40 D7 36 2A 93 F2
 D7 52 CD 33 38 FC C5 A1 B0 81 5F A4 E8 0F 0E 55
 0B A8 45 40 3B C0 B9 A3 F4 7D F2 DA 9D 23 31 C4
 73 AE 1B 16 3A E8 13 82 10 0A 02 7D 28 A9 44 7E
 8B 65 46 47 6D E0 96 CD 4E 7F 76 49 BB F4 3F 8A
 5F 52 FA 67 85 A9 78 13 55 CB A4 F1 70 06 06 97
 F4 84 A6 00 CA 8F 30 1E C1 DA AC 18 2E 53 1F 73
 F4 1B DA 39 4E 83 A3 3C 28 0D 44 A0 AF E4 04 28
 F8 82 EA 3C 7B 4A D2 3E 83 87 01 05 EA 56 3B FF
 39 56 B9 26 53 DD 03 AE 08 37 E1 EA E1 68 1B 21
 86 C8 05 A0 E7 EF 0F 15 67 A9 D3 AE D5 9A 54 1D
 0C F5 41 96 5B F0 B4 A0 8C 4B D0 B7 12 EF 9C CE
 40 83 2F 3A A9 08 B4 F9 D3 F2 41 2B 2D 17 EF C4
 FA 01 D2 B3 CB 48 AA CC 73 54 DB E1 BE 53 59 2C
 8C 29 71 BA 4C 9B 31 CC 25 FA 6B 21 F1 AD 3E 58
 8C 5D AC 83 A8 B7 00 C3 5E D9 AD 44 20 12 07 52
 68 6F BF E8 DA 11 81 90 45 56 F3 29 8D 34 80 BA
 5F 3D 86 A4 54 61 83 D2 7E 2C 97 23 2B 3F 62 1F
 BA BD 00 32 85 B8 69 C3 F1 AE E9 E9 D7 0B 8E F1
 CF 3B 61 3B B3 7D 17 DB CD 20 25 F0 3D EE EA 13
 B3 6C F6 21 97 A6 9A 4A 87 34 62 87 EC D1 62 35
 12 D9 44 A8 B0 F7 FB 39 62 00 51 01 E3 B1 10 8A
 8E 19 1A 2B D5 05 6D 68 B4 4C 9E E5 F5 BB 40 EA
 89 08 74 23 04 83 43 9E 57 4C 5D 33 8D 29 75 08
 81 0C 84 28 7B 5A D3 93 EC F2 CD B3 2C 7B 8A A6
 4D 1C BD 96 CB 70 FB A6 25 A1 DF F5 DD 12 D9 7C
 90 36 E3 E9 AA B7 1E B6 EB D4 3D 0F E2 A2 5F A8
 C2 70 8D 0D 1D AA 7C ED 78 D8 6D 6D FE 0C 36 F8
 3C 29 DF D5 56 B3 84 FA 5E 3F 89 48 EB 3F 85 2B
 59 C8 5E 93 47 BD 34 C6 48 5D 33 46 A5 B3 4C A3
 4A 35 D8 9A BE 0E EE 73 03 93 82 B4 86 9B 4F C8
 61 12 91 18 63 65 B8 A3 FA D2 C4 76 31 FC 8E B5
 E7 33 24 52 BB 9E 6F C9 8B 97 3D 8A 50 32 99 25
 6E 4D 98 CA 2B 09 43 60 0A CF 4E 48 2B E0 F0 0A
 CC 1A 0A 9C 17 9E 5C 48 2C FE 8E D3 09 BB FF 50
 E1 67 2B 2C 5E CB 62 BD 95 88 9C 8F B5 C8 8A B1
 7D 58 6C 84 39 F0 73 FC A9 F8 31 75 28 E0 64 32
 3D 43 F4 2C 07 94 2F B4 8F 40 5C D9 17 5E 3A CF
 C0 90 96 C5 88 90 F6 EF 22 8F 56 B8 FD 86 0E A4
 38 60 42 6D 96 7E A6 B4 95 8A 7A 41 CA 0E AC 6A
 58 01 A4 96 41 DA 19 11 83 30 57 38 CB B5 55 F2
 82 2A B5 7A A5 97 68 A7 EE E0 8C 62 01 F4 7A A0
 53 B3 88 39 47 04 72 C5 36 E4 C8 27 97 6E 76 F5
 5B FC 34 6C CB 39 49 C5 6F D1 5D 3F 9C 38 DC DF
 8C 94 BB 3F 8A 1E 04 79 61 EA 7E 2A C6 69 95 70
 31 58 80 32 EE 08 95 40 FD 17 09 2A 30 7D 8F 31
 14 38 7C 11 D3 8F F7 0E 89 5F 7A 35 A9 11 E1 34
 52 66 48 72 EA F1 4E 06 83 CC A2 6A E3 AD 88 CC
 1B 67 02 08 5D 7C 23 A2 7F 20 FB 38 2F 35 A5 0F
 6D 3E 21 8B 3F F8 E5 38 94 76 C9 9C DE 06 17 12
 5A 40 D2 B4 A4 2F DD 84 C2 5B 68 8E 80 E2 6C 7A
 5D CC 61 02 31 10 67 5E A0 AA 18 5C 25 48 D8 C3
 54 B6 70 FB 03 47 70 F1 28 E6 CF 89 4A 86 C0 ED
 53 B6 53 01 55 51 80 CA 66 9B 4B DD 4D DA 25 D5
 8B 5E 58 FC 3E 29 82 C8 7A 7B 42 6C 75 16 19 2E
 CA E3 06 1E BD 90 C0 AE 84 B2 F2 A3 4A 1E AC 4E
 B7 51 18 92 55 73 9B 42 CE FA 6B 41 76 69 0B 0A
 29 15 F4 F0 55 95 16 09 52 2C 52 B2 B0 75 6B 77
 7C 0D F2 52 01 47 2E 2D 36 B5 A5 21 A9 91 EE F2
 DB 25 4F 59 B2 63 A0 E6 AC 30 67 1E C0 7B 39 B4
 C1 AF 3D 14 26 CA 3B 00 08 25 BB 91 61 51 4E 6E
 AB 08 72 85 C5 AE 8B 05 30 33 71 60 0B 88 55 4A
 88 D2 A6 B3 06 D6 AD 9F 3C A9 1F 6F B7 3F B8 DE
 1B 5E 02 DE E3 60 40 BB A1 B0 7B E5 FD 74 C2 C1
 9C 65 EE B3 7C EC E6 A0 DD 79 3E D3 86 02 25 35
 06 32 E8 28 F4 0E E8 48 56 0A 74 17 AE E7 6A 23
 DC 9B B8 E8 4A DD 7D E5 63 20 31 E5 73 E0 31 7A
 1D B0 E8 BC CC EE 90 FA 06 1C D1 1A 11 D1 4F 22
 12 39 A2 A5 E1 C4 21 2C B5 B7 AF 61 EA FF 46 52
 66 F2 06 8B 50 03 DC 2C C2 5D E9 77 6D BC FB 58
 7A 5A 52 35 FC CE 0A AA 18 48 58 2A 90 5F 6C D8
 78 03 B9 54 07 41 01 91 5F 7A DE B1 98 A9 FA 53
 A7 33 9A AE 58 8F B9 31 96 2C CD 4E 6F 92 61 1D
 5A BF 03 42 BC 11 61 0D 1C 67 94 B5 FF AD 56 94
 98 32 AC 1F 2B D1 7A 42 36 56 A5 DC 74 E3 4A A8
 F5 D7 5B 22 A7 02 F0 79 BE F2 A3 0B F1 93 0D 39
 F5 E2 35 F9 91 9A 0D 40 71 E0 AC CE B8 85 D0 FA
 CC BD 4D B3 C3 F0 DB 1A A3 AA 6D 5E 22 C5 EC 46
 C8 22 4F 99 C8 81 CC CA 92 A4 29 61 D4 40 3B A9
 2F B0 A0 DD E8 04 42 51 C1 98 92 64 2A 1E 1A 07
 23 49 62 7C 8E 6A 04 27 E6 1D C7 36 1F 98 17 84
 51 5F F3 AF A3 CC D0 E3 38 EC 19 CC CD 58 7A 65
 B1 2D 1F 99 0D C5 A7 22 77 C4 4C 91 C4 09 5B 1A
 69 51 8D 5A EB F0 82 8C 48 75 7A 06 84 7A E6 41
 5D 59 24 A8 FC 8F 08 92 26 D4 0C 56 A6 45 01 A9
 FC 08 40 41 6D 39 6E E0 CE 43 AE 14 91 7B F7 3D
 D3 05 F4 CB 32 FD DB A2 83 B5 AF 5A 7D DF B2 87
 59 7F AB D1 93 D4 95 36 DF 74 DA 8A 4E 96 B6 21
 23 9F 62 8F FB F5 79 C0 E4 CC EE EE 8B E1 A4 4E
 40 DF 66 42 64 53 C6 B6 CC 97 72 03 0E 17 C3 D3
 C5 B0 D7 32 E6 07 A5 03 A6 0D D0 85 D7 E4 3D AF
 4D 86 F0 19 6C C1 43 78 34 EB 24 87 30 23 C0 92
 F8 5B D0 3A B0 18 D4 E9 A4 97 55 3F BD B9 29 29
 FE 9B A0 45 A2 55 AF F6 31 6B A6 74 7E 25 1E 17
 72 3F CA E3 74 E7 7B B5 1A 62 90 0C 1A A9 01 33
 CA 01 20 64 E4 B4 BA 3E A9 20 63 38 2F 7D 75 58
 8C 3A CD 7A 23 A2 71 E8 E6 F0 B4 7A E6 27 F7 AF
 79 F8 B8 4E D7 C5 B1 AE 7C 34 28 AA EA F2 F0 2C
 17 09 F9 6E A9 63 12 29 72 0D 26 27 CC E0 9C AC
 FA C7 B9 2C 73 46 89 39 55 36 17 3A D5 FA 01 63
 F4 51 E3 07 7F 2A 4A AA 7C C3 26 62 8A 65 BB 4D
 32 16 79 32 CC 01 DD 8D A8 52 B2 84 45 47 2F A1
 B1 2D FE 60 C1 5D 9C 7F 3C 70 10 18 29 E8 C0 09
 58 6E 7C 18 59 7E E3 E1 F3 E3 A6 6D EA F9 CA 44
 3C 5B FE 6C A1 5A A2 60 11 68 F0 6B 08 F8 84 52
 2C 06 3C BE E7 09 CC A2 77 43 3D 5A 69 A4 99 B7
 C8 E3 09 E1 2A D6 FD 39 DA 4F 0F 61 F9 14 E7 DD
 5D 02 2F 10 83 78 B4 96 9A FE 91 A8 93 AD A4 D0
 A3 9D C8 9D 36 61 D9 8D 98 F6 CE E5 16 62 B4 67
 CD AA 2E C3 22 E2 DD EC F6 FD 2D 96 1E 7A BF DA
 96 59 DE 39 98 75 D8 24 38 C2 03 A5 98 C9 E5 B7
 25 95 91 01 60 37 C2 91 AC 75 48 98 F9 AD CF A4
 B9 58 0D 6A 6F D2 B0 7A CA AE 9A 47 03 AB 90 6F
 C2 F1 36 5D A5 05 3D 2A F2 27 45 24 0A DF 5F ED
 32 57 1D A7 59 D6 7D 41 2B 03 4C E3 0B 15 42 37
 36 77 41 A3 21 C2 6B C3 B2 A5 DA 8F 9C FB 85 E8
 C1 DD 78 65 4C 27 DF D2 BD 26 0A C7 98 27 7B 2C
 2F 8A 63 2C 6E AD 81 5E F3 CD 35 73 8F 97 B1 3A
 E4 09 39 9A 03 10 3A 39 75 5B 06 53 4A B3 1B 0D
 D0 FD B0 D3 41 E3 F2 63 37 F4 F0 00 01 6A 63 0A
 47 00 13 38 C5 4C 9A 29 B7 B5 65 A8 43 19 5C 29
 20 DD E0 EA A1 82 88 EF 8D B7 C2 4A A3 14 A3 77
 10 DC D8 98 F2 F9 E6 60 D4 E3 05 4B A4 94 DC 7B
 9C 37 17 F2 D4 D3 84 53 B1 9E EF 39 B9 5B 8C D5
 0C 1A 87 C5 44 33 48 C2 53 C8 05 01 E5 39 41 D0
 A3 62 74 5D 06 BF 22 C2 CA F3 6D 99 A6 CA A7 31
 66 83 54 C1 A0 C0 09 AD C0 02 E9 21 22 18 07 0A
 FC E4 57 77 7F CE B8 8A 67 A5 C0 10 2E E9 7A 3F
 1E 71 EA 98 AB 9B 38 95 C3 75 39 A1 A7 43 8E 0C
 4D 73 B6 14 93 9F 72 4D 6E F5 F7 14 36 98 19 8C
 43 65 98 2B 08 38 42 40 CB 7C 44 8B ED 7D F0 BD
 40 B7 25 4A A7 E2 9F 7C FF 8A 07 5C CA 73 16 E4
 C2 00 43 2F 20 3F 4F 4F B4 4F 91 C3 C2 2B A2 7D
 BA 54 AD D8 AA 3F 08 A4 FF 07 8A 29 F5 C2 2E B6
 13 76 1D C1 76 97 F8 8A 96 30 29 9D EE 00 9F 85
 2F 80 36 F3 C9 18 46 88 23 BB CA 99 05 73 57 77
 CF 2F D5 0E 0B FE 35 08 39 28 37 A0 CE 25 38 19
 91 C0 C6 4B 0D 12 5F 9D C7 A3 BD E7 49 6F 3A 79
 2C 68 95 2A 66 A8 42 6A CD 57 5B AD 53 C2 EF 00
 7F 5A A6 A8 2B 35 9C BA 5F 56 A2 6C E6 34 F5 BD
 27 7D 16 F8 88 F2 FA DC 52 0C F2 2A 62 6E 62 36
 95 9E 13 33 BC AC 52 BE 54 05 21 1D 5E E1 41 7F
 59 F0 17 58 99 9C 1A 29 FB 58 A5 95 A5 86 7A 59
 AD 1B EE CD FC F8 D4 D7 DD 53 93 A2 21 6B 59 22
 45 FD A0 C5 2B 4D 96 38 BC EC A8 2A 6B AF C2 A6
 B7 8C B0 62 A3 89 70 75 07 F4 D6 D6 42 D5 71 68
 D6 5C 1C 9D 14 94 54 E0 FD 80 E0 CB C9 A6 2F 9F
 47 C6 1E 54 FD 84 D6 2E 94 F6 DA 1F DE 6F 7E 2B
 80 29 83 65 13 67 47 13 80 5A 2C 8D 81 A3 83 CF
 67 73 7F EB 20 46 6A 3A 2D F8 ED 8D 63 49 6C 9E
 D8 B9 57 22 48 3B 62 F2 B0 0D 38 F8 D0 24 E1 05
 CE 6A B2 66 14 50 9F DD D0 3B 2F 8C 02 C8 54 1B
 F8 86 9D EF 14 6B 3A 42 C0 C7 AD 79 04 8F 49 E3
 FE 84 86 6C 27 B4 7F F6 88 6D 99 50 8E 3F DC 50
 73 B6 DA 58 83 CD 89 2E CF 58 0F 77 B9 BD FE 9B
 F2 CA 21 A0 DD 85 97 D7 4F 85 9F E4 C1 1C 88 94
 A6 AA BD 7C 54 5A 74 AB 28 1D BC 5E A3 50 C8 DF
 1E F7 6C 47 1D 8B 79 93 50 66 D5 7C DB 3C E6 24
 3E 9B 32 3E FE 10 94 DA B4 74 BB 6D 45 F1 6C 90
 9D D2 89 89 09 FE D3 2D 06 73 8D C4 E4 B0 F9 91
 D9 3D 21 00 D8 56 67 97 7E A4 5A AA 68 97 B9 EE
 7E B4 AA EB 6F A3 22 52 65 B1 A2 05 00 F2 B7 05
 A3 4E 9B 8B 5B 32 4C 6C AA 37 53 B7 78 2F 6F 20
 47 A1 CD 54 F4 AB 15 0B DB B3 BD 8A C3 4C 41 D1
 9B F7 89 7B F1 57 1F 30 0D 72 D4 F7 EE C7 99 BA
 7C 10 59 99 A7 90 35 B4 06 67 E6 8C 2F C5 30 6C
 19 6B E8 95 66 EC BD 72 F1 E2 52 16 17 04 64 90
 CD 58 BB 79 0F 90 D0 E3 BA 81 21 B5 9D D3 63 4D
 CD B4 51 49 A2 6E 67 9C 32 C8 C6 09 3E 07 93 B7
 D2 B8 18 AC E8 66 B9 9D 55 1C B9 1F 55 4A 0C 06
 F6 BF B4 2D 49 12 66 83 A2 55 F7 FA 37 9F FC EB
 E8 06 5F 4E 6C 80 1C BB E2 D2 57 89 14 57 B7 F0
 A6 ED 30 3E 11 0F 67 7F 0C C8 CD 7F C8 C0 E9 37
 A4 3A 4C A8 76 DD 67 1F 41 15 38 64 99 D3 37 AB
 A4 77 32 24 66 A6 DE EE 38 1D 9E C8 8D 0D 26 70
 1B 84 8E B2 88 DD FC 43 DB BB 61 60 37 0C A4 EB
 68 C1 64 36 42 41 9B A4 A3 CE 2E 11 40 10 51 EB
 7F 6A 71 E4 39 B0 97 C4 DD 48 C9 79 07 84 5C 3D
 94 4D 0A 48 84 A0 1F 32 1A 4F 6E 62 54 D8 C5 FE
 A6 09 A3 A6 2D E1 9F B1 A9 6A BC E4 B5 A8 70 18
 E5 0C F6 1B 65 C3 33 AB 1D F8 52 BE D1 D2 B8 F4
 91 6A E2 A4 A8 76 CC 6E A0 A7 56 9A BA AA 23 07
 29 A1 3A D0 FC B7 AB 4A D8 0E 95 C4 3D F2 6F 7B
 A3 A3 A5 58 54 A6 AE F9 03 9D B2 98 C3 AD A2 60
 EB A0 D0 89 E6 01 D3 70 55 AF 2D B8 A8 B0 66 AB
 F0 5B DE 6D 71 C4 36 0E B0 F4 A4 90 0A A6 6F BE
 DA A8 2C 53 64 C2 FF 66 D8 F6 D9 01 2D 5E FB 6D
 B6 AC A9 F8 62 78 B5 2F 10 B1 6E 5D 9A 3D 6B 4C
 8F EE 19 1E 84 E0 68 50 FE 57 3A 90 03 1E 99 8E
 5E 60 E7 A3 09 92 48 AC 45 8F 37 2A DE 5E 9F E9
 AF 2C 7C B8 42 F1 60 B3 25 E3 92 AD 17 CA 10 18
 DF 62 D4 52 B3 62 DB 38 6E 19 2B EB 53 A5 47 76
 F7 8C 12 C2 8F B1 E1 7D CA 71 D5 18 C6 20 FD 0F
 48 F8 57 97 7F 72 BD 33 21 F9 91 E3 57 C3 1D 9D
 1A 39 CE C7 C8 C8 DE 27 27 1D 13 4C 61 6E D3 4D
 86 0A 27 85 5E 05 97 10 F3 5B A9 55 48 DB CF 1E
 8D CF C0 A8 3A 46 C2 AE 12 3A 5E DB CF 65 B4 3E
 3C C8 96 A4 B9 B6 65 C5 77 B4 6B 3D 0C 2B 40 5F
 F9 FF CE 04 BA 2A 8F 77 4E 2F 53 6F E6 8C 15 15
 8A 58 56 09 F5 1C 86 58 0D 0E 28 B6 77 CA C0 9E
 BE 9D 17 5D 66 4D 08 73 E4 84 F3 EF 43 44 C8 1F
 42 FB 4D 95 0F CE 86 32 2B CA 3B 19 F4 4A EE 7F
 15 42 4D 63 D5 B2 8F 65 5E 0A A7 35 70 81 3E 37
 BA 2E 35 59 2F EB 56 66 23 D4 B1 CD 88 A8 65 91
 23 37 73 72 B9 E9 A0 F2 FD B1 77 CF 35 0A F8 2E
 DC A3 00 55 9E AD C3 E1 49 84 29 A3 11 D8 9C BF
 A1 62 2F EC CA 21 04 E0 03 C1 42 26 8C E0 50 79
 3A FB CA 87 D5 B9 D7 36 3A 68 CC 28 92 60 6D 19
 36 62 D7 64 61 36 B7 8D DD 95 69 92 43 D8 97 B4
 16 31 97 4E 7F B4 10 3B 6B 89 5F C0 38 CA 8A F2
 FB A5 C0 04 60 72 53 88 24 34 E6 45 80 7C BC 25
 E0 4C 77 A2 CE B2 2C CA 11 DA 49 39 16 F1 86 0E
 F1 A4 35 3A 2A D7 67 A5 E3 EE FB 24 9D 9A E1 81
 DB DC 3A 84 D9 FB A7 54 8A FF 68 BF C5 C1 56 55
 93 75 B9 2A E9 F9 EC C7 4A C6 DE 5A 4A 69 83 2A
 A9 F2 01 F8 68 C5 D7 C9 B3 24 69 77 AB 4B D1 86
 6A BC 4C 43 53 97 5E 60 FC 39 54 9D 70 5B E7 6D
 02 86 61 75 AD B6 7D 67 A5 9B 8D 64 90 8D 72 2F
 40 D8 7C B4 1A 13 BB A3 DA 78 64 5B 03 A0 91 7F
 9C 62 F3 AC 45 3C 23 89 2D 0A FF 87 DF 35 0C 5D
 83 3E 84 24 9A F1 DC D6 E4 D2 0B 37 50 88 22 D6
 C0 53 21 A6 90 D1 DB FB 7D D4 91 96 74 15 F7 43
 B2 FB 80 D0 3C 6B 60 62 A2 70 89 6F B2 43 97 B5
 70 5A 5C 47 32 56 FC A7 E5 11 D0 06 F9 E1 37 B7
 2D BC CC 1C 3E 82 F4 70 61 58 90 F8 39 6A 77 5D
 76 C1 A7 89 E2 2C 92 1D 82 68 4A F0 21 13 4C 67
 B8 A4 0C EA 98 1A 50 88 B5 15 E0 5E 96 BE 7A 08
 51 D6 C5 99 64 EF 98 DE 67 A5 F6 4D 0E 96 C4 A7
 E0 1D F6 57 E0 7F 2F 13 90 87 AF 45 25 8C 62 A3
 99 90 AA B9 D5 FE 07 2F 02 8E E2 37 42 1F 17 9E
 6A DB 0B D0 F8 E4 F0 5B CA 31 4C B8 82 C7 82 0D
 C3 76 F2 00 AB 42 BA 9F 5C 50 A2 BB 97 95 56 44
 F6 92 4D E2 61 E9 C4 E4 8A 1A FB D3 3E 0A A0 F5
 6F A7 08 45 34 3D CA ED 4B F4 52 C0 13 4B 07 FB
 12 06 2A 82 7B 93 C1 87 9D 71 DA F3 B7 C4 B1 F8
 8D 02 AF 83 83 80 FB 91 E4 45 21 91 CA 43 6E 79
 33 0C 49 4F FE 1E 7A 47 B3 54 7E 7A BC 6C 09 C2
 86 A6 2A DD 90 5C A2 23 81 39 70 3A 56 09 21 F5
 DB F7 F1 EB F5 60 FA 0D FA 8F 9A 63 A4 72 DC F8
 BF 41 58 97 16 EB 0C 00 05 26 86 86 F9 E7 D8 BA
 5A 5B BB 04 C8 10 CD F5 47 7F CA F1 6C F8 19 C3
 75 1C F9 AC 3F 58 EF 44 D7 17 82 13 62 6C 5A 38
 2A 31 2F AA 46 7E 51 C1 79 A9 E1 C4 D4 9D E3 DC
 82 8F 5C E3 EE 8F B9 CD E6 C5 B6 31 07 B2 6C F7
 EF 6D 07 8B 2E 18 58 23 4B 29 BA A6 48 BB 3D D3
 F7 8C 29 00 4F 7D 20 83 FD E5 8B 5C A2 D7 26 92
 F0 BB B0 71 AD 4D 6A FF 80 1B 33 03 41 FC 57 4B
 65 58 F3 EE E1 3E 3C 9E 62 55 53 D9 CE E3 2A 4D
 82 1C C8 DE C9 45 21 32 54 F0 A4 19 19 9B 9D F6
 BC 31 E3 8E 2D 16 9A 5E 1F 32 81 81 6F 74 05 AE
 89 78 0D 30 AE 87 D9 66 FF 42 CD D4 73 24 65 27
 9B 7C 36 EF 59 74 09 A6 32 6B 44 91 7C D9 7D 56
 1B E4 8F C5 87 00 79 A6 3D 1E 21 3F C5 D0 58 25
 EE 6B 24 D8 7F 77 66 32 C9 EE D5 F6 25 9A 8E ED
 3F 5F BA 1C 9E 1F D3 B0 2F 56 00 3A 64 B9 DF 08
 3A E9 29 20 03 83 AE 96 32 74 09 84 64 96 C0 16
 09 8B 16 17 EF A8 65 88 40 5B F2 BD 6F FE 10 79
 BD F1 F1 86 EA 6E 26 79 4F 3E 14 FC FD E7 CD 4E
 D4 A3 06 CA 2E 23 37 36 90 C1 04 14 63 DE 09 44
 57 5E 99 07 20 8E 53 21 E2 1D D6 CC D1 C9 09 23
 E4 F7 92 14 91 C8 78 52 00 01 B0 D3 C8 2C 4F 26
 74 EA B2 39 2C 62 25 44 29 D2 A0 AE 3D 65 9D F4
 14 99 EF 1B 09 CB 37 C6 E6 46 56 71 CD 7B 4B 82
 6C 96 9A EC A9 1D E3 F0 3A 59 04 DD C5 AB 0D C6
 17 06 96 2E C3 49 AD E8 F0 4C 7B 41 61 B0 D8 54
 E6 16 0D A7 B0 C2 BE 0A 54 10 79 3B BE EA D1 33
 F4 8B BB 66 1F 59 87 C0 7C 8B 73 19 AD 97 36 89
 65 C7 AF 48 DE A0 CC AE F8 79 3D EC 73 3C AB 3E
 45 ED B6 69 D0 61 56 6F 65 90 61 EF 2E 59 6E 98
 B1 C0 09 6B 01 3A 67 BC 09 09 9C 0C 96 C2 84 28
 C9 3B 09 51 84 A5 46 82 F6 DF 82 C9 0E 06 A7 64
 2B CF 5A A2 1D F0 BF D5 10 18 36 E1 A0 AF 17 F3
 3C 81 00 F2 48 A0 22 5C 66 13 35 7B 73 4E FB 8D
 E1 2E 9C FE 46 2F A2 11 38 3C E9 55 C4 19 19 D2
 A9 84 9C 8F B7 A6 71 3D A0 B5 FD AC D8 18 8E 22
 37 D5 D0 DF 96 4A 89 0E 00 27 B0 FE 66 EE F9 65
 93 F1 F4 8D 6C 17 4C 97 FE 56 BA 62 90 A5 EF 13
 9C E9 08 C4 49 C1 24 53 E9 84 C3 E8 86 B1 47 2D
 5D 37 1F 61 EE 7A 87 1D 74 D7 AC 49 12 37 76 DD
 5C C9 08 92 89 65 06 79 3B 89 47 09 59 2A 10 20
 69 87 CA 79 71 16 68 36 D6 5A BC C9 E0 06 BD 3A
 32 58 76 1D D0 06 BD 91 FE A9 D8 55 BF 92 37 5C
 24 AC D2 80 75 D4 D2 62 B0 FD 3F E9 16 34 28 75
 5D A1 A6 C5 9E C1 31 6C B8 1B FA 4E 60 7D B0 F5
 74 B7 6D 1F BF 6E 1E 13 57 94 51 52 90 5B 8E 7B
 90 35 78 46 5C 80 73 A4 48 AE 73 E3 9B E3 DF A9
 D0 3A BD BE DB D2 96 61 3B 0A 65 D0 41 C9 72 97
 BC 19 AA 7A F4 61 99 CF 0A 60 B3 FE 84 8B E9 89
 F8 8F 88 C9 A0 7C D5 31 4E 42 0C 5B 32 65 62 6C
 4C 5D 1C DA 2D 02 F1 10 17 F8 D6 B5 39 B6 C0 02
 CE 5F 47 85 89 ED AC 88 92 17 1D BF 60 3E 23 61
 AD 56 11 A8 86 D2 89 6C 03 95 7A 43 08 DD 8D CA
 C6 C1 60 4C DC 16 CA F4 BE DF C5 17 66 4E 66 A2
 65 CF 82 E7 1A B3 FD DF C7 12 8B 1C 82 45 A2 0E
 3E BF 77 C6 56 71 19 8E 12 45 34 6B 39 31 76 E6
 E7 85 88 96 B9 83 EF BF B5 B8 70 21 80 E8 BD DD
 65 DC 45 DF 2B 5D 6E C7 0A EC 6C 6A 40 61 37 98
 F9 34 86 1B CE 0E F3 0E 3A B7 58 C6 E3 D1 A1 2A
 3E 16 11 42 49 A9 71 4D 8F C4 BE ED BE D0 62 0E
 DB 7E BE 91 A3 EC 5F 42 BF D9 81 69 AD 65 7B 94
 4C EF 9B 13 28 0C 43 B5 3C 3A C5 25 8D 2A F6 54
 9B FA 92 3F F6 BB 5F C1 0F 6B D0 41 69 2B A9 85
 6C 3A FE 68 AC B3 A0 3B 9D 10 8A C2 51 17 61 74
 F6 8F 92 0D C0 7B AC EE 94 98 DE 0A 69 67 74 DF
 13 FD C4 5B EB A6 4C 70 66 42 00 CB 06 D6 3A 9E
 C0 42 08 D5 69 47 1A FF E8 64 DC 2F 50 12 76 BA
 85 18 ED C0 3D 98 1B C3 83 D2 AF 8B 10 47 C4 E5
 26 31 92 78 50 3A 75 1B F5 0A 61 80 52 25 5B A9
 51 3A FF 33 FF C2 9A CE 7A 9B C7 C3 F7 F9 C6 7D
 28 41 56 A9 FA 9C 21 F0 18 DF A3 96 4E 29 4A 30
 EF CA 96 81 CF 5D 68 D0 FC 29 6B 34 01 79 48 12
 85 95 EE 2A 87 1B 4E EF E5 39 F7 62 C9 EA 32 AE
 D4 B8 0F CC DB 14 99 F5 37 E4 43 A3 40 98 08 E0
 06 F6 0E 40 D4 13 01 94 FD 9A 66 83 77 7C 06 71
 AC C6 C6 2E 4E 3C 18 C1 27 47 04 7E 13 35 B3 37
 57 0C 7A 18 56 AA 28 69 19 65 15 63 7B 02 84 49
 FD 47 F1 71 8C 28 D1 E8 59 BA 05 4B 34 70 B0 51
 8D 59 6C 9D E8 61 73 C1 B5 1F FD 82 72 90 4A B7
 96 A4 A5 AB D6 05 06 6B 0D BE 0B 0F 86 8D 6F 54
 A8 BC 03 5D 10 90 33 E3 29 92 8F 17 A9 D2 7E FB
 5F D4 41 22 0C DA B4 3E A1 6A B6 55 7B 08 DE B9
 C7 FA 25 D5 88 C4 EB BC 92 6A 4D 68 F5 B4 B6 16
 61 8A 0E 35 8A D0 4B 30 A0 4D 6B 90 55 77 50 93
 CC A4 47 F1 49 1F 57 A2 A4 A7 87 78 F8 00 AF 84
 87 32 5F 72 E1 F5 C4 C3 FF D7 AD 22 0F 1E 83 42
 CE B9 14 42 56 E0 A7 4A 21 B3 DC BF EE 3B 1A D0
 EF 0F 6E 07 72 CE CD DD 21 8A 4B 02 56 3A A8 F6
 86 BC 1C 2B C6 A0 38 D6 7D 0E 92 3B 1F AC 48 84
 1D 13 EB 3B 13 FE 6B 89 14 E6 43 FF 17 A8 17 B1
 3B 6A 0B EC 49 52 CC 5E 95 21 C1 7D 74 D5 66 13
 20 4C 07 1F EC 08 97 E8 C5 5D 17 1F 86 92 48 ED
 B0 C5 16 39 51 24 DC CB 21 6C 0C FE DB 11 A5 72
 8A 81 C7 EA BF 75 F2 B8 1F 92 D9 21 6A B6 F6 D5
 B6 4E 63 CF 12 52 30 47 9B 75 E6 C6 EC 08 F1 00
 4C 2B C1 C0 D2 89 F2 E0 41 4C DE 87 8B 08 CC 9C
 49 3E D6 6C 93 40 13 33 AE 77 E9 54 66 15 D1 05
 AF 2D 29 B1 05 AE DC DF 17 E7 24 1D 0F 10 6D 79
 DA 32 16 44 79 56 24 27 4D 2C 4D 3B E7 55 A8 66
 29 97 AF FC 08 D9 24 5E BA 3E C5 03 FC A3 2F 3B
 BD 8F 96 9A D4 F6 B5 3B DB 4C 93 E8 92 6A 64 15
 4D 5A FE 7F 1D 17 2A BC C5 F4 FB 17 F1 7D EB 10
 67 73 11 72 71 68 2B F3 5C 9D 33 AE 18 18 4B 96
 E8 4E 3C E1 2E 6D 39 6B AD 53 FC 25 3A E5 BF 2F
 4E 90 DB 5B DB 2F 68 E6 93 47 BF 87 3C 50 36 EE
 88 E5 43 EB E8 AE C6 78 1F 68 FA 82 B2 C3 6E CB
 69 FD 89 CB 52 26 19 41 7E 77 0C 04 2B BB D2 AE
 D5 5C 60 80 4E 78 D8 55 73 4F 13 59 79 4B 20 0A
 E7 35 F7 42 05 D6 F5 E0 70 82 91 86 74 27 00 C4
 85 90 5D 3D 2D FE 90 C4 11 44 C9 DA 96 9C 67 2F
 CA 27 75 73 E2 F1 2E 7C B5 BC 5A 3F 05 F5 60 5A
 54 83 7F DE 1F 53 4F 41 19 1F 51 3F 65 73 47 2B
 1C B0 14 BF CB 1D C8 20 98 89 29 2E AD 00 03 45
 4C 7E 39 73 09 69 36 AB E3 6F 0C 23 9A B7 F4 FB
 22 6C 21 93 81 BE A5 BA 34 FF 01 CF 90 28 31 C2
 ED 8B B2 16 D0 40 15 4A E8 E2 C0 55 53 73 8D 76
 CE 0C 79 4C 39 25 3D FE F5 4D 00 8C 4F 09 47 AE
 0C F4 7B C0 9B B8 FC 5A 4E AC 03 90 0D 87 1F A1
 EC 3A 10 34 C0 FF 9B D8 1D D3 47 7F 37 DA B3 DD
 F8 15 11 61 A8 FE 74 2C 68 72 43 33 AC CA 3F AC
 2C D9 CB 89 DE E3 97 5E 34 A0 55 14 EF 3E 0C B2
 A1 B7 91 35 80 E9 72 FE 9C 8E 40 13 A2 BD D2 B8
 47 64 01 85 E3 3D 72 C5 5C A9 C8 D5 DB 47 31 98
 AE 7D 30 9B C3 85 1C AF D1 ED 8B 81 A5 6A 4B B4
 A4 FB BA BE 0C 54 F3 A3 33 37 5B D9 0B B6 36 B5
 92 F7 85 98 DC D8 67 B2 60 53 6D E5 34 3D C1 5F
 0F DB 18 FC AF 6A 6A 96 3B 3F 96 B5 01 B6 53 C4
 DA 2E BE 30 AF FD A6 43 E4 44 E4 D4 67 C8 B5 5C
 41 C2 AF 5C 5A A8 62 4B 8D B4 2E 69 11 5D 36 E5
 E3 C5 95 A4 B5 2C C8 F5 C1 BF 14 02 6F C9 05 57
 06 08 80 E3 D5 CD 52 3C 6B BD 03 ED 57 26 1C 0F
 2C 92 A1 47 FC 3D 70 66 B9 D6 35 12 14 DE AC 14
 E3 21 23 29 C4 14 58 1E F8 13 55 AF 21 53 CC 3B
 28 5E 57 B3 20 54 CF 5E C0 36 39 96 82 17 2D 95
 B5 88 65 19 85 F3 42 C5 FA D9 03 2A 3A 31 72 6C
 EC 90 41 81 05 0B 10 4D A3 E2 DF C7 69 AD F9 63
 1D 80 6D A6 FB AD 55 0C 98 3B AF BA C8 33 16 25
 61 5C 9E 6F 19 33 AF CC FB 23 5A 2F B1 FC FE D6
 59 27 A9 34 93 18 18 24 3C ED D2 25 56 B1 C7 A7
 8B 48 61 20 81 5A FE DC 52 AC 6D E8 3B 54 7C 8E
 D4 ED 1A D2 4A 2B C4 C0 D7 3F 12 F6 90 72 65 27
 5A 2C 35 19 32 6F AA D9 6C 66 F9 94 78 9A 2C FA
 C8 DF 2C AD E3 6B 32 2B 4A B9 20 14 31 E4 F8 E6
 C2 E6 FE 6D EA 12 A4 2D 8A D9 9C 4C 74 85 1F 57
 7A BA 4D 89 18 78 E1 C6 E8 B8 FB C8 16 A3 09 FC
 A9 9A B8 09 6C C6 DA B2 2D C3 8C D3 C9 A5 BF 81
 21 A8 01 DC 8D 5E 3F 20 BF A0 11 14 EE 6B E0 A4
 EA 19 58 04 B9 AF 5F 8B CF B2 34 86 71 8A D5 E0
 AD B5 27 67 9D AD 78 F5 7B 8F 2A 03 2D 94 3F C6
 99 59 0D F5 73 4F 3E 5D 75 8B E1 F5 71 E8 6A 0B
 C1 11 9F 13 28 9E ED 70 68 A9 FF 69 C5 EF BE E5
 32 B5 02 39 3E DB 5C A9 58 6B 7F AE B3 65 3C 2C
 0E 9F 01 CD CF 0B E7 28 04 21 E2 48 DD D9 4B 3C
 75 94 59 69 49 B0 7B 1B D9 1B BF CE 8A 19 6E A2
 0B FE 6A 81 CF 51 8B 03 91 F3 51 28 BE D8 73 35
 A3 31 C0 90 7F CC 1A CD E9 EC 03 98 88 3C 63 07
 95 80 A0 2E CE EA BD 6D 59 21 2F B4 3C F3 16 EF
 58 BB 24 C1 1B 34 3A FD 81 2C 1D D4 16 B2 90 21
 0B 40 72 82 70 6F 80 3E 22 17 92 BA 47 DA 2A 45
 68 24 3F 8E 9F 8A 1F 1E 2A 35 48 FB E8 7D C1 4A
 8A A5 05 A3 6C 8E 02 CC 66 31 DC 3E 3D DE 42 89
 27 EA 68 C7 40 DA 10 AF D9 5A 7E 1A 1C CF 2B E9
 62 89 6B 97 CF 50 1B D1 7F DF 6D 57 A5 30 D5 56
 35 37 DA 9A 46 E0 2E 91 CA 92 6D 2A 94 49 76 84
 56 0D 9C 5C 18 01 62 D5 6C 64 3A BE 06 6F 9A 56
 3B 8F 8B 40 4B 77 57 56 DF CC 89 69 60 EE CF CF
 0C 3C C8 F4 5D 28 69 2D BF 0C 8E EB 0F 64 07 2C
 5D E3 0F 2D B2 3E C3 71 21 72 9D EC D1 F8 C9 B1
 59 30 A6 1B 01 EF E7 89 AF 4C 6A F1 63 25 CF 50
 95 CE 00 B6 3D 6D 05 5B D1 0A AD 8F 6B 8C 01 FB
 DF 84 AD FB 1B 9B 22 F1 9F C7 55 99 94 B6 E0 6E
 D9 5B CD 01 9B 20 E8 FF 4A 56 D2 07 7E B9 85 20
 08 64 4A 37 A7 A8 CF 0F 6B D8 8D 5E C5 6E C8 DD
 A4 1A 3D BE 5D 73 15 49 FE 6E 02 42 12 17 60 B5
 8D CA 94 A3 36 4C 27 F4 86 BB 6A BF F0 84 6E 18
 73 7C C1 F4 E0 7D FB 60 C8 B5 C9 2B A5 28 D8 2C
 3D E2 13 A2 2C C1 27 27 82 A2 FD 8F 3B 92 CF DD
 D6 77 D3 EF 20 16 18 BF F9 68 CB B1 27 D7 84 B6
 40 A8 78 BA 87 ED 46 65 DF CC 03 12 AA 48 79 49
 8D 5A C3 8A EC C5 E1 23 27 57 C0 BC 74 B4 3C 15
 B7 9D 92 31 BF BB 6B BE BA 03 D0 4B B3 95 7A D8
 39 13 61 6F 82 0F 03 B1 F9 68 35 AB 2A EC A0 AC
 F4 FC D0 9C 6B 7A 5E 2F 29 EB 44 3B 86 39 D3 FA
 E8 7A 76 74 33 CB F6 7E 48 E0 10 CF 21 88 70 09
 D7 AA 3D 2F 11 5F 3B D0 41 C4 20 0E 33 AC 56 6B
 71 B6 B3 7C 4A AF 23 6F D9 94 90 45 80 77 5D 44
 AC 63 15 E9 AF 60 70 58 9D A1 85 71 B6 BD 6D DC
 91 DF 98 25 10 87 EA 12 D0 25 39 7C 97 60 D4 ED
 B8 8F F6 05 3C A6 07 8E 67 64 BB 77 7E 20 C0 85
 5A F3 09 37 97 9B AF 1E F6 78 E0 A3 46 4D B2 84
 CA E6 24 3F DB DB BE 68 FD 42 2A 3E 2F 4F C7 43
 31 AE A2 A6 73 36 AF 1E 9C FB 76 20 78 B6 80 2B
 01 E8 D6 40 C6 6B C3 57 D1 E8 CD F0 DD B6 AB BB
 10 2F 35 39 68 A3 F2 17 93 39 3E 81 D9 4F 21 61
 4C 6C 3E E6 21 6E 42 12 A1 F8 19 CE 0E A4 9C A2
 00 61 D2 79 43 5C 5C 6B 85 6F 67 2B 1F E7 B6 B5
 8A 98 62 28 8B EB 7C F6 9C EF A4 C3 5F 8F 16 C0
 A9 2A D7 DF 2E E1 F4 4A 88 8F 14 3A 56 A8 ED AA
 D3 50 61 C6 22 8B A6 DB 1D D8 16 5A 90 4E 99 A9
 0C 51 D3 1F 17 24 C7 5C B5 FD 9C 73 E8 88 F5 E0
 95 31 10 BB 03 BC AF 4F BC CB 76 2B A5 B0 16 AD
 51 65 82 6D AD 4D 8D 30 78 F8 C7 6D B6 D5 BB 76
 DD 8F 96 0C 93 3A 8C 27 A2 A9 8E 94 C9 BB AD 08
 BC 10 AD 96 19 18 A8 4A 73 57 72 08 00 6F 76 61
 A5 61 CD 82 EB B2 98 1F 42 02 4D BB F5 E5 FA 60
 5C 5D 06 B5 B7 65 64 09 4F D8 01 10 9F 87 F6 24
 71 B2 E2 23 BB A3 8F C0 CC EC B1 93 F6 F8 75 8B
 F2 D3 67 61 DC E5 8C 22 B3 9A 98 96 12 E8 58 24
 7D 0B 8C B5 06 71 4E E3 67 D8 5D EF C6 50 F6 DC
 32 52 17 49 53 39 E0 10 3F F4 27 EB 36 D5 B0 B9
 82 86 73 59 92 41 CD 58 F5 6D 1B 9A 81 8E E5 D0
 33 D9 0E 7F 13 21 D5 07 E1 41 A9 20 7B 34 0A FD
 B0 95 B0 3D 6A A5 28 AF 18 26 68 4A 9D 2A B8 91
 45 F7 57 11 09 24 B5 42 2D 10 46 AF CC BE BA 57
 28 8E CE D7 D1 7D CE 95 BC C0 2C B7 C7 80 81 B7
 C1 37 AA 96 01 2C 2F 12 D4 1F 5C 02 5E 7A 74 F7
 21 5A C8 FC 2F 1D 22 6A C7 D5 3F DB 22 B9 7B 97
 78 F8 63 4F D2 4C 93 21 EA C6 2C 12 D8 F0 41 34
 46 02 B5 CC 6A 5E 98 DA 70 D2 8B 08 2F ED 9D 1F
 A1 7B 17 AF DA AA DA 01 0F BE 83 B1 0B 01 0B 8C
 80 91 7D 28 E7 CE BF B3 12 6C 97 A2 69 41 CC 22
 30 80 6F 42 F3 27 1C 03 0A 09 C0 07 C1 17 F7 30
 64 5C 0C 36 3D 04 32 4E D8 3F B8 AC 35 BB DB E7
 64 65 B6 5D D7 80 0E 8F 8E 29 3B 1B 45 D7 AD 25
 06 71 E2 59 B5 EB 25 1E B1 74 11 09 7E 0B DE 74
 6D B2 F0 CF 17 2A DC 7C DD 0E 41 18 15 8D A1 86
 07 20 35 71 13 24 5B 98 CC D1 12 7C D7 8A E1 F3
 38 A9 EB 10 C6 96 EC 8F A3 D9 55 E2 E4 F6 83 5D
 9C DF E7 29 04 4D FF A1 21 20 00 40 BE DB D4 03
 25 6D BE 3D BB 82 71 1D 5B 03 32 E2 99 D6 46 C2
 EA B2 2F 17 63 0E 2C 41 44 11 56 E8 9A 30 74 93
 9B 10 17 38 EF AA C1 59 79 C7 88 73 BC 13 BB 39
 DA 4F D7 49 7C 04 AB C7 95 7C 33 86 14 58 0A 62
 DD F4 60 CE CB 7F 87 63 AF FA DA 0D 43 1C 5B E3
 88 2F FF 79 C4 F7 BB 43 FF 10 FF E7 74 86 2C 87
 F9 C0 0E 91 37 E5 29 82 4C AC 47 68 43 F7 42 FE
 FA 72 82 43 F4 F6 E9 B4 DA 27 F8 12 F1 C1 59 17
 19 C1 98 41 DB 38 5F F9 5A 49 28 03 07 2E 91 A5
 22 6C 13 FF F9 E8 A2 24 4C E6 33 8A D3 32 3E CF
 A5 7B 78 C4 2E 0F 94 02 B0 19 7F 87 8F 73 E8 6D
 72 6E B7 0C D1 35 BB CE DF C0 A0 86 A5 1F FC 9E
 FE A0 62 52 61 D6 79 8C 39 9B D4 EB B7 E9 3E 35
 DA 17 8A E9 39 CC 71 65 C1 0C BB 6B AB 63 A9 E3
 41 C7 C4 AF CD FF 79 71 9A E1 FD 55 AC 2B 38 78
 03 79 52 08 01 1A D1 EF CC 71 B6 0D 68 F3 7F 9A
 0E F8 D6 0B 87 28 A4 6B B2 E4 D5 00 C6 30 A6 D7
 43 0A DD DF 04 A4 D9 EB DB E0 8B D7 02 93 B7 CB
 96 EA A5 F0 35 03 46 41 CF 51 A8 C9 D4 99 7C F8
 ED B0 23 49 2E E2 9D 32 55 28 38 0C C2 45 91 6A
 E8 39 49 29 57 0F 8C 83 64 D8 F4 C6 91 F7 3C 55
 93 3B 42 BF CB 8C 23 09 48 23 03 60 0F C7 A3 A5
 0A 20 9C 46 10 0A E0 90 0D 61 2C 8E D2 E9 9E 8B
 47 E3 6A 87 59 48 EA 9E DC 33 3F 23 68 D7 8B D0
 3F 8A 8C 8C A7 24 2B 32 D3 27 DF 35 D0 9A BA FB
 B9 BE 52 F0 07 72 1C F5 7D 30 36 30 68 57 B0 AC
 DB 05 08 D6 58 71 2D E3 AB 56 E3 32 61 79 64 CB
 55 40 D1 43 FA 8F F4 7B 1C 60 CB 9F 2C 21 71 5B
 05 BC 05 DA 7D 60 08 F5 F8 33 F3 1F 2A A8 1A 16
 1D 8D E9 13 6F F4 48 DF 5E D5 3F F3 C7 DB 53 E9
 FE 45 84 A6 96 58 C1 F4 EC 2B CB 00 CD D2 69 7F
 37 2E 21 4B 40 F9 9D A6 B2 A1 19 AE 93 B5 B6 FB
 B8 4A 00 2F B0 9C 35 40 78 51 F5 0D 3D 31 10 AD
 8C F2 84 72 E6 EA 1C E2 F9 6A 2E 65 30 46 4A 40
 89 B6 5B 72 FA 14 43 5C 63 DE 75 C7 C1 0C 4E AD
 38 CA D5 A3 14 C4 D7 89 89 5F 91 8E 75 71 3C F9
 43 82 4D C5 2B 0A D5 52 CB 6E F5 12 8C 89 FE E2
 08 76 0F B6 BC 60 5D DF 0B FC 94 41 A5 F7 39 14
 4A A1 A8 E1 69 46 24 23 67 99 4C 5F 8D 90 D3 81
 5D 15 9D CF 7F E1 BB AF E6 86 2E 23 9A 3A 83 AE
 C7 5E 3F 84 18 59 49 EB FA C1 6C D1 EA 9E 47 7D
 20 8D A1 FD 08 78 C0 E5 12 42 C7 60 24 54 86 98
 9E BD 06 91 B4 A1 E1 F1 C1 FB 2B D0 3A 82 7D 73
 76 C4 ED 82 AA B6 C2 DE 78 F7 44 CA 04 AB 79 76
 35 E8 03 13 8D E8 BA 1E 5D 16 5D 24 C8 66 A8 B7
 8F E2 F9 3D B5 50 71 85 07 7C FA 04 D1 89 A0 D4
 ED EB 7E 66 BC 4D 20 2B E2 D7 54 54 92 57 AA 4C
 B9 6D 21 D7 15 1D 84 40 DC AB CA 3D B7 A8 3A 9A
 83 04 4D 21 75 EF 62 AF 68 DB 12 6B D3 79 D4 3D
 12 D0 05 8F ED 44 8F 3C FF 66 A4 F8 6B FE E5 55
 FB 90 83 71 7D A0 F2 2A 4D 01 9E E7 50 77 2A 15
 2D F4 47 FB E9 F0 D0 05 85 ED 31 1D 4C 02 97 21
 3F BF E7 0E CC 7E F1 DB 1A CF 88 5D C7 11 52 EF
 52 B1 BD 1D 9C CF 79 8A 62 50 96 68 42 80 8D EE
 73 30 3F 42 BA 7E DA DA D2 44 9C 2C 3F 74 96 A1
 E7 00 D2 79 29 AA A8 43 6F 1E 7F DA B2 D9 52 CD
 47 FE C8 81 B1 A6 B6 85 DC 21 80 16 1C A9 2D 11
 19 64 8B 6E 30 A9 9E 48 2A C3 52 FB 5E AD B8 B1
 8A 96 0D 7F 86 FE 39 1A 93 DA 53 22 BB 32 23 62
 96 EB DC 9C D5 C3 06 8D 19 C3 55 7A A7 BA 19 44
 CA 5C 01 A7 96 35 4D 55 67 36 69 D9 B9 5D DB 94
 44 83 8D D5 40 F3 69 34 C3 3C 13 EB 9F F2 66 95
 F5 59 31 D1 BF 67 C3 E1 53 15 32 5B E9 E1 1C 1E
 B1 9C D8 D4 1D 8F 47 FD C5 E0 7B E5 BD 8A 20 0C
 87 C7 F2 4E EF 4A 28 CA EF 56 37 26 1E 59 B2 42
 67 08 EA B7 B7 19 82 90 32 B9 80 73 DD 12 5F F9
 8F 19 7E F8 05 5C 47 C1 C8 91 1A 52 E2 74 7C E6
 02 5E 0C 45 6F 3A 3A 06 1C A5 D4 50 76 1B B1 40
 88 58 3D A2 29 DD F2 E0 26 B4 E3 7A 7E D6 98 56
 5A B2 AB C7 85 8E C9 50 B2 A2 FB 85 2B 26 54 1A
 C6 A5 9C C1 9C F4 26 09 EA 72 EF D7 C8 9C 07 42
 B0 07 FB A6 37 EF DB 72 74 88 54 4C D3 5E D2 41
 05 F0 0D BA DA 37 6A BB 0E 9E 9B 97 9B 7B D9 82
 9C F1 31 1C 27 A1 07 EB 0B 52 0D 3B F3 70 9C 3D
 0B DF 41 47 2D 4C D7 0E 9C 3F A1 32 0A B3 13 CE
 48 E4 77 EA 2B 82 C6 78 2A 39 73 1C 58 CE 4F A9
 6A 28 A3 FB 8C 0E A6 F8 A0 52 FB 23 7E 86 00 44
 3E A0 6C B2 EC 0D 29 2C 6A 02 29 C2 A8 53 DD 96
 48 A0 7E EA CA 49 04 14 B2 D2 CC 04 56 1F 9E 60
 EC 4C 0A 03 40 48 AD 55 6A 72 B4 91 E9 08 2D AA
 BA D5 36 23 11 47 E1 C0 CE 33 F4 A6 4C 06 7B DC
 43 EA 14 13 33 47 CD FF 19 16 51 0B 4A A1 92 EB
 82 B2 A4 37 3D 3D E0 A5 BC 9F A4 BC 69 82 8E 81
 E8 A1 2D C3 74 08 17 12 87 71 00 D8 EF EF 00 79
 6F EF 68 AD FA 95 BD 55 72 C4 14 B3 5D 1E 84 1F
 B8 0F B6 12 22 54 D9 BB 17 62 23 5A C5 08 65 07
 A2 64 0E F7 1D 1C B4 E4 65 19 20 D7 56 DF B2 8F
 47 AD C4 AF 9D 4D 45 1C 71 AF 14 A9 0D 3A D5 53
 2A 98 25 1C 46 A7 87 F4 A9 B0 CE D2 88 ED E6 3E
 49 39 7D B5 FB CA E2 EA 46 FC A1 60 68 D7 0A ED
 44 08 07 2B E3 B5 C0 CB A5 28 A2 1D 5E C7 8E 92
 F7 56 26 F8 6E BB F4 4B F9 F2 27 16 73 E2 CA 49
 9E 80 19 46 B1 89 32 AA 8B 2A 4A 30 F2 BA 26 0C
 94 E7 76 B8 8A ED 2D 51 D7 75 9A D1 50 8D E8 0A
 ED CA F1 AA BE 8C 22 3D 97 70 3F CA 65 BB 2A 52
 14 CD 6C 73 71 A4 C9 57 AB EB EB 21 57 3B 7D 5A
 F8 B3 9C EC 39 F9 4E 53 61 31 7F F5 12 6D 28 C0
 80 BE 42 B4 41 13 B1 BF 2A 69 55 45 25 47 13 21
 99 6B FA A2 D0 20 FD 0C 09 EA AB 75 F6 8A 11 9B
 76 F9 7F D1 D8 05 49 86 79 06 49 9D 01 86 7F 9B
 9E FA 98 F5 05 0B F7 B5 EF 66 CE 08 FA 37 38 B0
 AF 44 12 02 50 D1 67 10 08 8A EC A5 F4 E1 33 7C
 D0 D7 7B 93 43 9F 1B 6E 03 C9 F5 AC 15 72 89 26
 0D 31 32 F6 CD 27 AB 4D 42 BE C9 37 98 59 E1 CC
 20 06 AB 60 61 D0 FA 20 B5 ED 14 52 E7 55 9D 5C
 4F 4D 8E 74 23 C3 39 9F B1 99 54 EE CF CC C6 DD
 71 5C 5E 73 34 F8 AB CC DF AD 0A 74 F1 A3 32 96
 ED 16 62 CE 45 01 10 DB AB E1 0F 02 95 2E 20 E3
 7C 80 A9 C4 E4 27 33 39 57 EB F3 51 10 69 F0 C3
 B6 85 EA 50 10 F3 AB F4 F9 76 D6 C3 8C 87 D5 EA
 61 9E 24 D6 28 2D B1 6B 13 00 91 FD B5 7A C9 1C
 E1 4F E8 D1 B2 BD 7D 23 D7 79 E1 09 76 52 BF FA
 A1 9A A9 46 82 EA AC BB F3 56 D8 20 B1 9E 53 71
 9B 2C 7F 24 0D E3 20 DF 28 22 A3 FA 03 80 A5 3A
 8B 05 AD AD 3F 6A 68 66 74 50 07 BC 13 C3 74 78
 51 3D 83 F2 EC 96 56 11 48 2B AA E5 E1 64 60 7B
 3D DE B1 FE 9E 58 CA 49 C5 4E 78 CE 91 70 A8 60
 C1 43 D7 CD AF 6D AC FD E0 B7 E3 5A B6 11 17 2D
 59 A1 CF 05 BB 5E 88 EA 9C A1 02 F4 9E DC 3B FD
 37 D6 01 59 2C 8E 82 4D 46 1C 71 6B DC D1 04 64
 38 66 2A C4 85 44 25 98 CC 7B 1C 14 AF 24 0F E0
 8B 24 34 2D EC 3A 05 A4 62 E0 22 07 5C 37 35 5F
 1F EC 6F B7 8C 31 BA 2F 7A 99 C0 B2 F7 25 E8 D3
 09 B5 C7 55 CD 37 64 B1 55 15 A4 B7 23 D4 B0 70
 BD 9D A1 4C D6 E0 05 A0 4A 74 66 8C 9B 3B 26 F0
 A0 99 98 62 DD 49 AE 4C 42 9D 2B 2A B2 95 F2 AD
 B8 FD 1E A1 55 5A D3 FA 83 BE 32 E0 41 23 F2 2E
 67 AA E8 94 33 7F 59 A7 15 82 54 6F E2 45 8A 1D
 F7 EA 92 E9 9C 72 C2 DA 4A DF 1B 86 36 A4 18 8E
 FB E7 E9 14 76 82 F3 5F A2 91 4D B8 94 2E 10 27
 94 06 07 39 28 E6 06 F3 EA 2B 6A CE EC DD 30 18
 F2 54 61 01 42 51 96 AE 88 58 B6 71 B0 6D DA BC
 D9 7B 9A E9 61 C4 27 18 A9 1A A9 3F CF 3B BB 7F
 A2 F1 56 10 3D C5 12 F3 44 25 82 BD 4B 3C 47 49
 8A 38 55 A5 2E 72 A5 75 0F 73 75 6A 02 E3 02 52
 57 39 04 0A 58 97 A9 7B 6B 92 F0 C9 A6 FA F3 78
 11 FE D8 03 7C EF 6A 26 CB 0E 03 5A 27 64 B0 58
 66 80 4F 16 B6 68 21 E5 16 D3 83 0C 75 16 09 C4
 05 53 50 BC EB CB 73 03 DF 42 54 2A AE DB 85 07
 A0 DC AE 93 43 C3 1C BF F4 A6 55 8A F4 57 D7 79
 51 B2 3A CB D0 D5 0D DA 2A 03 70 1A 11 0D E2 14
 30 3B 0C C9 33 7F B3 34 86 02 41 63 27 45 3E A7
 E3 16 77 2C 63 20 9D ED 9E 5F 0A AE CC 33 99 68
 7E D0 A0 06 37 92 6C 6C 29 D3 F2 C7 B4 DD A9 F3
 C7 8A 03 B5 FE 43 47 12 89 B3 93 5A C9 1B CD 83
 45 EE 01 0C 6E C5 95 34 CD ED 19 04 92 B4 61 3A
 EB 6C 7D B8 03 50 3A 35 29 93 04 EA 7F 46 67 C8
 E1 79 4C B2 F1 D7 2B 40 B3 3B F6 F1 3C 0D C0 AE
 CB 75 57 EF D6 30 F3 34 5B 7C 39 E8 78 EE A0 25
 C4 A3 07 45 EC 11 F8 AA 74 6A 7F 4A B0 09 F5 CB
 B7 B2 35 E3 B1 51 37 3D 1F E5 24 A8 D0 EE 81 62
 DD 65 DC 3F 90 74 36 96 CF 95 1E 81 5E B9 F3 7E
 DE AC 2D CE 1F 35 71 85 A9 58 B0 33 20 6E 0B 01
 35 FE A6 C2 54 71 1C F7 25 FB 33 7C 69 04 6D EC
 AC 6B 20 A4 51 2F FE 1C BA 90 EB 49 A1 44 32 8E
 F7 20 53 05 96 11 8D 74 7D 77 E8 67 F5 A4 6F 4A
 5E 7B 64 C9 1E 1C 2B 33 23 D5 0C A9 DF 56 C1 B1
 1E 9F 53 E7 1F 7A 64 2D 87 05 8A B4 81 52 BA 6B
 66 AA 0F FD 60 A3 CF B4 82 77 68 06 F7 20 D7 24
 2F AD 0D 77 2D 82 18 ED D6 F7 07 A7 ED 1D C4 0C
 4D 79 72 27 15 D3 B2 48 52 9D 40 79 60 D8 9E 5D
 53 39 52 FE AD 4D E5 C9 4D 18 66 CD B3 4D 1F 8B
 DA 60 65 C9 65 93 FE 6F B9 A3 9C F6 33 4D 1A 99
 06 C0 79 3D A8 A4 DD 0D FA 9A 4B 12 70 3A 47 D3
 EA 4C 07 E1 A8 4A 07 26 FE B3 52 31 97 0C C8 D3
 A8 E4 0F 3F 7C 70 10 44 4F C7 A1 9D 5E F1 26 AE
 94 40 74 5C 81 43 B4 4F 53 0D AD D5 46 D5 88 39
 63 4A BD 4B D5 DF 7F 4B 43 78 71 AE A5 16 62 61
 63 8A 14 80 C6 A9 AA 7E 0E 87 64 90 D7 58 DA 14
 AC 4A 84 19 08 82 E2 D4 83 D6 C4 8E D8 69 12 52
 8D 8B 3C 32 A6 7F 06 FF 01 9E A5 89 2E EF C1 FF
 E3 88 8D 81 56 78 5D 0E 51 75 48 72 76 84 7F 82
 5E 0A D2 A4 86 19 B4 17 CA B8 A1 09 B8 0A B0 FA
 F8 F4 A6 B5 3E F9 8A C7 96 FC 50 53 70 9A 7A 61
 DA 09 3A 2B E8 14 E1 A0 B9 14 37 28 04 0F 70 19
 63 5D 24 80 31 47 81 C6 FA 46 F8 1A 06 83 8A 41
 2D 68 21 5B E1 74 1B FD 25 0B 37 F4 E4 44 E6 F8
 07 6D B3 62 54 43 F1 83 9B BD 04 A7 79 B0 03 4D
 DC 6B D9 70 B7 4E D4 46 F8 03 D7 42 C1 BD 9F A4
 73 12 BA 01 6B D4 6C 40 B6 8F BF 2B 94 13 9D DE
 AC 65 B8 F0 27 75 8B FE F1 2A 97 7F 39 1E 7F 2E
 1F 7E AB CE C7 25 30 AD 76 48 4A C8 56 DD D2 A1
 D7 9F 07 4D D8 37 C8 85 23 C7 8B 53 6D F5 B0 4C
 1C 3D 79 0D DB FD 31 73 E7 E1 37 C0 E3 EE DB F7
 22 40 C2 27 5D 66 82 15 6C EC 6F A3 6A AC 32 0E
 51 D0 FE CF D0 96 5A 73 F6 77 DD 2F 12 79 9F 11
 4F 23 CB 27 A1 36 10 60 8E 7D 53 45 20 30 8F B3
 3A FC 82 A0 1F 76 2E 06 2D E7 E6 87 6A 7A D1 4F
 05 F3 A4 56 B5 62 60 3D 0E 9D B6 AD 0A 36 94 C6
 26 E9 6E 17 21 E5 46 64 D3 3F 41 95 6C 56 11 5C
 D7 15 2D 17 B6 78 60 15 F8 E4 29 BD 62 26 92 E1
 B7 A5 A9 74 B0 BE 16 99 E2 05 52 04 AB 0C B9 18
 4F C6 3D 49 50 BD C5 BD 61 2C A9 FA 0F 07 4E 45
 74 D4 6E 71 00 28 DD 54 8D 6B A5 61 59 65 22 74
 6D 9A 16 88 70 E7 00 D7 F1 A8 AD 2F 61 7B B5 F1
 40 6A CE 27 D2 4C 85 92 3F B1 75 9B E5 B0 D4 45
 91 E4 F6 39 64 B6 B3 62 B8 0F 51 97 50 99 AE EC
 34 DB 01 F4 C0 57 4D 81 27 2A E5 2A DE A7 71 90
 37 C6 4E 75 99 F7 70 B5 AD 6E B2 09 A6 04 92 28
 61 E8 60 B3 79 49 79 08 A7 9F 0D C6 37 01 94 2A
 5C A4 D4 CB A5 BC 21 57 12 83 74 09 10 5D B9 AA
 C0 CD 47 D9 7D B3 9F 5A ED CA C5 E0 36 58 DC 85
 E0 A2 E6 A3 1B 8B 6B 1C EB 1E 0E 76 D4 AF 77 7F
 2A 9F AF DC C0 DE 3D 33 D1 2F 97 7D A9 33 C6 B2
 98 F7 1F 24 F6 5E 05 7E E5 96 86 2F C4 C1 10 A3
 AD B6 F8 D2 A8 39 4A E1 60 00 BA 89 59 2E 53 30
 70 AA 41 D2 DF 80 C9 95 48 3A CA 7F 52 06 E5 64
 EA 9B 77 DD E6 66 26 C8 FA 80 BC A0 EC 85 09 8F
 4F 40 66 31 B4 EE DD EB 56 EE 82 82 61 84 6D 0A
 C0 D7 30 EF 46 C5 02 64 68 C6 4A B8 CE 4B 87 7F
 F5 3A 0B 42 17 E0 87 F3 E3 61 16 29 29 A2 42 3D
 79 0F 70 EE 66 2D 22 3C 4A F1 CE 5A EA 1C 83 44
 A3 E6 98 18 84 C3 93 1D 2C FA 30 35 6D 78 CA 69
 1A 3F 4F 9E B8 3D D3 28 FC D6 88 57 D0 B5 12 94
 47 18 80 7F 06 9F 0B 5C 3F B4 EC EB FE 2A AD 42
 C1 C0 3F 6C F8 CA 67 65 20 1D F5 CF 51 BB CF 55
 C3 73 4B A3 DF EE C4 DB 57 EC 22 86 0A B4 C0 2A
 37 F4 48 2E 9D 21 FC 31 CF 22 B7 06 3D 3A 70 15
 D3 B1 1C CA C7 82 85 43 EC DF D1 A2 14 BB A0 67
 70 CB 75 2D 20 EA 54 0D EF A5 71 9B AF F7 32 60
 4B A2 6F 7A FC D1 F2 CD DB 50 02 5F C9 50 28 8F
 93 FE 96 FD 54 B7 89 9F C9 E8 25 AA AA 58 D7 9D
 16 E5 A5 BE A1 90 28 B7 EE 7C CD 69 1D 3D C4 82
 52 4C 54 54 E6 DC D6 AD DB 43 42 87 7F AE 4C E6
 9E 0A EB 30 8F 56 88 F0 56 59 B1 FA 73 1B CB 7D
 9B 72 18 25 C6 EA 5C 85 89 76 B3 FD 42 EF 33 6D
 A2 06 0D 2D 51 BC F1 34 DC B5 8B C1 04 9B A1 F2
 6D 2F 2E FD 6D 87 B4 D8 31 01 D8 7B 72 AF 77 49
 58 38 54 B1 A6 7E B5 5B 62 94 1C 15 86 3D BA 5B
 3B 3F 50 6C 21 5D 7B 95 9F CA 08 3C 95 0F FB 40
 56 99 97 EB B3 A2 E2 3C 22 41 49 B0 A4 09 76 65
 AB 96 D8 3D 83 95 4A B0 98 F5 AC 82 69 89 3A 78
 5F 01 8F 48 1A 50 30 69 6A 90 A1 1C 41 12 07 76
 AD 0C 3D 3E A7 B5 90 DD D8 F0 A7 EC 14 FC 21 72
 57 05 58 6A C1 63 05 18 A2 87 3D 1B E6 98 D8 B8
 30 B8 F1 F3 BB 1B D4 22 0F F5 41 18 9E 27 24 18
 FA DA 03 E5 52 9D A9 58 95 68 3C E8 24 E1 83 63
 B8 91 02 33 4E 93 B0 32 C6 7B 35 59 D0 8D F4 58
 D0 5F 01 8F CF 7A 10 96 3B FC A1 1A 6E B9 78 79
 D3 FB CE A0 1C 5C B3 64 A3 1E A4 71 53 8E 01 0E
 4F 84 0F F4 0E 21 62 6B DC 3A BA 75 85 80 E6 DC
 35 E9 85 CD 15 8A 3E 8C 25 9F 7A BC 23 FB 37 2C
 D1 F5 4E 38 7D 58 A4 FF 16 E0 82 E7 62 A4 76 AE
 CF 99 E5 07 1F 5F 9C AD 10 CC EC 0E 12 C8 2B A9
 D9 3B 59 92 59 55 B3 92 79 BB 47 02 41 6A CA B1
 EA 26 3A B6 E5 6D FC 09 52 8F 4C 0F 16 3C 14 47
 CF 1F D3 B9 12 74 81 2D 60 86 96 AD 86 BD 6A C4
 C7 8E 23 9C D8 03 08 29 21 BA 74 0C 5E EA 68 6E
 2A 04 BE AF 0E EA FB F5 F2 A4 5E 40 F2 70 51 2D
 2E A8 F2 1C EF 44 CF EF A2 4C F1 5F 3E F0 FC 61
 E5 BD F3 6C 19 E7 9A 6E E9 5A 6C EE DE 65 72 9B
 58 9D 80 A1 6D FA 8A 1A 0B AE 30 62 EA 04 0F C4
 02 57 D5 0D 08 A0 95 E2 1D 46 0D 1E 33 58 06 19
 43 69 56 6F B7 B0 13 36 71 44 B6 B5 6C EC 39 B8
 28 A1 FC 2E 59 5B E1 A3 86 68 B8 6F 7D 24 A6 8B
 DE 5D 5E 2F 32 89 25 D4 B1 98 D7 32 EB 4E 82 C1
 DF 53 F7 41 17 ED F2 7D 29 8D D9 07 17 A3 3A B9
 09 6C 01 70 19 3A A6 53 FD CD E1 D6 CC C4 FC 05
 7C E5 D4 B2 7D BA 52 D7 B8 AC F4 82 0F 78 17 1B
 FE B5 4A 32 1E 01 E6 73 3C 1B B2 E2 11 B1 EA B1
 10 2F B9 16 C5 B4 6B 4A E3 06 38 53 47 09 A8 C7
 94 FA 9A 47 AA 9E 32 1F DF 88 FE 2D DE 69 69 5E
 6A 99 97 D0 E6 E2 56 A9 F2 3A D1 6D 98 91 30 E5
 DF 1F 9A 30 61 4D 34 74 C6 76 61 D7 6F FB 92 CA
 16 52 C7 37 BA AC CC B5 AA E7 F4 4E 5D 0C 89 CC
 AD 85 E2 D5 DA 6C 89 8B 4A 3E 9D 3C 1B 84 F3 20
 FC A9 DD 92 63 04 4D 25 13 6B 8B 88 3D 03 32 F6
 BF 0B 04 42 43 7F 4E 6A 4F 9E 68 13 57 DA 76 F5
 F7 AD 5B 29 C4 B4 B2 35 97 6F 16 14 74 9A A1 7E
 88 53 13 DE 9F E0 98 FE C6 A4 96 2F F6 0E 11 14
 DE C0 CE 0F 02 7C 41 54 C1 A4 EB E1 9D 54 33 35
 50 44 6D CA 1E A0 3A 44 F3 59 35 C8 7A 8E 87 2C
 D7 8E 6B 66 C8 0F 7D 87 01 67 43 05 94 0A 6B 78
 2D C4 0B E5 B1 67 FE 16 C2 BE 54 37 0C 1F 18 D7
 A3 F1 EA 8B 90 DA 05 43 59 97 AD 56 2E E7 ED 38
 C9 FB AD B7 53 0F 0C BC BD C1 23 E5 20 74 E5 2B
 E4 3D FE 98 17 2A 63 9E 8E 73 F6 0D F3 26 E1 B6
 A2 B8 5E 6F 17 B2 FD 47 E4 84 36 3A C0 D3 F0 02
 69 F5 37 52 B8 C9 29 E6 BC 8C 66 59 51 08 75 55
 FF AF BD 44 C7 78 14 F1 0E B1 B0 A5 81 91 B5 E1
 7D 12 EA 36 CB 93 CC CE 1E E4 51 0E 48 D3 93 F9
 53 84 FC E2 B9 83 DC 10 DC 58 8C D5 87 7F 01 5B
 FE 3D 24 FB 49 68 1B 0E B6 DD F1 02 33 C1 96 DA
 09 D8 6A 19 A2 A4 9B 3E 93 F8 FD F0 03 5D F2 B8
 FE B0 54 4C 9A 0B 51 4F A2 C3 F6 56 67 1A 9A A4
 A0 F3 97 7F 38 78 30 92 98 41 F3 78 B9 98 FF 63
 4B A7 22 C7 0E 03 28 A2 9D 78 BC 64 68 52 27 1E
 3C 21 41 BA 8E A3 A4 F7 F9 49 9A 92 33 91 DF 5F
 29 2D 4E 33 DA A0 BD 8E 27 EA 2A 74 46 8E 7D CE
 9F 94 E9 53 7C 4F 3F 84 40 B1 D0 64 4B 0C B6 73
 C9 85 82 A5 47 B3 BD 82 C0 20 43 2A 2E 5A 64 EC
 9E 14 99 97 18 5B 67 DA 3E 93 51 9E 30 0C 06 3F
 AB 63 01 87 1F 42 27 20 8E A1 88 CD 53 D5 0F D9
 3A BF F9 E9 A7 30 35 6E 55 0B 57 F4 52 85 E3 45
 A6 59 B0 E2 72 A4 CC A2 D0 84 1F 08 CF 58 74 34
 09 DC E7 1C 48 1C 77 C4 3B EB F5 FA C5 8E 02 77
 C6 E1 31 AA 1F D9 6F 7A F8 3A B0 73 37 36 17 2B
 D6 EE 24 0B BB C0 0E F6 2F 11 7F 17 94 B7 D1 3B
 D4 67 4A D1 AB 96 6F 7D 3B 0A FE 05 7A 6F 5C DA
 D1 86 45 F9 72 99 75 67 A7 59 1B BD E9 5E 25 68
 1A C9 64 40 E9 8E 2F 85 11 7B F7 82 3E 87 35 B4
 57 3F 1F 9F 49 20 23 63 F7 25 96 71 AB BE 50 5E
 15 BB B2 6D 38 1C 5C 8E 80 85 01 B6 16 B1 5A CA
 AA FD C7 36 6F E6 78 12 FE 35 52 4B 96 16 4F C4
 20 C4 BE A4 D5 D6 D0 84 3E C2 17 7B BC B6 40 F6
 3F D8 9F 37 C4 3E 33 D5 29 B3 CA 55 A8 35 26 76
 9D 99 A9 C4 A1 6C 74 E4 59 E1 AB BF FE 9A AB 89
 FC F9 FF 62 4C 15 92 4D C5 28 1A D6 7E BC 60 E3
 AA 62 1C FD EE 99 6B 02 49 1C D6 C4 74 19 62 61
 0F 60 A3 10 EC EE 56 7D 66 2A 61 76 FF 1E 92 BA
 D0 35 C7 F4 F1 C8 58 77 09 78 1D 2C AC CC 30 67
 EC 9C 98 3F 40 0B 16 1F B7 07 4D 7D D1 D3 29 D1
 48 00 9C 66 71 B9 E1 2F 4F DD DB CE 90 56 7C 7D
 CC 23 9C 27 48 04 10 F6 7C DE EC 26 79 CA 0F E4
 59 B2 EF 09 54 2E 30 F4 B6 A6 0D 6E 31 FC B7 08
 2B 76 00 D0 49 E3 8D 8B 06 A2 B8 48 FF 77 F3 E2
 8D 6D 1D 99 93 8C FF CA F4 7C FD B0 0A A1 08 A3
 51 BF 5B 4A 08 5F 34 24 67 4B 90 D4 EE 3B 07 97
 C6 D5 92 8B 2C A8 BC 5E 4B 6D 22 12 D5 A4 53 3F
 58 66 91 39 34 4E AF FF 17 C7 6A AC 24 7E 0D 4B
 9C 86 F1 AE 1D 6A 95 5D 81 99 F5 A6 DA EA 66 40
 C3 B3 D3 6E CC 25 6F 39 9C 2C B0 35 0E 2F 40 F3
 A5 B8 C3 D0 7D AE 39 31 06 20 DD 04 AC 02 14 B4
 07 10 BC 92 13 56 9B 5A 7A F1 44 19 46 17 EE 1D
 B4 9E 3D 00 08 FB 74 D8 AC 60 61 77 B3 7C 29 8B
 C7 E2 2A 37 5D 47 69 75 5E 14 78 CA B5 A6 D8 8A
 52 94 10 C4 BB 6A 36 EA 38 D9 DF 3C BA 20 09 C2
 9D 10 4D 50 53 93 DC 67 3D 7C 45 18 B6 BB 66 E1
 39 B9 9C 05 A4 A0 FD 05 63 54 EE EF 95 34 D7 CB
 61 B2 E5 90 66 37 28 0A 9A 75 CF EF 5B 5D B2 AB
 91 12 FB 57 48 85 ED 34 08 76 98 6A C4 BC 04 7F
 95 F6 9D 2C CE D4 4B 56 24 63 92 0B 7D 47 92 B4
 1F 40 1A B9 4D 03 CE CB 96 09 EF F5 A6 A9 E4 23
 6D 57 6C E1 35 CF 5B E8 65 06 92 ED 33 83 CD 47
 73 C1 E0 43 31 8C DF B0 4B A6 B9 8A F3 29 20 BE
 A6 29 5C 28 DE 6A 3E 26 71 FE 31 D0 18 B7 DE 7E
 38 55 01 3F 7F FC F6 B7 64 D6 0F DC DE 31 35 C5
 7D 52 6A D2 21 E6 6B AC 4F 0D 53 EE B4 43 53 BF
 45 E1 45 4F 61 50 DE B6 1E 98 C5 F6 A9 0F 84 F5
 ED 30 34 C8 48 F5 5C 78 4A 2E 84 AF 2D D1 98 D7
 9B 10 62 E6 F8 6C 54 72 29 1E F3 D6 95 1A 8A BE
 EC F6 80 4C 20 C6 8C E1 5A 56 CF 07 97 25 29 57
 B8 20 22 00 A9 24 81 C4 E3 8D 42 BB 43 31 ED D9
 9C 86 F2 F7 05 BC 3B 9B 88 1E C4 E9 3D AD 38 EA
 33 F2 4C 79 18 E0 20 96 A4 DC B4 D2 37 DA 96 D4
 19 15 17 58 8C 5A 9E 8A 5B 4B F9 33 A2 DA 00 91
 42 F6 26 1C B3 A4 8B B9 20 E9 DF 69 D2 96 21 C6
 79 34 BC C4 28 3C E5 AC 91 CC 0E DE 20 2D 6D A9
 96 9D 69 D8 60 E7 0B 87 B1 AA 5A 29 78 0D 51 F0
 F9 2C 9D AE 91 A5 DE C2 EC 4E B6 43 29 80 65 D5
 2B 7B 5C 70 87 94 62 C8 23 D5 FC 08 5B DA E3 D7
 27 FD 60 A7 22 D0 B1 09 65 19 AC 8F 04 AF B0 28
 5A DB AA 46 9E 82 BA 7A 74 84 42 F8 AF 97 BC 08
 00 19 FE A0 96 AD 8C F5 DD D3 1F FF 08 3C 2B 4F
 F4 F2 55 01 96 5D D7 C0 57 39 FB 72 2E DC 9D 29
 F2 E0 9C D6 80 83 98 A4 BF AB AE 26 CE 62 5E 60
 C0 4E BA E2 6C F3 A2 78 36 01 30 F9 30 A0 CB 8D
 CA 3E 1E 5F 8A 3F 50 77 68 FE D7 CC 23 40 37 17
 1B 6E 3A FB 74 03 4E BF 50 33 D7 8A 5B FA B8 35
 83 6F 0A 1D 4D BD B0 3C 2F 22 83 77 B2 B2 8F 8F
 6A 8C 24 D9 97 62 B6 42 E5 5C 5E 3F 04 14 21 4C
 6B 8A E7 5B 40 ED 06 4B BB E3 2F 88 42 EC 57 9F
 C9 77 CE A9 F4 87 C5 96 A8 F9 F7 CB 0C E4 43 D4
 BC 11 E7 55 1F BA 4D 8D 81 ED 5E C5 5E 79 B9 15
 1D 42 A1 1F D0 40 16 49 06 F7 79 3C EF 37 0C 06
 50 9E BE 7A F0 17 DB 8A E5 86 F6 48 88 90 36 7D
 8B 8C 68 FF CF 78 1C 9A CF 24 58 F6 FF 25 BD AB
 81 88 90 5B 3C 35 91 48 9E 49 9D 23 A5 DC F9 DA
 5F 4F 5A 60 B6 5D AD CE CF 63 B4 3E 9B EA 4D 96
 71 8B 5B 10 40 83 7B 74 23 5A E9 2B EB E7 13 45
 FE 7B 60 9B 5D E3 7B 36 6A 19 84 50 37 E0 68 BF
 85 DA AF 95 CA 9B 98 10 EA A5 F1 66 CE 95 0E E2
 56 36 5E 1A 87 3E 28 B7 5E 1A AB 8A B8 2D E4 C3
 F2 F8 31 91 1B EB 7A 8E B0 1D 06 68 01 53 03 13
 E0 FC 84 97 B8 F5 87 75 A3 89 7F DB F1 4C 35 AF
 D7 9E A0 CD 9D 86 EF CD 1C 32 A3 3E D4 C4 E4 EC
 22 7C B9 A6 99 78 BA 82 E9 E5 F6 45 FE 4C DB D1
 A6 08 04 10 A4 24 2D 8F D9 80 61 D8 60 CF E4 1F
 01 E4 89 56 02 8D 18 4A 30 B6 C1 19 85 03 E7 EA
 89 7C 09 03 79 C4 8D 93 63 6E 2A A9 AF 95 73 B1
 51 B6 22 49 C0 B3 D2 DD A5 7F 3B 34 7E 4C 52 81
 E8 09 85 EA 1B 59 32 6F 59 15 93 DC EC 82 6C 02
 E2 B6 2C A8 BD FB A6 83 94 79 F3 3D B7 98 57 63
 44 ED 65 00 66 8A FC AB CA 31 7F 22 AB F9 84 9E
 7C D8 AF 79 D0 69 B0 80 0B CD 30 96 68 60 20 6D
 3F 5C 91 5A 78 69 5D F3 3D C9 AA 3A 07 67 BD 66
 CB AE FA 2E 10 2F 56 CD 11 5E 4C B9 37 33 EE 76
 B3 28 81 A6 F3 38 5A 19 A8 C3 CA 7A 64 3C E0 AB
 CF F7 56 91 AD B0 44 E8 4B B1 7E 14 1E F5 4F BF
 CE 2F 1F A6 B1 A6 B2 D0 CD 5A 59 6B E7 89 DC 0C
 26 08 C9 65 43 8C F1 62 1A D5 08 14 0E B4 62 FB
 41 83 89 D7 8C AA 23 7F 41 47 7D 88 F7 25 9E 8E
 7D 63 A8 3F 45 78 29 7E 73 7F 4C 78 DA 34 0E 60
 70 83 3A A7 5F 46 B3 1C 0D E5 10 9C DF 0D BD E5
 94 63 7C AA C7 00 59 42 69 F0 71 2F 84 0D 70 8B
 3C E1 7E 87 42 44 08 4E EB F0 D4 34 D9 F2 E7 49
 0E AE 8B 94 CC CA 6E FC 1A 59 C3 E0 EF 97 B9 3D
 97 B7 37 A4 EF CF 4D DF D5 58 EC 26 40 FC 26 E5
 FE 7E A8 55 0A D9 A0 CA EA 42 89 3E 98 ED 52 1E
 A7 77 C8 11 85 23 2A BA D0 27 FE 75 1A 81 BF 24
 E2 4F AA DD AA 28 DB F2 F8 6F A1 83 47 23 4C 36
 6B 01 8C E3 12 3D D5 65 7F 71 5B 77 E0 5C 27 F4
 14 96 D3 71 43 A8 C6 2E 31 22 70 10 E2 A9 37 8C
 09 43 2A 2B 9A 11 51 FE 84 7B B9 53 5A 53 62 C3
 9A 3C 61 90 8B 4B C2 B0 7B 2A 9E 97 C2 85 13 16
 41 EE 4E 2B 9D 30 B4 85 94 22 D2 38 7E A7 67 E4
 D4 15 68 19 61 47 D1 7A B9 43 3C 66 7D 34 4B 48
 81 FD 34 C0 88 6B CB 9F EF CE 2E 0F 11 17 EC 6C
 13 CE AB 3E 62 84 30 69 A7 B5 C6 66 F8 2B 3B A3
 B0 60 1F F3 F8 AB 52 9F 52 EF 43 8F 0E B3 18 E0
 3E 62 8A 48 20 B3 31 1F 54 55 FA EA 10 CE DB 91
 1B DB 15 2B 61 4B 65 B5 B4 3A 4D EF 8F 81 69 0F
 8C 6B C5 EC 5F E3 8C A3 FE D6 A4 B5 42 0A 77 1D
 CE 5D 76 35 CA E2 92 18 52 3A C1 8B 26 CC 59 3B
 2F BC E4 3D 58 0D 24 BF FE 78 67 C2 9C 5E 00 33
 C3 E5 A5 53 0D 64 A7 35 8D 24 26 3A 2A 7E 03 47
 54 70 BC 60 44 4A 7A 1E CB 7A CA F7 21 A8 52 41
 03 C5 76 A6 E2 9F 07 1F 1D F3 AD 87 5B D2 F3 DA
 CC F4 2B D0 7B 32 07 70 70 C1 A6 E6 FC FA 33 BB
 B8 FB C6 30 F6 76 C6 77 6C 00 41 F4 B5 3F 72 B1
 66 44 CF 68 D2 B0 5B A2 3C 74 5C 8F 2E 62 A1 79
 5C CF 02 85 96 7F 45 31 BA D3 8E B7 19 FA 3E A8
 C7 0B C7 4D B1 AE 54 6D 35 1A 3C FA B5 5C 73 C2
 F4 E2 F5 7D 80 A3 CA 85 68 2B EE 00 A9 A6 08 86
 97 6C 29 85 0B 4E 12 5B 56 1A 1E 0B A4 D6 01 71
 5D 8D 60 F3 43 4A 93 72 16 85 D4 A0 50 9F B1 E2
 C4 56 0D 35 46 3C B5 38 6C 13 CB 97 86 DD 87 EF
 3C E6 82 15 FC 6D 40 AA C5 31 2B 2A 87 1F 6D 73
 D6 89 45 94 13 55 E4 6C AE 8E 25 64 FA 2C 85 3B
 EB 63 E7 4B 71 D9 8B 6A AE DC 5B B7 AB AA C6 12
 8D 73 37 DA A2 D1 13 A6 9E D7 20 10 13 40 C2 F4
 A6 FE F3 C3 AE 6E 18 36 01 5A 0C 1F BA C4 32 D5
 23 DE 06 86 A3 82 7E 4B 59 CC 93 C7 24 91 C6 B7
 CA 2B DC 3D 98 CE 18 8C 28 07 62 34 21 1C D0 9E
 EF 92 3E E0 6E 53 B4 E8 7F F0 8A 77 F9 AE F0 AB
 C2 2E 0D E9 B3 77 FB E4 56 99 C4 34 91 BB B9 2A
 F5 C3 75 61 EA 51 5B 29 9D E2 DC 0F F9 49 9D 44
 DA 1B 5B 48 0A 32 4D CB 99 22 EC 52 69 13 DB 0E
 0B CC E5 DA EB 8A E5 4D 3B 9A 66 99 A6 45 DB 18
 15 CC 83 E4 8B C7 DD E6 27 D7 A1 0E 7E 05 80 83
 F4 02 51 97 8D 27 EC 0A FE ED B1 C3 06 26 04 FE
 F4 A8 51 82 A6 55 4A 24 3F FC 00 70 16 6F BD 2A
 B1 D2 51 13 6C 0F 1D DF AA 97 5F 3B 10 D2 E5 24
 DC 0F 4D 3E E3 A7 EA 10 C2 69 E9 61 1B BF DD D7
 B1 1E D8 CD 50 D6 65 D1 03 A3 26 65 81 49 0B 25
 5A E3 EC C0 32 2C 6B 62 99 C7 08 BB 07 BE 7B 33
 26 E8 D9 F4 F4 3F A7 33 5C D3 05 96 22 AE 8E E4
 89 64 F6 4C B2 C5 E5 BE 80 D5 01 22 75 31 9D 1D
 1F 41 2C C7 34 86 62 6F 53 C7 60 78 71 F3 BB 46
 D5 6B 6A 38 E4 0F 84 F0 A2 79 B3 59 7D 93 76 98
 D8 B3 A4 38 F2 BB BA E5 74 08 F6 1E E2 68 5A 7F
 0D C0 1C AC 69 A1 28 CC 09 8B BC F9 0E 4C 44 CC
 22 2D 6C FC 14 DD AD 83 2E 20 C3 8B 48 7B E8 BD
 F5 5A A0 21 90 A0 26 C8 11 68 25 F6 A2 19 A5 DC
 26 E9 99 88 09 91 A1 0D 07 73 EA EB F7 3F 30 FD
 8F AE 97 C5 5A 1C 83 75 92 CB 67 8F 24 10 62 DC
 87 8E 11 87 07 A2 8E D0 17 FB 83 B2 29 66 15 72
 EE 03 84 FE 53 74 C6 B2 AD E2 23 E1 72 A3 1B 00
 7A E2 24 BE 5F 70 47 D3 1C A6 74 45 23 DA 82 34
 25 61 CF DC 49 19 EE 5F EA 5C E9 0A 2B 4A C7 75
 FE E1 42 9A 11 AC 57 99 0A 80 EE 01 34 BA 32 2B
 45 69 93 90 77 14 43 45 BB 48 64 43 A9 8C 07 96
 DF 0B 1D E6 AD 77 FB CF BC 63 4D 4E AB 51 C6 7E
 05 FC C7 DA B7 44 CC 2F B5 12 13 81 FE A9 3D 8C
 3A 1E 10 76 78 72 13 BD D7 B1 0C F4 EE B8 EC 51
 BD 46 9B 44 5A 96 1A 6F 3E 02 07 64 11 C2 78 58
 29 28 24 3F 90 BA 0D 49 6F 53 79 09 60 52 BC 34
 36 24 8A 66 62 DD 44 07 81 B9 38 CB 26 6A 1A 4A
 FB 63 7A 45 C5 46 93 F1 F2 F0 6F EB 34 4C A3 FF
 FF FA FD 30 AF B7 AF 05 BA 24 F1 95 CE 1B 42 49
 5A 24 3A 5C FA 66 33 03 D0 75 ED DB 9C 1A E3 5F
 55 88 C6 BC 86 24 E2 79 F0 5C BE 83 9A EE C0 C3
 30 DB DC 6C 60 5B 72 AD 2A A4 22 B6 F0 F0 F1 F3
 1C 12 EB 39 6F 15 7F D9 32 7D CA F1 45 E0 06 40
 91 BF F8 3E 5C 87 6C 3D B5 2C F8 2D CA 84 94 6F
 C7 0E 74 23 0B A5 AD 47 FA 6E 8E C7 88 2F 33 E5
 C6 AB 88 DE 70 45 F2 A9 39 F1 B8 A4 05 54 54 E7
 C4 0B 47 2E FA E3 2E A2 53 34 22 3D 0A 52 6B ED
 4B 86 62 B2 8B B8 76 58 3A 91 6E 55 E4 D5 8B CD
 1F 0F 2D B3 13 93 CB F7 4E 18 9D FE 56 03 DD 10
 15 62 CC 90 7D 57 74 B4 DC D2 0D AF 8C CC 59 A2
 27 A5 BF A1 5B 27 59 71 2A 56 37 8C EB EF DB 0B
 1B 76 61 E2 F2 1D 4D C7 FB BE ED AB D1 AA 8E C3
 45 90 15 8A 3E B8 FA B2 08 CF 94 82 DB 14 3A B2
 78 93 38 7B 51 65 46 B8 3C 4B DE A8 1D 0A BA 14
 93 E0 97 19 AE F4 FB B2 25 9A CE 34 C1 C0 0C 2B
 6D 62 ED 59 C7 4E 81 52 F0 4D BB C2 3F 1C 01 3D
 74 A2 96 0E 3A EB F4 C0 C7 FD 80 1B B7 98 35 E5
 AC C7 B8 60 2A 91 2A 2C 72 8C 5F A4 A0 AD AE 45
 B3 82 22 D7 C6 4C 8B 51 40 02 FC 5B 59 6F F1 D1
 01 C9 1C 80 44 4A 29 41 4E 1B F9 D3 AE D1 A5 CB
 22 C1 CC D7 CA 7F 91 56 D0 14 85 DE A8 4E 1B 9A
 EB 70 2C CD DC 62 A5 06 58 2C 6E 93 59 CB B2 6F
 A2 E5 A4 94 22 87 D7 51 AC 41 1B A1 C9 61 9B 7E
 3D 41 9C 3E 7D 06 9E 18 37 FD D5 F3 21 3C 2A 37
 2B E1 17 E8 80 00 E5 2C D3 C7 36 27 7B A0 45 9C
 3C 16 6F 7D 8B D1 C3 CC 75 7B 74 4D D5 69 E4 B4
 50 DE D7 F4 69 19 1D DE 4E 73 AD 60 BC 59 5E FF
 46 C9 5D 45 24 F5 F8 37 F1 E8 12 DF DC DB 7B 4F
 BA EA F2 EA FE E2 B3 D6 2D AC 97 D6 D9 DB B7 6C
 8E 2C 1B FF DD B0 C3 17 39 83 B6 80 A9 79 C3 DA
 7E D3 5E 06 78 C8 03 23 F9 35 51 59 C5 2E F7 34
 C0 63 9B B2 19 B4 DA F4 27 F8 7C 97 2D 7D 06 70
 9B 2E 45 75 4F 59 AB 65 82 73 FA FE C0 21 A8 90
 85 C1 9F 83 A8 2A 72 29 50 99 A4 61 6F B6 29 5B
 77 A3 CE 6E 90 24 60 C7 76 CF E8 0F CB 18 BE 13
 62 DC 70 28 6A 3F 42 E2 45 4D C7 D8 C7 8F D0 D7
 CA FC 48 01 BD 1C 35 F7 99 28 23 D4 B3 12 C1 82
 8E 94 84 18 4B 35 F1 36 F4 00 55 47 A1 4A 9D 1D
 20 92 09 BF 1B F6 3A 50 03 67 C5 BA 2C ED 03 68
 91 8F 82 66 C1 F5 E6 DF 3E 3D 75 CE E4 A4 F1 F5
 26 3D 3B AE ED F5 AF 2D 0C 99 39 82 E3 4C C1 C8
 87 BC 18 84 22 13 D8 A5 65 B4 DE 92 67 45 31 08
 38 31 89 FB CE 21 78 60 1C 83 9E B7 84 5B A6 5C
 02 98 41 7C 5E 40 7B 9F 45 42 EA AF 4A C7 17 D4
 D5 7C DD 4C B8 BB CD B5 1A 6A E2 49 E7 9E 6F 2A
 62 F4 20 96 0E C4 37 64 B5 C7 DB D6 0A 24 79 BE
 7F A6 5C 1A D1 4E 2D C9 4D CA A6 B7 5D DC E7 00
 47 FB FE 4D F9 24 C4 09 D4 A0 A6 6F 47 9D B7 90
 3A 59 61 60 4E 61 06 DA 45 29 06 76 1E 1C 49 3E
 83 A8 1C 0E 65 3D 8E 89 3C 7E 51 1B 93 7D B5 D0
 F8 6B 50 B8 87 58 70 2A BD 68 DB 9F B1 42 47 EE
 48 EE C3 37 DC 32 73 19 34 FD 28 9B EF 68 EE 4A
 57 DE 78 64 22 C6 8F 76 60 F5 32 E6 07 7C 81 A1
 1C 1F 3D B2 A7 AB 1B 32 4B 39 CA E2 1A C3 33 B6
 A7 B0 BE 50 84 62 62 49 A5 E6 0A 26 1E 26 9C 0F
 3C 63 B3 46 FA C4 A6 AE 85 70 01 9D 81 01 5A 90
 44 76 DC 8D E3 66 29 71 2C 73 6F 57 13 17 A9 10
 E3 FA 89 A2 3C BA 1F 99 ED 86 AC EE 27 7D AF 81
 4D 35 74 21 34 A0 5C CB F8 1C 95 3A D8 65 46 D0
 B6 F9 E8 9C 78 B8 AA 99 CB 9C C3 09 35 AD 59 FB
 19 07 6F 45 FA 92 92 5A 6B 39 B1 D3 E9 5A 87 71
 F5 34 F5 DE BB 5F D9 AA FD 08 F9 B2 02 3B 00 99
 A0 0F 6B 85 60 D8 10 EC 25 30 25 E6 9B BA 75 1E
 68 14 D8 89 F4 65 90 CD 10 D0 CF 68 AD 55 56 69
 B4 3A 84 35 8C 99 7D F1 BB FB 0E 50 C5 7E 1F 75
 65 15 B2 7C 88 08 D7 7C 1F 94 FA 2A 5F 57 6F F3
 A6 D2 11 90 AE A0 37 46 89 25 13 BB DE 61 1E D5
 77 44 FA FB 41 AA E2 5D 6D 17 2E 8D D0 E7 6E 79
 05 C6 0F 89 D3 90 0C A7 1C 52 BC C0 3C DD 0D 13
 FE 81 33 40 BE C0 0A 43 BE 7C 9D FD E3 4F 86 11
 D1 92 A2 2F 4B 71 29 FB FA 8A 95 4F DF 3B F0 6E
 0A 2A 8B 8B 02 F2 87 1A 8A B3 DC B3 69 43 9E 9A
 A8 9A 68 28 04 FF 09 36 B0 32 5D 08 DC AA 33 91
 D3 DD 3A 32 A9 32 C5 EB 1D 2A E3 5C 3E 5B B1 75
 6A 5B 91 8B F3 F8 EA C2 89 72 E3 92 0A 14 0B 92
 3A 3E 80 FF 3D 1F 9E 6B 51 D8 DC 42 A0 E8 37 C6
 09 4F 5F DB AF 6B 72 9E 2E 6A C7 17 DA 8A BF 56
 85 FC D7 8E E3 B9 D6 2A 90 53 70 12 CE CC AB EE
 FE 98 EA 2F 8F 80 8F 74 7C 4F 55 D3 97 F1 B0 20
 11 65 13 00 E2 81 69 2E BB 9F 16 8B EE B7 AE A6
 9E 2B A5 2E B9 7D D3 35 3B 11 CD A8 A8 B7 8D 72
 BC DE AA C3 79 98 57 49 38 1D 8B A6 86 0D EA 33
 DE F2 D8 D2 79 7C B9 34 E5 C2 06 87 49 CF C7 AE
 6E DA 73 FB 27 9C 73 A9 8F E9 78 82 75 BF 57 58
 1B 92 ED 2E 2E EE 03 60 0E C9 FC ED 76 68 9D 94
 2F 39 25 71 5F 7D 47 E6 E8 E7 8B F9 69 31 82 87
 72 64 B7 68 24 72 91 E7 18 C2 7F B9 8C B5 BD 44
 D1 32 0E A2 FF 54 3A BB F4 EE ED 4F E6 BB D7 E6
 84 5C 8C C7 D6 54 57 3D 1B 58 45 E5 04 43 1B 66
 B6 C3 EE E1 63 3B EC 07 E2 4C BA 98 F4 33 CC 6E
 DF 57 87 29 12 40 63 5F DE 5C 40 72 24 73 C8 0F
 12 C9 2B E9 2A A0 BA 5E FB AF ED 69 3F 2D 21 FC
 08 82 2C E7 6A 78 2C 33 3F B9 9C A0 7A 32 97 01
 26 78 74 6D 3D BF 6D 30 AF 20 55 44 27 25 49 2E
 E4 C3 09 2C 1A 3F 49 CE CD 7A 88 F9 B4 DF 07 88
 51 AF 13 E6 0C E5 E5 8C 10 26 AA 89 B0 E8 B5 B4
 5C A3 19 42 55 55 A9 B1 64 34 04 CE D1 8B 3F 8D
 B4 0C 88 13 9F B8 DE 21 14 FC 24 07 9D 78 39 A1
 74 E6 0D 89 D3 32 C9 FB FE 1D 5C D1 27 90 3C 7D
 53 0C 33 65 5B B9 FA 5F 8E D1 83 3F 27 43 08 53
 B5 2C A0 5F EC 82 1E 25 C5 98 4F 44 60 30 89 F7
 ED 0C 5C 50 F5 0E 28 A5 E4 3E 2C 1D 03 66 60 A9
 62 15 2A F0 E7 9F 28 BF 4B FA DF FB A2 3E 30 01
 61 57 D7 AD F1 36 FA 22 D8 9A 03 28 5C E9 01 B9
 E7 D7 1F 49 A1 CE 2C 69 BA 38 04 8D 0C D4 33 8F
 48 A5 98 40 6A C3 50 CA C8 B4 48 33 30 25 01 D7
 28 86 20 79 0C 3E 51 8C 7C 42 FB B6 A8 E3 B3 7D
 AD 20 6C E8 A3 12 57 09 0D 64 AB 35 7A 17 07 A2
 04 42 50 75 83 D6 77 98 C2 02 45 FA D0 22 3F 3C
 32 18 DA 9F 2B B0 3F 80 57 9D 14 8E 2A 67 13 3E
 3F 8E E4 40 85 A7 28 6E B4 AD 58 82 F2 98 81 A0
 7D D8 4F 93 90 BE B7 5C 2A 65 CB 69 BB 85 BC 1E
 C9 98 DC 60 06 06 6A 5B 47 02 49 45 1A FD 63 0C
 F4 90 01 59 56 95 DA 39 FF 17 16 C2 6B 46 FC 37
 8E 18 5F CC D8 EF 2C 78 F5 4E 2D 20 4F 8A 7B B9
 F2 98 F2 55 11 70 57 85 2C 8B 8E D5 8E 65 C4 E3
 BD 22 7D DA 50 A6 95 5A EA 3E D0 B3 D8 79 4A F7
 D0 60 FF 6F 8C EF 7D EF 62 E6 7C E8 BB 04 57 DB
 F9 AA 9C 0E 11 31 89 22 BC 2E AF ED CF C6 C0 28
 A2 94 26 6F A5 15 B8 87 0A F8 91 0D 0D 90 89 AB
 B7 44 0C 82 F1 B5 B5 CE 7C BE 0B AB 9B 3E 39 CD
 16 54 A6 54 24 4E 55 41 0C 80 6D 6D 33 99 FF 93
 CD 46 EE 94 37 23 8B F6 F9 E1 E5 C4 F9 EC 46 13
 42 98 3A E2 28 BA 6B BD F1 0B E2 36 BE BA 18 B6
 A6 30 38 97 E8 88 D7 CB 22 9D 9A 58 E7 9D 1A 74
 46 3D CE F3 39 27 15 FB 53 D7 D2 93 22 39 3A A7
 13 F6 80 A6 AA BC BD A7 52 50 E0 56 62 22 63 91
 C6 37 AC 39 8C 31 04 C8 79 38 09 95 CE 63 B1 21
 F5 5D AC 95 A1 C3 30 39 14 58 61 7E 9C 0F BD EE
 76 A3 88 0C B8 91 84 BF 9A A9 59 4A E3 80 02 95
 3D 5E C8 4E 0B 14 38 69 9E 23 DE 22 6B 89 32 2E
 3E 73 FB 7D 67 15 87 C5 52 CC 0E 22 A6 2E C6 D0
 E9 9A 27 5F 5F 49 AE E2 A2 13 5B 5A 8D A4 A7 7C
 0C 0E 8B A7 16 EE D3 00 76 E0 95 67 F8 37 FD 1F
 0B 1D 95 98 EE 1C FF 6A 54 7F BF 8D 3A 77 1D 8F
 D5 10 97 D8 5C D7 54 BA FE A9 1D 11 AE 50 3C C0
 62 44 F9 4B 44 FD FA 7C A2 E6 24 6B 0D 75 DC 76
 A2 30 71 BF 14 1C 9E 4D 49 26 9D B8 77 4E 72 A7
 14 2F 9C 83 D3 61 DE 9A 98 07 D6 03 CE 0A F3 A5
 AE 36 01 6E 2D 4C 8E 4D 73 55 D2 D1 2D 6D DC 01
 17 CA B5 EB 0C 26 56 02 F9 56 FE 32 DD 42 95 B2
 34 AC D4 5F C9 47 84 C0 18 32 8A 2F CE 68 D4 5A
 31 2B 02 B3 0C 5A A3 7A 45 91 EA CC A0 D7 2C 30
 9C 78 4F 27 F9 5E 41 D5 CC 96 B8 47 8B F8 3D A8
 8F E7 3D 18 5C 81 5A 76 8D 94 5F 8D 5F 5F B0 C9
 F5 F5 3A BA 55 D2 6C E7 07 35 B4 76 29 C2 EF AA
 D6 18 7C 8E EA 2F 4D 68 19 5F 54 42 7E 57 8D 74
 7E 55 26 F7 01 89 0D BB A8 0B 8F DB 7D 33 CA 8F
 37 89 0E 25 3C 1F 89 A4 CD 01 39 56 0E 82 16 62
 FF 12 0C 48 C8 FF 25 5A AA 6C 39 89 C1 00 6F 53
 C0 00 9F 16 7C E8 91 C3 F9 5E 15 94 61 7A C1 4E
 84 A4 0C 27 D4 45 FD 03 8D DB 1F 1C 98 AF CB 39
 53 6B 11 3C 29 5B 09 8A 8F 69 28 A7 C1 F3 78 42
 D1 8E 75 FC 11 E5 F7 21 5B CB E5 09 63 1B 4F DD
 BD 37 B4 6E B4 A3 AB 45 07 69 69 6B 50 CF 8E 7C
 C7 8D C6 AF 39 3F E1 4F C5 30 18 6A 89 8E FD 5C
 C9 6D 60 5A 3B C2 ED 9E B4 06 C8 D4 FE 17 32 90
 64 7C 02 C0 8A 06 48 BE AB A4 AA 62 B3 76 6F E2
 33 62 8F C1 BC CA DB BD D7 15 78 8E 4C C6 D4 C5
 31 9F 02 8B 7C 68 3D DB 9D 8E D3 D7 9E 5F F4 1E
 8E EE 38 12 15 A0 03 68 E6 C9 59 9B 20 F2 21 36
 E4 0A CE 65 59 33 BD E2 D2 10 E5 C2 7A DA 41 35
 83 CC DE 4E AB 01 EF 3B 2E 51 98 FC A8 F0 AD 38
 F5 FC E9 E2 D0 BF A4 E4 D8 C8 B3 D9 07 6D 92 EA
 83 3F B7 91 00 BF 14 A3 CE 95 A4 63 48 B9 F9 5E
 E2 AE 92 D5 F8 BA 1A 47 51 96 56 8B C8 1B A4 CD
 2F 3A 71 22 93 14 0F 86 FD 8E 7E 2D 8D 33 F0 D3
 1D 42 7C 40 50 0E 46 8A A6 88 75 04 01 46 9B E9
 BE 82 83 66 87 34 96 CD 79 0E E1 30 1B A6 2E 70
 17 BD 29 CA 88 FA F5 48 0F 98 BA FE 0A 8C D5 70
 43 38 8C 34 74 6C 43 91 DC 5B D8 94 CA BC 2B 6A
 D1 A9 B1 8C 3D FB 2F 59 BA FF 1B 41 80 23 45 E0
 78 D9 14 2C 31 D3 94 84 CD 52 93 04 D0 96 34 53
 56 56 4B BE 7A 44 F5 75 49 DA DF F9 22 F1 10 0E
 B6 5F CD 46 F7 DB DF 1C C4 6E 61 35 48 F7 30 7A
 1D D2 62 70 76 15 36 B4 0B 14 16 C9 1C 01 40 17
 1C 56 7D 4E DE B3 B5 C5 7F 0A 57 1A 3F 8D 3A 49
 0F E6 73 F2 99 65 FA FF 78 29 4C F6 92 5A 17 9D
 34 7C B3 C2 C7 14 89 91 E2 89 D8 70 EC 32 0E 75
 E4 6F 6A 58 B1 0E A9 6E 8E F0 43 E9 0C E8 66 38
 C4 E2 92 83 DF 70 B9 13 F3 17 C7 D3 E2 5C 80 44
 D1 E6 9F C0 77 C3 B9 59 BC F0 7F FB 68 E7 D1 62
 D6 9E 19 F6 DB C0 DE 58 23 23 F4 77 4C CF 84 A1
 B7 6C AC 29 FC 63 7C AB 87 E3 14 70 70 A8 86 7D
 51 21 E5 9A A6 3D 81 70 BB 12 CA 8A C8 08 95 89
 DE 84 73 37 ED 58 7F 4F 75 B2 2D 9C BC 41 43 EC
 EB 95 93 B8 8E 41 4E 48 74 34 32 AB D3 32 2F EE
 20 48 5B A8 13 3D 73 9F D4 6D 28 7A C3 5B BF 50
 82 D3 80 34 4B FB A7 C5 2D 76 2B 7D 10 CA 3E 27
 67 75 28 E2 87 90 FD DD 98 95 87 37 4C 28 EA 36
 BA 22 D9 6B A3 72 8F 58 FB 12 1F 49 E5 9E 5C 78
 05 69 C1 6E 31 DF A1 7B C6 5A A3 71 2E 0B E6 4A
 AF C7 BA 01 8F C1 20 79 21 E8 14 FA F6 53 0C A2
 85 D5 6C 17 C3 DD DB 4D 83 DB BC B6 D8 A1 35 64
 A7 A9 F6 B0 F4 45 7B 75 85 F1 FA 9C FF 80 2C D4
 6B 65 66 FB 75 35 44 7C 20 D7 72 28 EE 8D ED B9
 18 33 CC EF 70 D4 5E EC A9 FD 55 27 98 F1 51 03
 ED 42 E4 AC FA 3C A7 7D 04 23 A5 D7 72 A9 42 84
 EF F9 47 0F B5 65 5A 4B 5F 82 89 33 F8 02 E8 4E
 72 CC 39 FB 34 AE 6A 3A 8E 26 D6 D7 35 B7 66 24
 F6 CF 5A 2A 2C A9 CC 40 5B DA 38 28 5F D7 BF F6
 F5 03 D6 7A 43 C0 18 57 21 90 C3 AD 7D 1E 98 95
 66 85 75 04 7E 03 D4 30 B1 71 CF 97 EE AB E9 B7
 72 C5 CE BA 92 5D B4 DF 2A 70 AA 98 A1 2A D1 96
 97 8C 4A CA 88 1E B1 77 23 4B F6 07 36 7C C5 77
 4E C6 93 F5 2F F8 86 05 25 65 AA 58 8A A0 4A 6B
 A0 E1 F3 A3 1F BD 73 CE 96 37 E0 E2 83 00 96 4A
 5F 46 D7 86 4A 1E 78 B5 93 2D 46 DC 1B 5E D2 0C
 B9 E8 BB B8 3F B7 D9 0D 63 66 AE 18 93 1C C1 D7
 69 34 95 A1 46 0B C8 C3 B3 B7 4C B7 75 4E 8B 11
 7E CF CA 1F 30 9F 7D A8 B2 71 84 1D C8 11 D8 7A
 E5 08 BE 5C 1A D6 AA 35 25 81 2C 27 41 AE 6F C0
 11 19 91 A4 77 80 1F D6 33 69 76 DD F0 2B A6 34
 F5 8A 36 69 4F EC FC 91 5A 65 34 FE EF BD 6A CB
 59 95 83 0A E4 8A A3 2D CE 4B BB 5E 08 73 2D F0
 A8 77 CC 36 AF 71 F1 96 5F F0 92 6E 94 A7 41 CD
 E0 13 29 E2 B3 AA 1A 57 6E 95 BE 43 46 33 17 A5
 7A 9D 39 3F 83 CA B1 F4 D1 BA FC 44 AB 67 36 91
 FC 65 58 35 FE 0C 70 3A 1B 4A AD 3B 93 8D BE CD
 60 A7 C6 27 D9 27 7A 9C 1F BE 27 24 38 79 F4 A8
 EC 70 1D 78 48 1C 3D 82 73 99 0B C7 0B AF 2F 73
 DF 7C 5E 72 C2 75 55 B1 FD BA 4D 0C 1F 2E 0D 0D
 1D 00 50 6B 62 83 21 29 56 3E 2C 27 CC 97 80 9B
 31 B9 64 16 BE EF 05 97 B8 D6 FB 56 57 77 85 78
 FA 2E 97 8A 81 15 DE 77 3E AB 48 AB 7F C7 05 AF
 67 FF D8 4D 29 7D BE 1D F3 70 25 AF EF 8E DC 26
 7C 79 99 7E 52 D4 01 72 58 9F E6 E7 59 72 1B FF
 07 0F 28 FB 76 15 CD FE 5E 7C ED E2 C5 DD C7 02
 47 C0 88 F0 D9 55 3A 51 75 06 4C DC 5A A6 5E F0
 7F 8F 5C D6 3F BE 08 0F D8 C8 B8 5E 1F 72 F1 7B
 06 F8 73 C5 FF 9E D8 14 7E 26 94 72 27 9A 0A C2
 9F 24 16 07 A7 E1 06 86 D9 53 60 DC 5B B3 13 DE
 D4 91 14 B0 E3 34 06 C8 25 B9 FE F0 E7 76 C2 39
 ED F4 15 D6 BB E1 22 C3 F1 B2 7E 15 39 CF 41 B6
 64 31 22 8E AB 93 47 0D AB 2F 0B A5 C6 FB F7 CE
 96 C3 61 F4 07 07 8E 67 48 EF 37 46 B0 7F 9E 43
 9B 58 A7 DF 80 13 0D 5A 14 61 27 2F 3E 6A AF 7F
 70 83 D8 57 51 20 A1 67 2E AF 65 03 F3 99 38 8B
 98 D2 20 7D B3 D9 F0 06 E2 84 9D 57 FE 1D F4 FA
 68 F6 8C C7 8F 4A 7D A9 6B C8 1C 91 F5 27 E4 E9
 79 2A 50 AF 09 86 54 A4 B8 E3 1E 7A 70 55 C8 2E
 DD 78 B9 1F CC 9C 2B AF E1 FD DE 19 89 A9 DB 6A
 F1 67 1D FB C0 24 BC F0 A4 B9 BF 44 D4 2F 5D C7
 E9 54 71 FD 01 7A 3A 3C BB 8F 82 D0 6E 1C 61 52
 E6 15 7F FB 83 29 F2 FF 25 4D E9 44 45 58 68 B6
 F5 93 89 B2 F3 41 38 C4 1F 3E 46 ED A0 78 42 04
 94 90 EC E6 4C 7D 34 39 77 07 96 B3 64 DE 26 37
 65 37 9F AE 39 4D 49 03 56 FD 4D 2E 33 C2 74 A2
 71 D5 04 02 B9 BA 14 D6 16 FA BF 4A 0A 82 84 60
 8F B1 A9 06 B0 11 C9 D8 95 62 7C 35 AC 8C 1B C9
 2A EB 6A F7 1D 9F C8 39 32 05 33 29 66 4A AD 31
 00 BA 83 E8 F3 4B 69 EE 8E C1 B1 D9 BE 11 C3 B2
 0B 57 62 08 5A 9B 9D 4D F7 72 AE F7 7E E8 5B A7
 33 B5 46 4F A1 1A B3 6A 05 EB 52 CC 9F A7 54 D2
 55 FE 14 69 3F 13 36 60 69 FF 5A 37 FC 53 EF 48
 AA 83 B4 BF C1 CC 4A 13 15 3C 0A 0B 6E CE 6D 68
 AA DC 8F 62 CE ED EB 49 E5 02 35 5D 0F EF BF B2
 E4 18 DE 48 76 73 71 56 07 A5 C2 03 C9 F9 1A 69
 2F 26 55 D5 AF 96 1E 42 B7 A2 9F 68 10 3D 47 76
 CD 85 61 95 12 A2 00 56 E2 39 F3 F2 19 C9 EF F0
 D2 43 8F DF 36 8A CF 1B 30 5D D1 B5 B1 15 60 61
 1B B3 ED AE B4 9E 0C 5D B1 4F 27 F8 C8 FC 35 4A
 95 BF 50 E4 3A 5A 04 34 63 3D 20 13 6F F2 5E BA
 CB FA 6E 40 F7 D0 35 A1 EC D4 D7 F9 C4 2C 93 41
 F1 EE 40 28 4B 68 01 27 E7 6A 91 60 D2 20 3F F5
 51 6B C2 85 F7 7C 0F C9 51 FF 51 6A F4 5E 42 35
 37 6E DD 48 31 5A 30 70 5C 25 A9 E6 D0 B5 04 D4
 CC C6 F2 C2 B8 86 AF 8C 29 39 CA C2 2D 0F 52 20
 44 04 5C 68 0A 27 D3 8F EF E9 4B 7D 2E B0 1E 4C
 F3 BC 3E 9D 1C 0F B6 D1 37 5B F7 00 65 98 9A 23
 8B F2 F3 B8 58 1D 24 B7 AB 30 AB C3 6A EF 83 DE
 8E FA 1A 18 76 86 65 3C 3F 6D CE 00 C3 70 96 02
 64 A0 64 A0 51 53 E5 92 3E F3 6E 64 97 0D 4D 86
 33 AF E7 74 5D FF 7E 64 23 9F E6 B2 EC 91 EB F2
 A8 1B D7 E4 90 E2 99 25 2D 68 BA 10 40 2E E0 4A
 C8 A7 83 8B 53 F6 AD 62 07 F1 CD 2E 9D AC 1C CB
 B0 D0 B3 23 79 A9 93 1B 58 B6 69 93 66 CB 4B B5
 34 4B 16 3A F6 CE 12 D9 FD 61 EE FB 03 CF B5 3C
 AF 3A 7E E7 92 EB 19 32 02 A9 88 77 AF 24 91 0C
 06 52 1C FD 1C CA 3B E8 B6 3E 69 46 43 61 88 76
 11 E7 66 6C B8 1A 8D CB 45 E5 BE 19 60 EF 99 00
 E0 BC 5B 04 E7 1C D9 07 F7 1E FC 19 62 E8 B3 D1
 9A 34 AA 76 4D 72 96 6C 9B A8 19 0C 84 C6 99 6D
 03 81 E8 C9 C2 DD 95 B2 3F 5A 56 42 75 9A CA C7
 77 88 E9 BC C3 F9 84 FF D9 E0 3A AE 2C 0A 3F 63
 D0 64 D8 E0 7C B4 FE 6C 5F C4 BA 79 28 66 30 D2
 9B D2 47 E0 B5 AC F2 EA 10 26 E0 B3 03 80 1A CC
 3E 16 B9 70 AA E5 0C EE 49 0F BE 48 F7 F2 6E 47
 25 68 3D 63 95 9F 0B AC 4C E5 64 54 1D 6E 2D C7
 F0 CA 7A B5 3D 5C A4 42 9B BE 45 09 8D 37 7C 3D
 67 18 75 DC 30 E9 62 6F 82 8B C3 2B 3C F6 D6 97
 E5 F2 43 C2 A3 D2 C7 5A C4 D8 56 AF 7F 62 B4 D5
 78 37 7E A4 21 1E A2 CE 9E 87 13 DC BC 2A 56 69
 E9 AE B3 59 EB 27 83 E0 B3 CC 35 6D D7 ED 64 CF
 FB C9 0D 0C 96 6B E4 50 32 54 57 66 45 2C A2 60
 B9 20 E2 87 EC A1 C0 22 BE 47 82 CC 39 55 9D 17
 ED 47 DB 4F 19 E9 A4 F6 65 25 9A B1 86 FA 53 FB
 54 48 70 2D 10 8F E9 60 1B DE B4 D4 98 2E E0 93
 19 49 F2 4A 2F DB 6C 40 2C AF 94 F4 FC B9 5E DD
 86 22 32 16 3F B2 38 48 2A BC DA 92 A9 57 DB BD
 E0 D4 AB 55 AE 58 E8 73 EA D3 22 03 85 8B 54 D3
 7A 33 EC CD C9 C9 BE 35 77 2A 70 65 8C 68 89 91
 34 0F 4E 70 68 DB 0C 89 2F 6C 97 1E 59 32 D1 D3
 33 0E F0 79 CD 2A 06 6D 96 EB 97 50 76 80 B4 E2
 D2 43 35 C7 F1 00 D8 CE 35 1C E7 0C B1 A1 18 72
 B0 01 ED A0 F6 8B B5 A1 2A 90 EF 0B 9C 9B 81 C9
 B8 4F A6 32 B8 17 95 78 5C 3F 45 C4 63 FF 6F 40
 F6 77 25 87 12 E9 54 3A 47 2A 2D 51 B2 E4 64 9E
 A1 3E 82 2D 29 99 6E 6E 35 D9 B8 A1 18 B4 5A 9E
 94 EB BC 3C 72 31 B9 21 D0 F9 3A B0 CE B2 15 8F
 C3 FE C9 45 2A 49 AB 43 02 F6 89 E0 AC 42 A1 45
 13 C5 9A BE C3 44 0D 23 74 84 E0 CF 92 FD 02 0C
 B0 6E 5F 94 FD C5 22 76 70 9B 59 5F DB 7D 83 CC
 CE B8 64 BE DF 35 84 2C 2D 74 4E 7E AD 0C BD ED
 87 A9 29 35 31 D0 A4 3B B9 10 40 77 B8 2F 3C 4F
 44 B0 77 5E 07 C9 B7 B6 94 6B D0 47 62 F2 5D B2
 5F 90 2E 6C C9 3D 6F D4 C5 6E 33 1D 81 15 7A C3
 36 7B AA C1 B8 9B 1E 79 A5 99 3C 42 F0 CF BD 53
 5C A4 94 F5 3E B2 BD 5B F4 8B 14 B2 EE 53 06 23
 92 5A AB B6 8B 74 7B BE 2E C5 6E A0 35 65 03 0E
 88 00 21 A9 5C 21 D4 60 8D 78 9D BA 4D CE 75 9D
 E0 61 AA A6 82 DE C9 5C 91 20 EC 1B 39 49 FC 42
 76 7B 6A 74 FD EA D9 F9 9D 89 11 B1 DC 7C 0B CE
 D6 ED B5 2F E0 24 4D B1 A1 36 FA 71 5C 34 46 4C
 BA E8 61 F1 97 5A 4E C4 79 EF C4 B5 70 B2 60 43
 AB 91 74 8E 71 36 7F 91 D2 AF 89 61 D8 9C 9D 37
 E0 56 3D EC 32 FF B4 EB 3C B8 0E 96 EF B1 81 3C
 15 39 98 BD 66 FE 62 F6 C8 4A 58 A0 EB 63 EA 87
 EF 77 9B 24 59 50 95 D1 C1 97 80 A1 A3 69 AE 01
 60 15 86 EC AD 9D 3D 64 1E A6 61 D3 7F FA 80 7D
 87 C0 A2 F1 5D EF 3B 12 91 3C 27 CD D8 90 DE 6D
 DB 93 A4 8E 13 C9 B0 41 0E 84 B4 D6 27 AE E6 D7
 82 55 77 99 B5 B2 5A 61 51 91 D4 1E 4A 8C 9D 5E
 09 31 19 15 24 C8 30 9A BE AE 1D BB 7A CE AD F6
 7A BA CD E0 19 1D 5A 33 D2 36 A8 3F AA 86 C0 0A
 36 0A 95 E1 1B B3 4A 6C 04 A4 6E 36 58 59 28 83
 F5 1D 85 D6 8C 95 9D F0 61 F4 0F 26 32 51 45 9D
 84 45 4C 4A D8 81 75 DE F6 9F 34 28 28 94 77 D8
 23 A2 9D AC 83 29 8B 43 05 21 84 3F C5 7A 0E 5B
 DE 51 0C 15 85 C9 22 BD 25 1D 5F 30 A1 07 84 F3
 78 6B E8 8C A7 31 F6 CD 30 8E A5 E9 6F 9D 4B 3E
 3F BD AC EA 13 AE A3 24 E2 D5 E7 E0 C7 FE 64 0A
 94 9B 2C 5B CD 24 0E BC 1B A6 73 60 90 A1 20 27
 FE 22 66 AD FC 5E 2D C8 AD 54 CF 7C 0E 39 44 A1
 54 6A 64 66 63 D2 77 5E 2D 1E F8 8C 73 18 77 6C
 9B AF 23 5D FC 6D BC 4B EF CF E8 68 C6 E3 45 15
 32 E3 47 91 A2 5C 33 21 99 82 FC BF 1D 0A DF D2
 73 18 78 FB 63 86 E2 26 18 C9 BA BD 2B 84 75 87
 9B B4 32 94 8A FF 07 84 B2 48 5D D6 13 E6 18 03
 74 87 58 F8 A7 7A B5 3D F6 F2 5F 9F 67 44 D2 8E
 BD 37 FE 8C AE A8 20 A9 AF F6 4E F3 A5 11 AC BA
 3E A0 28 3E DD C8 BD A8 57 D6 06 A0 E8 A0 B2 B1
 30 18 FE 88 E5 A6 4E EF 5D 75 31 C9 49 0B BE 67
 F2 C7 57 A0 79 B3 1E B5 7A E2 28 6E A0 C0 D4 90
 C1 75 6D 15 29 32 E4 3B 82 92 51 5C 79 FE 41 F3
 83 13 77 8D BF D0 2C 40 AF 1B C5 77 F9 58 19 4D
 F8 31 BE D0 BC 78 23 FF 9E 52 33 FD E6 54 90 D3
 DB 59 C2 AA 57 36 E2 F6 91 FE 22 B6 2E A9 2E DC
 0E D0 B2 62 F2 46 F6 DF 7E A1 17 D5 FB BE D6 A6
 CA 83 E5 7A 98 06 57 C4 92 79 D3 93 8A 48 E3 F0
 15 C3 E6 C9 24 4E 42 14 98 67 C2 7E C6 46 8B 9A
 DB E6 A2 A7 8A B4 F2 A6 ED F7 79 D9 6C 9A 25 78
 1B 62 7C 18 EC 69 2D 1C DD E8 F3 51 17 6B E6 48
 7D 86 09 D6 4B 4F 3C 26 69 50 02 86 8B F0 05 62
 0A 8F 51 40 2F E1 CC C4 CB FC AF 9E 4C DB BE 3B
 21 A3 AC 03 FE 6C 75 41 57 FF 0E FE 1D FD 6F 26
 C4 C0 EB 7D 92 BB 58 75 08 56 31 ED BD 93 F3 B9
 A1 2F 67 72 04 07 63 48 49 95 F4 B6 5A 24 14 77
 1B E7 D4 AB AA 9E 8B 97 D1 68 86 AC 0B B1 DD A1
 F5 64 8F CE 9E E8 1F 6E B6 77 1B 07 4D 70 EA 29
 73 45 30 DE 33 66 97 ED B0 46 AB 96 E8 58 41 66
 20 07 58 5C 54 DE 6C 10 63 45 2C 97 C3 56 64 13
 41 1A 4B A0 6E 6A 52 46 93 A1 30 34 B7 48 AB A1
 6C 10 85 EE 97 0D 8C 5B 2A 99 D3 52 77 13 1D 8B
 10 09 12 BB 22 07 DA 22 B7 7D 03 A3 60 47 9A 16
 D7 2E B5 35 10 BF D7 62 9B 44 74 DB 87 89 C5 2B
 44 DA DE A3 36 BF 74 53 AE A9 A5 55 26 73 08 47
 D7 47 58 41 FA 73 3A 89 9B 21 A5 E5 D2 65 C5 B3
 CC 01 C5 71 44 35 E4 1B 07 0C 32 2F 61 7A A1 E6
 DE 1A 4A BB 68 64 2B 3E 2F 0A B9 8B 94 A2 2E 78
 7F 85 EC BC C0 DF B5 BD BA 32 01 E8 FB 38 85 0A
 9C 5B 4D 52 76 AE AE 15 90 81 73 39 5D 8A 92 3F
 73 18 97 F8 58 3C FC 89 77 6E 59 69 B0 27 1A 36
 85 17 A3 99 E9 31 84 8C 92 1C 2B 5E 11 25 94 44
 E5 77 EB 54 66 F8 96 B6 A5 8B F1 AA 70 01 6F 76
 24 ED 5C A1 16 4E 3F BA CC 14 6D 57 BB 8E 29 00
 F3 BC B1 83 08 BD 0F F2 5D 5B 19 FC 1B 2E F2 90
 FF DB 73 22 BE B0 21 02 11 88 DE BA 64 E6 51 53
 DA 53 7A 5C C6 8B 05 B5 7C E6 9B 00 87 E2 13 82
 2D 8B 8A 64 E9 E8 43 C2 E1 FC 58 1C FF 43 A4 71
 2B 50 93 74 D7 36 44 BE 4C 4D F9 BB 4D 3C 46 CE
 87 EC DF 63 B4 7D 95 54 CC 5A 77 75 9C E5 C3 6D
 3B 81 4B 2B 1F EB F7 9F 12 C3 F1 FB 79 AA 3D 15
 7B EB 79 E4 D1 75 BB FF 2F D2 11 5C DF 77 87 84
 AD A4 97 E7 A4 8B B5 BE 2D 46 B6 24 A5 C2 DF AA
 AC 46 17 1E 75 22 42 48 67 06 96 13 80 70 F7 AE
 D3 3E AD 7C 7A 3E 00 4A 7F 21 1A D0 44 F9 EA 3D
 D1 88 29 DD EA 79 A5 1E 20 22 E3 1A EF AD 11 05
 79 12 85 35 38 04 65 BD 3F C7 E2 30 38 4D B8 7A
 16 73 C7 05 33 2C 5B A6 C6 5D 83 6E 5E AB B5 1B
 F0 C1 54 A2 84 83 EE 2C 7F 84 12 95 24 08 19 83
 73 0C E2 0C 8F CC 77 50 57 7C 9F 2D 69 A5 8D 3C
 E0 85 AD 23 45 2D 27 EA 73 2E 68 24 25 AF AE B0
 17 85 64 8B 35 34 11 20 15 9D 0E A4 70 3F C6 4D
 BE A0 B6 3C 9B 96 71 AB 10 F6 B0 D1 D0 21 95 A8
 F8 68 0E 7B C6 6E 34 6B B8 35 0F D4 00 39 36 E1
 93 EA 91 2D B0 5B 5E F7 62 37 BB 0F 58 63 B4 CF
 7A 65 76 9C DE A8 0F 65 39 27 A6 30 0D EE 5A 3B
 09 B8 12 94 76 14 CC 49 A8 17 7A 0F EA 78 F5 6C
 6D 7F F4 79 03 07 B1 E4 E6 3B A3 FF 4D 1F CC 4D
 BB 9B B6 7A 49 BF 81 91 36 D3 01 EB 5A 27 10 3A
 D6 5B B9 78 F9 1D 8B 22 E7 39 63 8E BD CC 64 4E
 88 89 EF 30 AC 3C 28 47 6B E1 DF 0D 64 DD DE C6
 CF 77 95 38 C5 CD 93 E1 06 7C 9F D3 6B 4B A4 A6
 8F 40 94 8E D8 14 89 3A 33 64 92 8D E1 9D 80 20
 7A B4 BC CF EF 35 A7 D4 4B 4E A4 32 97 86 7C FC
 7D 9B 8E 9C F0 25 49 AB 7F FC C5 2C C6 23 3B 30
 FD BF 92 D0 8E CF 49 36 8D 6C 7C C7 1F 1D 1E 81
 82 A8 BB 6D 3B D1 B6 F9 B4 3D 36 30 7A B2 DE DC
 1A A9 3A 17 5E 04 46 38 EE C5 E4 49 AD EE 56 93
 F7 F8 D1 72 DB E0 5D EE CF A8 3C B2 B3 07 C2 95
 3B 18 AD 82 F0 01 BA 57 DA 80 96 79 5A B8 CB 82
 F7 A2 F4 A8 43 B0 94 86 3F A2 87 22 88 01 B5 1D
 2C 3E E9 90 61 76 C3 D1 38 36 FD E8 9A 0E DD 97
 D3 4F 03 8B 1D 63 38 E3 07 9D 5C CC 3B BE BB C2
 57 CA 6B 5E 28 BA 00 78 15 41 B4 25 18 27 49 DD
 54 4C 19 DE 2C 14 0A 65 71 8D 99 2A C4 4F C0 BB
 6C 1F F1 C0 CD A2 7A 0B EF 94 B4 EF 2C A3 7F A2
 95 7F 12 F3 30 B7 AC 94 31 6A DA B9 35 95 E9 D7
 71 58 53 2B 4C DF 0E DF E3 0D A6 58 32 8A 5F 13
 53 CF CF A2 37 9E 71 84 DA 0F B6 CB 47 11 E7 DF
 BF BF 83 F1 D3 B0 9A 87 5D E3 AE AF 7D D7 3A 85
 B4 6D 6E 13 CA 21 D5 C2 ED AD 42 27 67 6E 3A CE
 D5 9B CB BE C1 4B F7 1F 84 D7 34 4B B3 CF 1C 46
 98 08 5B 94 57 37 76 A7 35 DC DB 25 F5 DA 4C E2
 43 C9 E5 9E D8 AA 78 19 AB E0 3B 49 C1 30 0D F1
 7C C9 69 B2 03 17 BA 4D 67 4C 4E 38 13 70 0E 2B
 B9 AC D5 D3 D3 14 1A 6E 35 71 26 99 CB 38 04 2C
 30 19 E1 0A 36 9F 4C 9E 83 C3 03 1A 61 2B BD 2B
 07 4E 5A 14 5B C7 F0 E2 FA C9 F8 9F 27 71 93 97
 8D CA 8C 7C B0 29 45 07 4E 79 17 08 D7 0F C5 CC
 D5 A8 18 0F 5D 56 1C 02 4C 03 65 90 51 61 E4 C0
 57 AE F6 33 61 BD 23 CA 74 A7 2F 38 D7 46 5B 69
 0D 98 87 CE FD 55 77 E0 D4 28 E1 B4 5F 6E 25 6D
 70 1A E0 FD 8F B2 71 2C 71 6E 4F 79 BA 6B 50 6B
 F4 C1 3F 88 C3 2D D5 AB E7 EA 24 F0 5C AC E2 4F
 FC 0F 0F B7 43 97 80 B6 44 81 AF FD A5 03 9D 4B
 40 0D 6E 2A C6 5F C7 0B 8A 62 14 B9 45 92 F5 10
 EE 7E 81 A8 71 A0 72 B0 6C FF D0 47 AA 4D E4 F7
 C0 D6 B6 F8 23 E8 29 0E B6 A0 A1 A1 BB 2D 2A 08
 8F 1D 42 0C A9 25 AB 53 4C 33 2E 3F C3 7C BD E2
 DA EE 53 E1 C8 3B B7 22 EB 8C 19 C7 18 81 C2 AB
 82 D3 15 5B D7 83 3D EC 26 23 63 7E 3F FE 25 F8
 77 97 47 C4 69 48 AD 27 4E B1 1E 15 15 EF 6F 6F
 05 7B 5F D8 5B FB F1 03 E7 1B D4 E9 48 53 98 67
 99 D4 A5 14 B6 61 76 B4 7D D8 A3 7F 34 4A 2F 29
 58 4C 43 82 A6 4C D2 18 E0 F7 01 8A C7 21 F2 4F
 6F 40 B2 A9 20 99 F1 20 2E 40 F1 BB D6 AA 89 54
 C5 06 74 A8 F3 3D DF B3 C3 81 61 E9 FA 85 5B 01
 80 C7 D6 E8 6B D0 66 7E 2D 7A B8 C3 3C 05 69 BB
 AE 65 82 C2 BD 72 DD C3 4A DB 9A FF F8 40 48 32
 1C 5A 7C C4 70 45 72 8D D0 8E 28 33 6F 7F 90 D3
 30 65 39 7E D1 1B 56 E7 AA 20 59 0F 7B 60 7F 1D
 27 56 CD 98 83 67 DB 5B B0 EB F8 D5 5B 67 C6 1E
 19 1F 67 4A 9A E7 DC 53 9F 5C B3 08 24 3B D8 91
 2D 6B E0 31 05 B4 D9 73 9C 50 19 CA 73 17 BA 29
 2A C4 2C 33 A9 28 E7 7F 84 DE B1 F9 79 A4 22 CA
 F1 AE FF FD B8 38 CC DA A9 85 46 BA 5E 6F 17 5E
 5F 60 DD 01 4B 91 AE 80 FE FC 14 12 67 9C 76 55
 A5 0F 44 23 A5 98 E5 E3 C6 24 47 90 2E 6A 20 24
 CD EA 1A 08 88 AC EE D3 D4 4B A4 2C BB F3 D6 0A
 27 75 4D C4 3A 3A 40 D7 8F 7A 84 57 47 60 95 A9
 B5 B3 70 E0 46 F9 63 A7 25 D1 BF 75 83 30 C5 6B
 99 47 66 57 81 F6 DA B2 36 E2 F2 F3 72 D5 86 E0
 08 25 C1 8E 19 44 A6 13 89 52 25 07 E1 49 B7 01
 57 93 7E 6C 2B 8C 47 64 BD 83 A6 F7 02 48 F8 88
 11 AE AE BA 80 DF FF 8D E8 7C 9B E0 FD 15 15 E2
 F1 88 AE 85 2D 12 BF 3B 6C D0 BE 47 2F 6B 06 4E
 BE 4C 03 75 4C 17 EA 63 9A C7 4E D0 10 98 8B 28
 F6 59 89 05 8C CD 32 5A FE D6 5C 10 54 FB 7A D2
 E6 E6 B3 7C 18 1E 2F 39 4A 39 3E 84 D6 DD 20 A4
 E6 4B BB 01 E5 51 9E 70 41 6A 9F 1B 67 D0 1A 1F
 6F 6B 33 20 82 0A DF 77 45 55 C9 C2 BB 49 56 3C
 11 8F C9 2E 12 8E FE 7E D6 2D C1 F6 19 EF 50 33
 24 27 BE 36 60 6D F2 51 70 97 57 FC 3B 86 92 41
 F1 E4 B6 AC BC FD DE E3 84 5B C5 C2 B0 22 88 08
 50 F1 18 36 BE F6 AA C4 E0 5A 6A F7 DE 32 AD 7B
 11 EB AD 1E 88 25 CE 77 36 CF 8A EB B9 C3 2D 1D
 B5 1B F1 AE 0A 2F EF E0 DF C7 CC 7A F5 1A E6 4A
 74 4E 57 FA 27 25 5B 1C 20 C2 C6 41 54 81 E6 5F
 7B 43 12 E7 C5 F0 69 77 0F 4C D6 11 29 C3 66 CB
 23 17 09 43 FA D5 E5 96 82 7B B2 F9 42 48 56 BE
 6F E3 11 D1 98 FF 1F 33 B0 08 C6 61 19 6D 11 0C
 69 8B 24 04 77 15 8E 42 3B 18 8E 4C 2E B5 68 89
 9D A2 48 4A 95 63 E6 DF 75 EF F5 4D E7 FF 00 F0
 E5 9A 19 91 DE 04 56 4D FA 92 14 1B 45 E9 13 F2
 5A 11 31 98 53 B1 E3 D0 CF AC C8 36 4A 70 41 47
 F3 56 AB 37 31 A5 D6 88 B5 CB 1F 03 6B FE 4A 97
 3D B8 A3 0B 2D EB EE ED 49 BE 5C 3D 3A 5E 05 90
 CA 67 CD AC B4 FD 2C DD FF 1C 1E B8 37 D1 FB AC
 B3 E8 6C E0 CC B4 F5 D1 21 C1 5B 56 D0 11 69 06
 DA 66 FD 9B EF FA 31 83 F9 1C DC D2 8E 2C 8D 93
 1C 83 BD 14 3F AC 08 69 CB 06 AF BA 2C BC 05 01
 25 75 3E 3D F2 7F 0C C3 8F 67 00 09 27 0C 70 8F
 2D 1D F7 C4 C0 68 94 13 F8 28 F7 45 00 E6 D9 B5
 18 D0 41 59 28 D8 86 5B 41 D9 09 5B 87 23 2A 5F
 ED 4B D3 2E 51 A3 53 B4 4D D3 09 34 64 68 9F F3
 C6 0F C1 5B D1 25 95 89 AD E3 FC 38 04 23 E2 A7
 9B 66 E5 4D 66 55 1E B4 C1 79 F6 58 A1 C8 45 A9
 E2 D8 F1 9A 85 3D 31 28 84 9C 5B ED 13 98 6C 6A
 21 D6 40 43 B7 4A AF F4 60 2B C7 96 51 C1 F2 7F
 8F C7 82 EA D9 D0 26 D5 98 6F B1 14 BB 49 D3 F4
 74 DB 25 99 6D E9 22 D1 D8 3C D1 E8 44 9B 9E B2
 81 0F 5A C9 AB 71 7B D5 B4 DF EC 40 A5 FA 36 6F
 60 D1 7F EB 32 7A 4E 56 EC A3 40 44 F0 FA 6E 52
 6D BC 9B 8E C3 D7 09 BD 35 BC 0B E9 62 BF FC B0
 50 E9 48 0B 26 63 B1 8A 47 2F 60 BA 60 DF 6F 94
 81 5D A5 F1 FD A8 1A 57 2D 2F FB FC DA CF D7 C3
 05 82 2E CD 27 16 1A 87 26 36 5C 8C 97 10 9F C9
 9F D7 E9 AF B2 F9 61 0D 71 98 90 C6 37 22 47 53
 57 D5 EE B1 F2 DE 19 49 73 25 35 A0 E8 F6 69 67
 C0 69 32 ED C3 86 5A CF A5 E2 7A AD 57 18 36 3B
 30 31 F5 D3 C8 41 0A C8 44 D4 52 9B BE D7 8C 7A
 8D E5 79 30 05 05 F0 5C DF EA 76 C3 85 B9 8C 1A
 A1 E8 07 FE CB D4 89 89 81 DD 1A 1A 09 0A BB 45
 A7 E9 25 3C 11 47 E4 ED 1E 86 92 F8 FE 59 67 D9
 C7 CD B6 2E B9 B3 F3 D6 E7 39 AB 68 C3 45 19 CC
 93 5C 55 97 88 59 F3 11 EB A3 A6 F6 A4 29 6F 1B
 DE EC E6 22 2A 02 49 96 AE 0D 70 69 0D FB 49 3A
 7E 54 A1 8D AD 94 64 F9 CC 4E 5B 3B CD 6A 28 32
 D5 B4 A7 DF 0F 19 F9 0B A2 48 BE 7C 0F 71 D6 FF
 24 39 98 71 CD A7 96 D0 A9 F5 FF F7 C1 29 7D 13
 E7 EF CB 80 8F E4 86 0C C1 1E B6 98 5A 55 3A 1C
 3D CF B9 DD 88 5F EE 3F AC D7 E4 30 9D A6 03 EB
 7A 46 37 8C 2E C1 C9 FB D2 06 B9 EA 34 4D C3 3A
 B5 D7 77 5D 80 7E 42 A3 7C 15 6D 94 C9 A9 1A 6B
 8E 1E E8 3A 02 33 87 4B EB 89 13 E0 65 31 4D 0B
 12 EF 93 F7 E3 77 F7 B5 EC 48 05 4D FD 93 D5 70
 F5 76 A7 D7 52 43 AA 4F 1A 66 48 DD F7 48 04 01
 E8 69 55 D3 3B 6E A8 47 F8 83 FE 77 37 05 64 76
 A9 89 11 08 53 3D 9C 15 FF 07 A8 E4 93 A3 B2 FD
 5D 41 46 51 C0 C9 F0 9F A9 35 76 03 91 18 FD 2F
 A1 30 8B CF 46 B6 C0 A9 41 82 4E 0C CB 81 2B 3C
 18 94 07 23 25 FE CB 5F A2 AB 97 34 87 25 E7 59
 8B 68 12 97 AF AF C1 1A 5A 90 64 52 4A F2 2D 8D
 0F 55 0A E4 D1 7C DF F4 1F 1B E0 0A CB 91 B3 CC
 A1 5E DE CE 88 D7 1F 9B 4B 15 34 83 AB 1C A1 FE
 21 D2 E5 4E 4F 43 3D 9F 7A 0A 68 06 BB 83 8D 76
 F4 D3 62 97 FD 16 58 EB 46 42 B7 24 A0 76 AE AE
 3C D8 65 F2 26 78 E1 4F 9F E4 06 DA 0A 41 E5 2F
 D5 82 63 F7 B4 78 C6 7C 5F DB 64 ED DB EC 04 53
 D6 AA B2 79 BC 4F 30 DF 2C 31 D0 29 63 9F 16 CD
 91 83 58 0E 4E BA D4 52 D4 F4 38 CC CD 02 92 03
 47 EB 6C 87 18 FD D9 49 18 9E 1E BA 72 C4 E0 A0
 F8 CD 7B A4 37 87 E5 6C 98 CE 94 0E 5D 25 CA 11
 07 A2 76 C4 1D 56 08 CB C1 0D C4 E1 D3 16 9C B8
 F6 4D CE C4 3C CD 49 E7 58 0B 75 01 0A CD 90 BB
 44 CD 30 E7 10 37 62 5D 09 4B EF 11 13 15 59 B0
 94 B5 AE 5C 31 8D EF 30 A6 CF 97 02 B8 69 01 0D
 ED F7 CA 5E 88 62 FF BD 03 46 19 8C 85 8C F5 C9
 C1 F4 12 9B 16 C7 24 1B EC B0 C7 4A 8F 87 BA 35
 0D 6C B2 83 CB 6D 78 CC EB 87 05 D0 44 77 35 8D
 5E 52 CB 4A C6 46 C4 5F 76 A4 6D 5B 4F 88 44 4E
 69 F3 70 3E 52 47 D5 62 E3 73 AE 4B 49 EB 6F 3B
 D2 94 55 BC 9D 2B 29 A5 3C 05 C9 31 EF 51 09 A4
 B4 05 09 88 41 F0 52 57 11 A6 AF DE E3 C5 98 F7
 48 B6 D8 74 1B 06 0F 5F EF A8 D0 B4 62 0F 26 41
 15 CB C4 75 B8 47 CB C2 0B B9 59 D3 97 C7 DF AD
 95 1D E8 8C D8 B1 BE D0 DD CD 37 B0 C0 9D A8 EF
 69 08 0F 0B 64 04 34 51 D3 A9 DF 43 FC 2B CC B5
 2F 3C B8 D1 DD 98 4B EA 7F C4 8A B7 66 94 D4 62
 11 F7 F3 54 05 A1 FE 24 A1 7C FA 2F 89 59 26 7B
 B2 57 48 DC D2 B5 05 26 A3 28 2B D9 04 F2 4A 5A
 52 4E DB A0 53 E8 06 39 A5 2F 8E 56 43 B0 2E 25
 E6 03 6E 49 E0 B6 05 41 78 2C 63 1E 73 F3 FF CA
 3D 8D 0F 9D E8 FB 28 ED 3E CB 18 72 A1 D8 2E 28
 19 EC B0 6D 37 90 A7 10 FA 0A 7F 10 43 3A 81 3E
 0E 73 33 76 57 8A B4 ED AD 6E 9A BB 74 77 85 A7
 13 E5 10 8C 61 C8 4B C3 36 19 A5 AD 3A A7 28 2C
 C6 8A C8 14 3A 29 76 36 1C 31 B9 46 2B 41 BD EC
 5A 70 BD F0 50 FD 00 D4 86 63 FA 1C DB 44 36 41
 58 B3 04 28 14 9C A3 E6 A6 A2 0B 94 D3 99 D2 7D
 24 BA 1A 09 97 89 05 66 5F 04 79 C8 1E 9C BC 57
 C7 3C 77 E2 A0 F6 CE 43 3F 70 8E 70 50 59 14 41
 8A 99 E3 FE E2 59 27 F2 7A F3 E8 75 4A BF 38 31
 93 63 66 67 3C B1 17 B0 96 74 71 52 24 6A 5D 26
 CB DC 48 78 48 91 E8 7F 6F 07 1E DE EE 5F AB 92
 F8 87 36 C9 5E 30 03 85 B6 DB 83 2E 7F 71 F4 CB
 C7 E3 C6 9C 17 FF B9 83 AD 56 D6 D0 31 D0 27 42
 F9 BF F0 25 D0 61 6A D3 4B C0 29 8D 21 13 41 D6
 98 06 F3 6E A1 7A 58 83 A6 FE C4 52 78 66 8A 86
 46 00 9D 19 64 22 CA 73 61 1A 6B 50 C2 25 5E CE
 30 A6 C8 D3 DC 21 33 9A C5 5F A4 67 27 B2 0A 52
 C1 1D B5 68 5D 65 4F F9 DB 63 FF 72 49 56 D8 97
 34 5B 29 40 5C 3B 4C E9 8B 34 62 C3 FF 0C 3D 4E
 CE A4 E2 C7 78 F8 4C 77 CC 6C 94 A4 27 66 5E DA
 DC 5B 19 B8 67 B5 8D 3D 0C D3 CE 3A 57 7B 1B 55
 88 1B 95 68 D7 7A 8B 9A A5 AC 00 27 F4 34 1E 32
 12 F9 B8 9B 82 4E 2D D6 9E E5 85 7E A9 09 2B AA
 50 FE 31 0D CE 27 E0 51 F8 19 F3 86 CE 3F D4 E4
 0A D7 58 BE 8B A1 D3 88 7B AA AF 57 75 BE BB BE
 DA 7C 67 B1 27 FB F7 AD D5 AC F0 F0 F7 B2 2E 06
 E7 16 41 A7 E4 33 D7 4C EA 43 37 5E B0 15 AC C9
 57 82 12 6F 81 3C D4 59 84 9C EF DE 44 4C 1E F7
 70 66 E2 AD 0D 35 E8 D1 33 04 66 E2 0D BB E0 2D
 7C F3 64 5C DF 0E E7 13 7E 73 25 A3 E3 89 F3 EF
 2B 87 3D 11 94 DD 4A B9 DE 66 A6 B8 DF AA 29 AF
 33 60 B0 A0 03 AB 18 E8 6F 06 21 60 6B F0 F0 29
 6E 22 EA 6F AE 96 51 79 7F 2A 4B 62 C8 0E 66 98
 71 63 98 4E D8 81 A4 6C C8 84 7B AB 8F 75 57 21
 40 00 5A 28 4A 02 EF A7 32 1F EF E5 78 A9 94 BB
 F3 E5 45 D9 F3 CC B5 E7 C1 A0 6D AB 62 AD 78 46
 00 EA 23 0A DB F6 CB 11 BF A4 49 EA B9 BA E3 57
 E3 D1 C2 DC 11 85 E8 25 CF D7 44 7E A6 8F 55 04
 C6 B6 39 64 0C FB 9C BD 7C 11 4F CE 30 6E 6D AB
 61 08 24 A5 C4 8F 5B DC 4A 40 19 0A 3E 38 89 AA
 DB D6 7A A7 73 CD 9C D6 01 3B 43 62 A1 DC 11 7F
 2B 7A 0B D4 7D AE 00 C9 CA E2 D3 5B C7 D5 5C 4F
 32 F6 8F 19 6F D5 D4 3B 76 1B 54 B4 0D F9 C6 FC
 D2 A1 42 DB 01 64 E6 C7 B8 49 24 34 7D C6 B8 47
 BD 48 54 4E 0D 09 E9 B9 50 58 FD 8B 9D DA 20 79
 AB 90 95 65 45 65 A5 EF 5C E3 31 4D 53 F2 FB C4
 02 75 60 8E 81 5A C9 BD 10 8A 6F E2 DB F9 D1 FA
 27 47 85 89 1F FA 3E B3 2B 94 6D C8 53 0C E0 40
 1A EB 7B 10 91 A1 52 D5 C4 6F C8 D9 9C 66 CB 3E
 50 17 60 EA 7C 34 23 EF 4B ED F5 2C 91 08 53 1D
 E9 44 EE 13 7A AE 7D 46 EA E5 B3 04 A3 CE 35 2B
 36 23 BE F0 8A 32 24 6F EE D4 CD AD 38 00 11 EB
 8F BE 1C 08 06 69 71 49 DE BA 05 12 4B 82 28 17
 9B 51 27 A8 32 EF 42 06 D0 04 15 02 FE D6 61 D8
 52 91 52 0A 94 34 FC 90 C6 61 58 66 8F A9 8F 61
 8E 16 3F 78 30 87 93 DC 79 11 C7 F8 84 F0 A5 4B
 03 04 F3 6C B0 8D 6D A1 3C D9 17 83 D7 97 8D FA
 C5 78 3C 34 2B 9D BA 29 CD 8A D9 BB 1C FD F8 17
 91 FD BB 5A 9F CF 7B AC 7C 35 70 C5 FE 93 D5 7D
 90 BC B5 22 82 25 5A 42 1B D5 C5 9C 9F C6 80 48
 87 49 05 98 96 B8 78 95 BA F6 EA 22 12 80 80 DD
 A8 0F EA EE E0 A4 01 75 30 8A C5 AE 1C 1A F3 41
 4C EF CB 9B 28 80 D5 80 5C 5E A8 EC F1 24 60 8E
 6D 44 CC 80 F5 A9 7B FF 2A DD 7A 2C 65 E7 F8 84
 8A 66 40 E9 0E 91 39 F3 78 96 8F B2 D9 16 21 73
 6E 72 50 5E B2 B7 56 A0 63 EA 72 FB 09 8B 1C 19
 76 30 CB 0B E7 CD 5F F9 F1 B0 7C 93 E1 97 E1 0B
 4C 42 68 BB 0C 19 E2 28 74 47 0C 23 BB 8A 7E E8
 02 EC 95 EF 1C B7 D4 F5 67 D4 A5 17 E5 D6 22 9E
 E3 45 50 CD 67 81 0D DA 39 6D D5 F8 11 12 6D A1
 1E 2A 7A AC F3 83 B9 C8 5B E9 51 7C 01 FC 7E AC
 9B 6D 05 DE D2 89 1D D1 F3 2E 68 D2 36 BB 67 03
 59 79 F5 A5 3C 10 D9 03 CF EE B6 A6 43 B4 2E D6
 FC D6 0F 71 26 00 BB 52 E9 60 5D FD 21 E5 07 77
 F5 2F 28 AD 19 9F 49 9A 1E 6F 8B 3A 29 D2 85 8C
 19 1B 4B F5 97 16 9C 3B 1B 67 D2 FB B8 1E 54 5D
 32 BF F5 AA 63 C5 29 1F FF B6 23 E1 CD A3 46 24
 B0 DD 88 F7 58 ED CE 26 43 6B 7F 61 80 E9 00 F8
 94 6D 1F 73 C4 FB 17 E3 D7 DC 24 34 C9 EB EA 59
 34 10 3F 23 53 3F 6D EE 5F 28 62 D5 F3 50 C8 D7
 47 D8 3B 58 02 96 C8 89 9D 40 5B D7 CF 9C E8 D3
 F9 21 CD 14 E2 6C F4 D2 7A 4F 2A A3 BD EE D6 03
 4C 9A 94 9E FB 2F 4C 85 44 59 62 90 34 B8 C9 AF
 4C DC E6 47 51 82 90 E3 E5 E8 88 80 E4 E5 6B 56
 7B 52 6F 75 C9 2A EC 57 25 B1 5E 63 2C 90 DB 68
 AE 06 76 CD 2B B5 2C A7 97 18 9F 74 20 56 84 90
 D5 1F E6 8C C0 51 0D FA F3 F6 EE EF B6 C2 43 44
 61 DB DB 65 6C 6B D3 9C 0A 95 24 89 07 C5 F3 E1
 D8 93 4E 87 52 2F 6E BD 29 4F 32 CB E1 C9 DF 3D
 94 77 66 31 08 23 BC 63 EC 87 AF 8C 37 D1 F0 11
 1F 9D 70 DB ED B1 65 1A 04 99 E7 DB 16 E6 A0 9C
 A3 4F 97 40 65 06 D7 0F 2D 6E DD ED E6 8D 08 D9
 4A CB 98 3C D6 4B 5E 59 F3 8B B1 67 16 D6 EC 9D
 B5 B7 18 45 CF 60 6B D4 FD 36 06 72 29 46 4C C0
 04 AB DD EF BE 2F F0 E0 4D 4D AD B1 E1 C5 E9 97
 15 C9 B7 17 B7 AB C0 43 56 CC 1C 9E B3 5B B5 74
 FE E7 2B 76 1C 9A 07 A2 E0 3B 5A 1D FC 55 C4 3E
 D6 AF E4 A2 F1 FB FB 49 04 B7 09 23 EC 73 08 17
 34 1B C6 70 2F 3C 18 70 68 37 AA B0 B0 5B 4A 05
 E7 53 3E C1 FD AE F4 9E D2 26 1D FC D5 18 12 60
 12 8A 44 6F 57 1C 20 E9 CC A7 39 52 99 36 2C C6
 81 31 FE A3 A4 2C AC C2 4B 34 53 9C 53 D2 9C 44
 D5 56 2B 26 7C 75 66 50 16 68 C8 0E B0 59 23 8D
 D1 3D A4 0C 22 9D 69 77 EC 58 D6 73 7D 3F 29 43
 E3 99 AD 05 D5 02 C3 A8 D3 F3 B6 F9 21 6D 32 44
 63 B6 85 46 E4 B6 E3 6E AE 6F 3D 01 E8 06 19 16
 8C 37 A8 4D F4 8B CA F3 F4 88 A9 7C 10 84 3F 44
 3A 70 32 E2 67 2E F3 7E 33 E9 1F 18 4D 68 5B CF
 EB FC DA 61 6C 1C C3 1B 85 B4 8F 34 AB 36 21 45
 4C 70 3A 89 2A 9D 76 FB 69 C3 12 B1 37 FC 62 9B
 CB D8 77 38 AB 68 86 BB E5 F5 79 24 B6 7C 43 37
 42 0B 3D 3C 82 E6 FF D0 DB 92 E0 04 82 F0 8F 26
 18 B4 B1 AE 48 E7 42 97 F6 71 48 CA E9 5D 29 B2
 4C F4 76 53 99 C9 6B AF 28 AF F6 0A E6 B7 A0 C1
 2F 37 9E 23 E7 5D 69 EC A8 9B CD 9D 5E B8 F8 24
 DA 1C 75 75 15 CE 40 85 A8 DF 78 06 F4 FD 99 3D
 2D 58 EB 70 3F D2 C6 9A CA EC 0B BA 8F BA 2A DD
 05 E4 B0 59 91 72 4D 86 22 45 7D A5 D2 91 79 71
 34 20 B4 D9 6B A2 1A 8C 00 34 0F 72 ED 28 A8 3A
 01 46 A9 64 D0 A1 A0 72 C4 AE B2 6E 31 F3 29 F1
 7F F6 F9 56 E7 9C 89 6E 8B C3 8C 67 E0 BE 16 E8
 D8 33 0D 9C 92 F2 11 9E 1A 11 53 1B E2 49 FE 68
 11 54 12 12 6D 64 DA FA 94 1D 75 00 63 EC 7C BC
 4E 5E 2C 92 46 65 E7 58 87 5F DB EE D3 51 63 99
 EC 1B 8D BC 6F 94 65 FB D7 ED BD 78 CF 99 56 C9
 DA EE 40 A7 61 F3 E9 48 F7 80 0E AF 1D 43 FF 46
 19 AA EE EF 50 F8 35 49 C0 C4 0B EE 8E 79 8D 81
 C6 25 54 8A 90 3D 1A 60 BB 66 99 B8 4B 42 DC D2
 B5 F5 7C 05 DB 32 85 A8 3D 0B F8 2F C4 8F 4C 60
 58 29 0A EE 2F DE 04 7C 1C 0B BC 07 AF 57 5B 99
 1B 62 AE 46 18 54 12 02 E8 09 AB DC 7D B7 E7 AE
 1E 37 1E F7 56 15 B2 03 B7 E9 1F 2B FD 02 CE F6
 A8 3A 82 B7 CB AD 25 69 7A 63 EB 51 B7 49 C8 9C
 90 DE A4 61 03 2A 4E AB 1F 79 98 DB 4C 02 49 81
 D0 CE 29 66 02 36 43 10 45 F3 91 38 96 48 31 B9
 6B 7D 0D 5B CD 30 23 4A 38 72 3B 20 3B F4 FD 63
 56 0D 2F 8B C6 BA B0 AF B1 88 D2 43 DB 46 8D 84
 7C C8 13 59 88 37 A8 1C CD E5 4C A3 6B 71 93 8B
 97 41 C6 16 FF 24 2C 6E 2F AB 6A 2B ED E3 76 9B
 68 46 10 38 AD C6 F3 CD F9 2B 95 F6 75 9D 40 28
 D3 82 CA 06 1C E8 FD 60 55 3A 8B DA 13 7F 4E 61
 D8 0B F1 18 86 2A 5A 2E 64 A2 42 D4 67 B0 8B D5
 62 19 6D 01 66 7E D2 1D 67 1D C1 37 EE CA F0 18
 3C C6 D1 78 C9 2F 1C D4 19 C5 2A 6C 1C 59 AC 42
 EA D3 5C 34 76 3D CA D5 12 B4 18 C3 25 5A D7 CC
 08 E9 08 CC 10 A6 11 CF 4A 6C A1 88 EA 77 74 55
 88 E7 EC 94 D0 E2 4A 16 6B D9 DD A8 4D FB FB 2F
 34 0A 70 94 7C 84 F4 71 36 94 D5 40 6E EC 9F E9
 67 1F 86 EB A0 1C 79 F4 C3 FA CB F6 77 25 56 0B
 2E 23 53 89 C3 38 18 E4 F2 A2 85 E9 FC F7 12 57
 A4 4D A1 E3 E5 CF 4E F6 E4 9F 6F EC 6E 68 95 9E
 1B 42 DE 15 4D C5 44 B1 EA F2 E2 09 03 5C 75 FC
 96 FD EF E4 71 27 1E C5 13 AE 54 91 8F D0 44 B8
 33 4F CC 3D 2A DA E1 1E 50 0B 2E 35 BC 72 3A 65
 14 20 7F F9 65 6B B4 FA CD 83 17 59 C2 DB EE 38
 BA EF 6E B0 53 97 BB B1 1A 62 0E 13 6A AC C2 B4
 6F D3 54 3D 41 C4 20 D0 1A 61 C7 44 6D 9C 95 35
 2C 0D 7C D9 83 E2 58 41 89 26 9F BC BA 61 2B F0
 C1 E5 B9 35 45 5B 7D 5A C6 0E 8E 3C CC 19 17 9F
 E0 FE 31 75 BF 6C 51 39 C1 56 CB 11 7C BC B2 75
 A5 DC E0 4E 6D 39 66 4A B1 3F AD E6 5E 95 79 4F
 FA E1 61 A4 4D 99 8D 2D 9B 64 B4 82 A9 2D 77 2F
 7F 73 A1 DE 57 82 CE 9D 29 23 EF C2 18 74 C6 5B
 3C 8C F1 39 8D 35 C3 71 DE 3F B7 29 41 C3 7D 39
 5F 9E 1C 49 CC 4A 0C 25 F7 E2 28 01 02 50 5F CF
 87 EE 51 FB AE DD BE 8C DC CB C4 5F F5 19 19 05
 50 48 30 0F 12 F9 99 74 F5 45 13 A1 F5 39 69 7E
 F1 F8 C6 BC 0E 24 A2 0A 70 60 DE 04 D6 EC 7B B8
 42 A6 FC CD 23 AD 07 F9 3B 4B 94 BE A0 05 10 19
 75 48 4D 57 3C 3E 42 87 8F A2 C7 10 40 8D 12 3E
 54 15 AB 5A 7B 92 22 AC 68 0E 70 65 5B B4 F0 52
 ED CB 38 EC 92 1D 81 81 21 70 B3 43 DA 8D 70 24
 12 E5 DB 02 6A F7 2B 82 5B 4A 16 4B C8 D6 7D 9F
 27 14 7B FB 78 2D EB 35 3A 66 CF 7E 36 93 FA 9F
 C1 99 06 75 D6 9E 1A 2C C4 98 4F 1B 94 34 5F F2
 4C 74 1A D6 87 7A 87 CB CC 3D E5 5A AF 63 B6 4B
 B0 08 C4 37 AC 36 BC ED AC 76 29 F5 06 F0 C2 C5
 57 79 9D 24 87 20 EC 66 0D 77 CA 5C C2 F6 D9 BC
 0B 63 5C 30 4E 93 72 7F B1 95 7A D6 A2 13 F4 09
 52 09 39 1A 98 12 23 EC 22 6B BF F6 0D 09 E7 FE
 AF 34 FE DA A7 59 E5 58 CD 32 9F 53 73 34 5E D4
 A0 EC 39 A1 35 B3 66 0C CD 9A 6D 46 12 6B 1F B6
 59 8C 84 55 00 BD 16 50 8D 39 DA A2 09 08 FB DC
 B5 DC 8F B4 95 CB 6E 7A 09 B9 AE 93 31 E7 6F D3
 87 0A 61 D2 9E 0F F9 CF 81 DD 23 41 39 4A 31 81
 CA 6A CD 0F 4F 29 5F 34 35 F2 0E EF AF 4F D0 1C
 D0 A1 40 95 C8 44 52 92 24 FA 33 8F 77 63 A8 40
 D3 48 C3 B4 27 6B 88 F5 4F EC 5A 1A 64 98 A1 0E
 25 E2 82 45 27 29 2C D3 A5 49 64 C1 3D 8C 2B 72
 F9 2D 0D 09 D1 DB 55 74 B5 02 09 0A A9 2A B3 CF
 F8 63 FF 36 9C 7F 62 89 A9 BE 66 F3 73 41 34 16
 1A B0 6C F0 9D 2F 88 96 52 07 BA 06 7A 5E CB 0D
 1A E8 89 23 E0 8F C5 E9 41 EF 06 AE A8 6C 1B 58
 7E B1 F8 AC 46 04 C4 FC 22 6D CF DB 2E CE 7D 6D
 41 28 C8 90 38 C2 AF 15 D3 98 40 E4 44 D5 69 DE
 4C 0A E6 8B B8 4A EC CE 5B 85 11 8C A5 99 D8 CB
 8C F4 36 A7 D8 A1 48 A9 F9 DE 26 3A AE 54 75 19
 B6 F9 D3 6A EE 92 30 FB 02 39 B9 53 E2 E5 7B 02
 13 48 9E 1F D9 D4 7E 09 A1 B1 F0 D7 6B D8 E5 A1
 A5 36 B0 81 E2 00 1D 6F AA B7 C6 82 DE CC FC 30
 0D 12 87 9C 9A 26 4A 80 FE 16 9E 59 67 5F AD B4
 42 D1 0E 34 51 34 F7 4B C2 CB 6D E1 0E 53 7A 38
 A7 F2 FD 87 BD 19 BD 47 78 3D 1E 70 C6 5C 04 D8
 E1 FC C7 ED C6 BE F8 6B 27 DB 92 7F C7 5E E1 1F
 6B 74 99 B2 59 78 20 A4 79 CD 53 C7 51 B9 4D AC
 F0 63 B7 99 90 77 4D B9 C5 96 C9 43 CB AE 59 1F
 00 BE 6E 0E 32 A9 CB 17 C3 A6 B4 27 97 2A 8C 54
 13 7D 11 46 89 9E 7A 97 F8 A7 D9 35 B0 64 C6 01
 14 10 6B 66 BD B2 B8 85 F8 82 69 35 8C EF 5C 72
 4D 6B 81 79 34 8B 5B 3C F6 69 0F 11 61 7E 51 E7
 5D A6 BB 01 E0 48 38 82 FC 7E 39 ED E5 70 86 47
 7C C1 5A 59 9E AE 90 4E 8B 92 6D 8C B7 04 B5 1A
 EE A4 4F 7F D2 EE E0 DF 16 2F D3 2E 8B 39 A9 CF
 1E 5E BA 32 F3 F9 72 E0 7F 9D EC D3 81 80 C6 4C
 9C 31 20 26 DC 9F 28 CD B9 04 88 D9 3C 47 3F 90
 94 E0 57 F3 13 C0 92 D8 25 B5 D5 2C 39 64 3D 53
 49 9C CD 38 5B 50 3E 75 34 66 BA 4B 21 F3 DF B5
 83 A8 2F 95 D3 CB EC 83 AA A8 78 11 06 62 5A 84
 E4 09 B1 9B F8 1F 8A 64 53 2E 55 04 74 6C 2A 46
 A8 D9 FE 20 8C B4 70 13 95 A4 9D 01 2A 10 BA 9D
 67 C7 7B AC C8 34 46 3C 7E 3A 25 B5 A1 C6 5A D8
 1F B4 EE 0D 43 80 16 AA 66 74 01 35 2B EA 99 3F
 AA E7 CE AE 19 27 39 D3 80 8B 20 36 1F EF 7D D8
 ED 59 78 CA 80 87 DC EA 10 CD 89 8A A9 FE 8A D7
 85 03 05 B0 95 38 F7 8C 89 AF 48 C4 C9 ED 92 87
 5E BE 44 0F A4 C3 03 62 AA 87 BD 59 AF 16 68 11
 9F B6 CB 5F 92 41 CE A6 B9 C5 9C ED B4 D1 E8 84
 60 05 DC C8 66 BE 18 E2 4F AC EF 03 E4 71 35 86
 45 E9 90 09 42 3E E0 7B C2 5D 74 DA 50 CC 2A CD
 CF D9 8D EF 3E 9C C9 A2 60 49 68 89 E3 AC 15 95
 B2 51 FC EC C4 5C 4E 35 EB 2A 45 DE 0B 6B F0 00
 22 64 28 89 98 F1 6F D9 48 41 C8 3A B0 C4 45 1D
 91 D9 6C 28 F7 AD 9A 12 A1 DA 73 AF F4 D5 96 1D
 34 68 E3 DC E2 6C F4 F1 70 3F B9 4F 92 A7 91 07
 4D 04 5B 3F E3 43 9B C9 10 8D 47 AC 16 B9 B0 CB
 B3 85 99 F8 34 CB 82 66 44 26 8F C4 24 87 C3 0A
 DE F2 A8 F2 5A D0 7C BC 0A 03 0F D8 18 9D CA 59
 5B 28 07 2A 6F 7B B7 CD D2 D1 F5 DE 93 C0 9D F7
 3B 3E 0C 74 73 87 E2 37 AF 20 5B F9 48 0E 0E 42
 46 89 29 C5 B1 1C BA CA C7 DE 4C 59 9F E0 BB 59
 82 02 5C C0 F1 E9 89 FC 7B 9B 16 85 5E 44 9A B3
 13 83 6C 10 48 57 5E 56 6D 8C F0 B2 7F CC FB 59
 68 8E 05 EB C4 91 9B BF 55 59 F2 8A 80 AB 6B 0A
 EE C8 A3 44 C8 FE 66 39 80 AE F8 78 8D 83 15 86
 A8 A5 74 C8 DB 63 62 06 CC 1D 07 8B EB 01 33 E6
 1D DB 70 B1 3D 79 F1 26 BA C2 26 30 4A D7 27 19
 2F 15 47 7F 85 E8 56 83 19 5B DC C1 5D 10 9D 9C
 D4 20 56 A1 C4 60 22 82 A7 43 E0 69 D5 96 D2 38
 C5 83 4B A3 C7 95 D5 ED 44 86 5E 6B D0 07 A5 96
 37 85 D6 E4 E9 9F 43 2E 71 31 D2 D4 D4 C7 F8 44
 D3 F0 99 72 D2 21 5B 9E 9E CE EB 55 D4 85 17 23
 5E CA 4C 35 59 25 F4 2B A2 37 04 2D 92 46 12 3B
 2A E5 C0 35 04 58 74 BB 4E 82 7E D4 F0 70 2E ED
 E4 52 D2 09 44 DC BD 9B 44 50 89 CD 7C 61 E1 44
 4B A3 21 D3 76 86 26 FC 70 DC 03 01 D9 4C 57 47
 1F 42 29 11 52 BB 39 83 2B CC A0 AB 7D 4D 37 D4
 85 95 03 D7 F3 59 B0 16 02 E9 83 C3 B7 9F 52 44
 EE 35 7C A8 45 7E 68 4D 41 90 C8 32 76 D8 3B F3
 C6 6C 21 ED CD C7 32 DB 4D 4D 6D C4 B2 F3 87 DE
 91 98 94 85 73 A9 51 CC E8 3E 47 DA C8 1B D7 93
 A3 E8 E4 56 A4 F9 61 13 78 F9 05 52 99 98 6B 7E
 DC F2 FF 67 4C 4B 41 E9 8E 81 97 8E CB D8 A1 A9
 F2 77 A8 8E B9 AA 4A F0 3D 48 0D 50 7A 59 D2 5E
 92 68 47 0E B9 97 C0 20 7A 2C 15 22 78 51 23 F6
 24 BC 8C 03 95 D9 25 C3 EE 12 28 23 DA E7 37 DA
 B5 F1 A7 96 29 6C 43 30 B8 12 04 8A A8 21 DB 98
 5D 67 66 AF 73 F1 17 F2 F5 24 48 E9 59 BA 38 28
 E8 F7 F5 63 53 1F 54 2A 21 40 F9 2F 36 74 66 E1
 AB 8C 8E CF 76 B7 73 4B 36 27 AB 6A F5 E1 3B 97
 1C 24 2C DD EB AD FF 17 95 18 9F 7F 9B E4 AE 60
 C9 D1 5D 9C 1C 94 D9 13 57 8C 3A CC 94 C9 42 F9
 61 82 A2 F6 2B A7 0D E5 E2 7D DB F3 75 DF CB 7D
 C0 0A 5B 41 7C D5 BE C8 8B 1D FD A7 C7 FD CD 39
 4F 53 22 3D A7 E6 FB 19 A7 44 B0 B2 DD 44 2E 0A
 1F 0B B5 D1 EE CE 93 8A 59 EF 42 7E 77 57 FF 12
 83 6E 0B 3C E3 4B C4 45 C5 C2 99 A4 15 9D DB 92
 82 34 86 65 8C 5D 0C B8 4D 5C AA 49 0F 54 B7 FF
 2C D8 6B C6 94 75 52 A1 61 69 D5 0A 60 AA 29 BC
 49 4D 29 0E A1 E4 E8 6F 97 9A B3 D9 11 05 68 94
 8E 29 54 A2 1E 80 C2 C3 9F 1E 79 29 61 39 66 50
 73 9E 2E 3F 7A CE 76 9B C1 01 74 8F 76 82 A6 37
 B0 EB 86 3E D6 EE B0 4C 4D 07 D4 F7 99 17 BE 49
 66 EE D2 AD 6D 31 8A CB B0 6B 5E E5 D7 BF AC 07
 0D AA B2 D8 50 FA 90 B5 C3 F4 1C E8 92 51 0B 4A
 46 89 55 32 5C FC AF FA 57 76 00 DD AB A5 5F FC
 18 0E F6 54 CE 11 4E 9E E7 67 85 53 B9 C5 76 DC
 B5 00 C7 92 B6 42 15 E5 99 35 EB 5A 04 DA 01 87
 8A 73 E5 39 5C 77 FE B8 72 92 F4 C8 E2 49 E5 23
 C0 10 40 72 FD 80 8C D6 BC E7 DA 85 1B 34 AC D5
 F9 DD 3C 09 29 D7 3B FD 27 72 69 6F 25 2F 7F ED
 AB 22 75 1C CE B3 A7 DE 57 62 E1 6B C3 A7 64 44
 74 5F F4 BD 1F C8 49 5A 3E 1D F5 B9 5D D8 5B 2A
 71 6F B4 DE 89 10 00 A2 0E B6 68 71 7D E3 31 C1
 4D AD 66 A8 C0 1A E2 57 BC E0 23 79 48 A5 43 AF
 A4 10 D5 3D 99 E0 9C 24 F3 7C 9C 05 3B 31 C9 A6
 E5 2B 09 7A 7C 85 B5 EC 56 3D F5 36 98 9F FE DD
 E9 69 94 F1 35 08 A7 70 92 32 CE D1 92 E9 B7 DE
 FC A6 FE 08 63 CD F3 E6 01 D9 F5 61 CD B0 8F D9
 85 2F 39 91 40 F1 27 E8 37 E1 19 0B B2 AB EA B4
 CF DA 90 FD D1 23 60 E0 0D C5 00 B0 2E C7 E9 50
 02 80 84 F3 76 36 E1 E6 9A C9 8D B6 20 E4 20 61
 43 A3 17 46 40 48 D0 A4 47 3F 2B 7D 7A 0C 5F 7C
 9B 29 17 DE 33 50 41 F1 96 8D A6 16 56 A5 E2 EE
 CF C6 98 28 38 60 BB 0B FD 6E 97 A7 92 96 31 60
 66 84 55 A2 CB AB 00 D3 49 2D C3 25 57 97 3B 3B
 AD 27 35 8B BD 15 99 9C 83 FA BF 85 6C A6 A0 FD
 47 51 93 64 AC 5D 48 7B 0B 07 35 7A 22 05 4C 5D
 C4 14 A9 05 6A B2 B0 07 D9 CC 7C 25 6B F0 54 83
 DC 8D BD 1B FB C2 D0 0A 27 79 E7 DE 16 C7 84 8D
 F8 48 D2 27 FB D7 54 4C A9 B4 4B CE 93 B6 C2 8A
 6F BD BE F3 08 03 CB 81 EE 91 3C 6F CC 4F E1 AD
 31 C1 00 70 AC 24 E8 1E F7 FD 7A 3C 99 9A 51 4B
 5A 48 3A CD EE 80 FD ED 59 19 13 52 CC 7F 73 1F
 B6 60 8F B0 B5 65 F2 1F 7E 18 DB 82 40 0A 9A 3B
 7A B7 7A 00 22 3F 63 63 DC 83 B0 C0 D2 03 AE 6F
 79 5C EC FD 6A ED 26 27 FE D1 D5 0A 3F 30 F1 8F
 7D 49 AF B8 AC 49 81 81 2E 17 E3 BB 1E 3C 46 1F
 41 8B 80 80 E4 51 C1 BA 54 12 67 76 67 87 50 D9
 B5 10 D4 A3 CE 84 FD 57 55 AB AF 5E B0 57 E7 FC
 98 2F A0 26 00 D1 50 43 C2 42 7C E1 47 A4 49 CE
 7E 35 B4 AA 66 81 5B AC 3A 77 03 72 EC FF 06 53
 6D 55 4C 77 59 BF 5D 0F 21 EB 30 19 DC A4 00 96
 61 46 6D B0 C1 47 2D C5 3F 1D 09 7F 0C 88 D0 F3
 FC 33 31 A9 01 4D 79 03 A8 A0 C5 AC AA 1B E5 7B
 3A 36 E4 07 8D B9 12 AE 9B 0B DC 31 6D 1A CC A6
 49 A2 80 64 68 07 9E E4 F3 4E E4 8C 45 B2 FC 55
 DB 5E 3D A5 EE 45 53 52 BE E6 9A 8E 12 99 9B 06
 F4 98 46 D8 2A 7D C6 11 AB 25 FA D2 6E CE FB D8
 C9 86 DB 30 21 05 FE E5 21 93 DC 4A 3D 4D 28 F2
 91 F0 4A F7 61 15 F4 26 5D 9B 76 0E C3 3C BA 8A
 77 89 F8 A0 53 DB C3 4D 55 28 48 D0 72 3A 19 0A
 AB DF 8A 56 9A 5A 97 0A 53 BA 68 A8 C9 E6 2A 07
 E2 BA C8 D6 D6 61 97 03 20 34 CF 8E 92 59 1E 3C
 9A 95 EC 4E 6D 54 FA E1 C1 92 D8 4A 3B 59 17 8A
 88 9E CC B0 F2 F3 8A 00 FB CA B2 FF 42 63 22 AA
 9F A8 C3 A1 01 A1 60 C6 3A 25 B8 B1 5E 90 80 3E
 09 CB 6B 43 62 F2 22 AF 3D 43 7A 44 C6 2A F6 45
 A9 95 AC 41 03 B2 7D 69 69 CC 29 B4 F8 1D 9F 3B
 7F A6 86 8F 16 1D E0 4D F0 B3 18 AE 67 1C EB E1
 84 A8 D6 0B 46 47 02 AF 8A 01 8C 42 31 78 D1 63
 ED 92 54 40 57 AC A5 36 A4 92 D4 B8 F2 0F 2D 4A
 B2 DD 5E C9 AB 90 99 E0 6F FB D0 29 13 46 33 CA
 9C 26 03 F0 80 6C 11 48 58 82 AA 6A 53 0A AD 05
 8D 32 FA C1 9B 5F E5 2A 9C 9D 08 AC D3 17 A8 F8
 5F 23 1B 67 FB 98 B8 54 AB FF 83 87 A1 BB C2 CD
 43 B3 BD 7E 85 9E F1 FA 8A 5C CB 4C 6B 30 88 DD
 6B 9E E5 07 1C EB 8A 57 64 1B 51 F7 30 54 4E 67
 3D 5C 1C 44 29 15 93 B3 46 7E 79 58 8B 6A 03 AA
 32 43 28 A0 59 3B 13 1E 64 1D 42 9F 73 47 E1 A8
 0D 1A 3C 7B 80 6A BA CB 93 A7 78 85 5C F9 0C 5A
 E5 D9 E0 AB 28 07 DA E2 BA 77 39 E0 D0 A1 89 F0
 AD 09 1F 91 37 4C 01 A7 C6 D2 45 93 32 08 DA B9
 4A 1F 64 C9 A6 2F 0B B9 CD 95 C8 99 CB 7D 0A EC
 26 D9 F8 62 08 E6 26 D3 6B F6 20 06 36 D1 00 E0
 39 FA 76 42 6C 3E FE 3C 66 3E 78 24 11 90 A6 C7
 82 05 F7 C5 65 B5 B7 74 00 B4 85 B8 C1 0A B8 D7
 27 DE 5D 93 C2 A6 30 0A D4 F1 40 3E 8F 1F 34 48
 03 C0 D2 2B 05 D0 22 E7 99 68 8C 17 95 21 CF BB
 40 3E 76 06 01 ED B2 F8 15 BE 96 0B ED 8B 71 FB
 34 58 3B C0 FA 84 77 9A 65 F2 60 CD 97 29 34 1B
 F8 F1 5D E0 19 32 24 D1 CC 06 96 4C 4B B7 BC 8C
 30 0F 36 36 58 00 88 05 1E 5D 94 BD AC F3 36 18
 84 55 15 EB D6 70 E2 C7 AF E3 05 D1 7B 6F CE 5B
 8A D7 88 F7 0A C9 B8 7A DD 2A C2 36 5A E7 CB 4A
 AC 50 CD 29 4B 51 AE D8 5B FC 7C B6 E3 BC 63 23
 8D B7 E5 1F 67 76 A1 71 47 E3 64 DC 91 3B 83 4E
 41 95 D5 45 24 12 A6 1B A3 DB A3 23 0C 5E B3 AD
 E6 62 A6 50 28 DA 0C E5 9D 41 8D 8D FA DD 98 BC
 6C 68 60 DD 48 BD 55 F7 32 A5 3E 6A 03 59 8A 2E
 83 AC 01 54 CB 8F C7 CF DD 7C FB CD C3 4E DB 8F
 AF 68 33 30 9D 73 9B D5 24 97 47 91 60 B9 DF F7
 44 B4 6C 0A FF 3F 04 EA 24 CF 89 54 48 00 AB CE
 C9 8E 6B E2 8B DB 1F 3B CB BB 09 E7 E3 29 A3 B4
 C1 A3 05 04 42 AC 5F 5A 1B 26 97 7A 87 89 53 A8
 D2 AD 6E 57 E4 FE 9C 81 1B 41 50 95 E0 19 DC D0
 B1 CF 02 F1 03 AF 5D 10 37 6E B6 09 74 3D 74 F9
 5F 08 8C 4E 77 04 F4 2E 4D 1E 79 6D AA 1D FA 81
 D3 06 EC 4D 85 12 DE 21 8B 79 4B 16 AB 78 47 61
 1D 63 14 F9 FC 44 AF B0 BD 04 FB C6 54 EB F0 C2
 A2 21 8F 80 FD 85 F3 C7 21 04 B5 72 E2 B2 EC 4D
 67 44 D8 C4 69 7B 79 50 2E 21 2A 3D 75 20 31 71
 E6 C8 2F 0A 16 E4 7D FA D0 05 3D F6 F9 25 CC 04
 1C 69 30 AF EE 4E 5F 45 64 78 66 1D DD D0 12 2F
 BB AA 99 84 84 A5 92 E3 0B FE E2 0E 9C 94 EF D3
 19 39 CA 6A A5 14 E3 D3 8A A3 B4 B1 73 66 60 DB
 AB 5C 5C 70 F5 BC 71 DC 3D BD 70 5A B4 ED F6 CD
 5D AE 6D 8D A5 53 9B BF D6 E7 E6 5E 0A 70 93 0A
 75 E4 92 12 FF A5 CA 34 5E 29 D3 22 47 9E 30 17
 ED E6 66 27 20 6B 2B 33 44 56 F6 91 D6 4A 47 F0
 90 08 6A 64 3D 73 CE 3B 94 D8 67 05 80 BF 39 BE
 A4 FD 5D FA 5F 4D BB 8A 2C E3 9A 5B 4C 8D BC 88
 2D A8 4C 23 A4 8D D9 43 5F 48 D0 1A 28 27 A3 FC
 2F 4F 78 00 F6 90 77 85 35 59 8E 5A 08 62 C6 17
 D3 71 E6 4F A5 C6 37 E2 3B CE 90 D2 7B CC 9D 38
 9B 44 D7 05 ED ED 7D 50 B3 61 27 FF 72 23 00 D3
 C4 6A 50 BA B3 5E 12 DA 84 D7 3C 54 F2 C6 CA 41
 13 6E F5 AD 0E 4C F6 55 AA 00 A1 67 0A 38 16 E8
 34 54 1D 5F C7 F7 6F 1D E7 2B 7E A1 65 48 A9 EB
 89 F2 90 B8 50 33 FC C1 FD A0 32 FA 20 FE 86 A0
 41 3D ED 01 56 C0 27 4E 4F 93 63 E9 F4 49 92 D6
 E3 40 0E 6E 05 D1 B2 59 71 51 16 18 80 B6 F1 52
 04 03 50 12 82 45 70 8E A4 16 ED 12 63 FD 7D 60
 06 4C DA 4A 8B CA 13 F4 DF B3 94 8E 09 D2 93 D5
 52 22 FA 09 98 09 22 D6 1B 56 EB 49 7D 0A BC EB
 FB FB DB B4 ED F4 A9 D5 FA F6 30 4B 18 D2 12 A2
 A0 A8 EB 8B 4F F2 12 E3 7E CA 05 3E AC C8 45 99
 21 3B E2 57 DA 12 B9 5D B2 DB AA 53 99 40 E2 E8
 E9 CF B5 9A B1 3D 90 33 BF DD CF 85 4B 65 7D 7A
 8A E2 EC 8D 75 3F BB 19 03 76 80 A8 A2 69 9E C9
 5D 46 26 33 F6 20 87 28 AC A2 72 98 4B 78 58 FE
 A1 EF C6 FE FE ED 99 69 14 52 47 D1 23 63 07 61
 DB 54 BD 23 95 37 79 6C 2B DF CC 4A AA 62 B2 57
 0A B6 53 CD F2 C2 9F 3F 5C 11 78 F1 DE 14 19 44
 B4 3B 15 AC 7B E1 74 92 4F 84 65 CA EA 53 44 85
 09 EF 10 A5 4A 53 8F E2 C1 F2 06 D0 5D 20 AC 7B
 3F 4F 36 28 A6 1B 8F 2C F9 F0 05 11 54 5C 20 FC
 84 96 7C 19 13 ED 39 8A D0 4B AF ED 1B C6 1F B2
 95 27 6C 50 D6 F9 FD 13 50 92 42 BC 74 72 4E 0E
 03 67 F6 4E 4B 5E 14 40 59 92 58 BE 6F 39 E1 93
 56 B6 54 B4 37 9C C3 54 47 E9 7F D8 D8 78 31 26
 E1 D0 7C AF 4F 3C 06 3B CF 00 2A E3 A7 47 4B 2A
 4D CA 86 EF AC B7 BF 1D 2C 5E 2C 47 2D E6 CF CC
 FC 86 34 55 84 A6 D8 F4 53 BC 42 4E A0 89 9A 86
 18 B9 14 A7 18 CC 3E 4A C8 95 48 F6 3F 27 DB 40
 41 BA C4 CD 9E 13 D5 E1 92 80 96 84 24 22 F9 40
 34 CC 2E BB DA 5E 8D 37 E5 CB 1C C3 E6 C9 7C FE
 6E A2 51 3F 2F FF 14 8D 87 E2 99 08 33 D2 C4 68
 45 AE 7F 0A 27 2B B3 07 AB 31 E3 C9 E7 4A C9 32
 F6 5C A5 8C 0E 05 08 05 2B 11 C5 40 E6 30 72 E0
 96 0A ED E7 58 34 9C A7 69 04 00 29 D3 22 24 C3
 47 25 C1 A1 9C A5 99 07 C4 E6 85 E5 DC 14 CF 73
 5C 6D ED 84 1F BC AC 5D 71 95 18 3B 73 79 0A 66
 EB 94 57 65 92 E0 EA 6F 26 C8 0D 4A EC 68 FF 09
 B0 3C DB EB F9 0A 31 06 63 C1 20 21 B0 C9 91 89
 BB 7A 74 B8 5E FA EC E2 EE BA EA EB 07 5D 5F 1C
 71 C8 1C D0 DC A3 92 C9 2F B1 20 90 35 64 0F BE
 4D 92 6D 3C EF 24 F9 99 7D 5D 53 76 F8 E7 8D B4
 0C BA 0B 54 A3 91 CE 3B F2 4D 75 87 F5 96 74 5A
 C9 A5 4C 2B DE A0 CF 34 81 EB 2F F7 86 A7 64 29
 C6 0B B3 0D EE D1 0C 94 60 DE 7B 0D 54 26 DC 42
 B3 B7 A2 52 28 32 71 3A 19 82 1B 38 69 FA DE 30
 79 EF 27 48 05 32 7B 97 80 20 9B 7F D9 97 FF 28
 DA 4B F5 CF 07 E7 F7 6B ED D5 42 9A A8 78 55 C9
 20 5A FD D6 AA 83 55 A4 80 94 0B 7A 63 56 06 F3
 C6 0B 75 B1 EF B5 62 82 83 34 65 AD 3A 9E EB 3C
 1E 85 78 1C 1C 0F C6 A0 4B AB 82 47 63 52 01 3F
 0C 87 62 8F AB 1D E3 69 67 28 78 79 95 B0 A1 3C
 73 FE 8C 78 DB B8 17 77 14 B5 16 4E 9B B3 FC D3
 1E 28 3E 7C 29 4F 39 84 68 0D E7 78 0D 42 64 24
 07 6D 4F 44 E6 99 AD 67 76 10 88 74 2D 6A 51 92
 1D BF 46 AF C2 A8 F8 44 C7 03 48 F4 1E E3 15 8E
 80 4D 79 8B FF 3E 70 58 3F 8C D2 F5 BF ED 83 8F
 38 41 6A 41 E6 D0 22 D5 87 E5 DF 42 EE 00 A5 51
 30 E8 1C B6 5F 4B B7 5E 93 53 D2 CC 4E 3B EB 12
 EE 3C C2 56 CE 96 67 2C B7 CB 77 47 4B 5B 5F C8
 C0 FD 62 15 11 3E F5 50 84 DC E3 F6 7F 34 B7 DC
 A2 F4 9D D0 06 47 DD 60 59 33 E7 CC 48 D0 C3 8C
 C8 28 33 D0 AF 4D 2B 27 39 D4 48 2B 76 9A 28 01
 E8 B0 7E 84 54 9A B6 C4 B4 4A F9 52 1A 68 D1 64
 20 DC 83 63 8F 3C 1D 8D 5A B8 59 DD D2 2E 03 04
 26 FF A6 E3 C7 F7 C5 6F 0F 5C 30 8C E8 15 24 4E
 D8 C3 F4 7D 29 75 67 18 76 44 70 B4 EC 5C 49 09
 65 04 3A 1E ED 95 D8 AB B4 E2 3E 76 1A B5 07 8D
 7A DD 3B D2 4F FD 02 D1 7A 26 16 4F 84 94 E7 CE
 E5 9F DB 64 13 53 2F 81 7D 37 7E FC 04 73 E4 B7
 DD 66 98 97 23 54 DD B9 90 FA 23 3C 6E BC 10 9C
 1F 1F B4 0A E4 08 82 A7 4A 8C 49 EC 0E B2 30 44
 FC 61 CB 6D 12 FB EC 5B 47 01 E3 31 53 67 58 81
 CA B1 90 38 E4 7E 67 C0 BC 12 D9 9F 92 A8 3B E4
 63 A4 0A 42 83 6C 3A 09 BD C7 7D 79 B2 66 43 A0
 BE B0 52 6E 98 3B C3 00 1A 75 A5 85 93 3E FF 9C
 2E 4A 6D 79 3E 62 8B ED FE FB 81 F2 F6 46 B3 14
 22 B8 E9 5D CB F4 18 EB 03 D0 82 69 33 3F 25 27
 48 04 2F 92 FD 47 04 10 3B E9 95 A8 E6 8A 17 1B
 86 BD 2D 5E 19 01 1C 60 FF 5B 6A 08 BE 8F C8 59
 2E 9D DF B4 62 5C 4B E4 48 8A DF 22 F6 C1 2D 24
 CF 82 30 45 A7 DB B4 6B 2F 1E 8D B9 72 38 26 B3
 7C EF CD 19 C4 13 99 0C FD DF CA D1 3C D7 23 6B
 24 AF D5 D8 FB DD B7 4F 13 18 25 D1 54 90 88 69
 E9 63 61 73 CB FD 5E 11 F6 F8 67 03 13 80 3C F0
 59 03 00 39 57 38 BA A0 68 DB D5 1A F4 E9 CD 07
 CB 95 97 28 80 96 85 DA DB 14 A5 5B A2 02 E5 AB
 1B FD 31 15 E7 A4 FA 86 4C 84 51 B5 6F D8 5E 94
 F6 4E 04 23 0B 2B 78 6B 76 A8 1D 43 52 F0 BE F4
 87 55 C5 21 34 E5 CE DA 69 83 2E 1D 24 ED 00 F7
 1A 49 1C 80 91 84 6B 62 AD FF 51 09 13 0E 05 75
 62 58 29 CC 35 D9 A2 7C 93 5B 93 DB 81 38 E6 D3
 57 8C E7 57 9A D0 A7 CC 84 27 74 47 D8 0C CD 0A
 B9 4F 91 89 9C 99 F3 90 D7 6F 3E 7B 73 83 53 60
 45 AB CA 2C BC 8D 8E 04 92 61 35 D6 5B B7 A3 6D
 2F 9C 33 D4 43 6A 74 D5 A1 C0 8E 43 49 2B 46 D3
 20 06 FC 38 6A 84 41 9E F8 AF 42 90 1A 32 22 1A
 55 AC 70 93 67 88 94 21 80 82 40 FE DF 07 81 33
 5F 10 C8 48 AA F7 0C 15 2F B1 C6 A1 42 87 6F 07
 F0 81 8B AD 32 D6 40 FB BC 1D AB 6A 37 73 98 D6
 94 E3 6A BF 58 74 41 8C 4B 3C 0D 3C 6E E9 B0 01
 1B 7A 5C 4C 30 B1 F4 F2 B9 D3 C3 ED A8 3D 86 18
 DA 77 5B F8 22 71 0C CF 5C 73 0F C6 F8 9A C2 5C
 E2 9E 0C 95 0C 0F CE D4 13 53 4E F6 97 5C 5A 91
 37 78 40 6F 63 5D BF 53 39 CD 3B B6 35 7E 81 F2
 58 97 3C 9D 4F 63 AE 46 3C 48 18 91 7E 43 51 73
 6C 35 1A A8 DE 8C 75 84 8F C3 87 B7 FA 03 19 AF
 9F 48 32 33 85 64 0D 0B B6 23 46 9F E5 5A 32 6F
 C1 F4 08 DB 54 27 63 57 BA D8 5E 2F 27 F1 B4 EE
 61 A5 F6 79 BF A1 89 07 B0 94 CE 82 62 FB 9A CF
 3F 95 0B 19 50 A9 95 31 6C 9D A2 BB A1 2B 0D A0
 CD 90 D6 82 28 AF 72 B7 20 0B 4D 9B 3A DB 72 97
 E1 FE C3 1D 27 16 7E 08 DC 5D 4B D0 B1 02 ED 78
 4D A6 73 7C 20 AC E7 8F 4C 8E F6 A4 7D 57 20 4F
 8D 3F 6C 22 CB B2 58 58 85 AD 18 1C A8 23 FD F8
 87 3F 69 85 93 5A B4 81 84 4D FE 01 FB 8A 09 7F
 F8 2A F6 E3 A5 A9 E0 7D 53 98 EE 99 FC 15 4E B1
 A6 81 DB 8D E6 EB 4D 3B F6 59 ED 38 30 B9 11 F0
 E4 B1 4B 7D 29 4D 64 0E 93 7B BE E8 E4 2F C4 6D
 AB 0D 85 18 19 00 F1 0B AC 73 AC 40 41 E2 D3 44
 8F 75 4A 60 D0 C5 01 60 61 96 61 AA DE EA 60 F1
 8C 95 88 CB C5 74 00 F8 6C 9F 4C 1F 44 F0 C6 BA
 26 93 DE DC 29 6E 5E 6A 89 11 F9 C8 2F 4E 91 A6
 A8 80 28 C0 6D 40 4A 77 F4 32 18 F9 6C C8 E1 50
 63 6C 93 43 FB 1E A4 93 8C 5E 43 54 FC 2D 70 3C
 5F F5 41 79 15 A5 8D E1 CE AE 5B 3E 32 EE 94 5B
 C2 EA A1 B1 CC 28 4F 11 8B 5F 9F E1 07 52 23 71
 3E 4E 45 6E 27 E3 90 65 81 5E 72 3E F7 9C A9 E6
 DF 3F 5D 67 E6 D6 D3 AE 94 24 59 6B 61 F3 31 E5
 F0 6D 13 53 E8 4C 4E 9D E8 FC 26 76 B0 9D 5F FB
 F7 51 5A 2B BC A4 90 87 F4 4C CD 96 1B 40 7D BF
 AB 98 57 6C 4A 82 61 DB BE 4E B2 29 20 EE 0D 03
 C4 5E 4B C0 BD 64 1E 4C 4B 9E 92 02 BD 0B 2E D4
 04 CE 43 E6 01 44 CE 06 FF E1 96 0B 87 E7 ED 54
 E6 47 56 C8 DB 62 17 12 C8 73 02 3E 08 00 C8 DA
 84 D3 D7 F5 EE 61 5D F2 F9 58 39 D4 53 AE 20 B7
 FB 0B 20 78 32 C8 44 1E DD 37 94 6A 6A 17 57 F4
 A7 D5 4D 11 D3 9A E2 AF 3C F7 8D F7 68 E5 E6 19
 B4 79 51 52 10 B7 C4 5F 26 B4 42 40 64 CA 1E 3F
 DD F4 58 33 DB 19 72 6E 20 5B F1 50 EB C7 A7 8C
 D5 AE CC B3 F2 91 25 54 D8 A8 45 5A C4 09 58 34
 CF 30 36 2C CE 9D 3A CE F8 33 3A F9 FD 4F F8 87
 1D 2E C2 57 07 62 1F 2F 96 5F D9 7F 1F 14 17 E7
 E9 71 85 A5 9B 12 7C FA 47 41 25 04 88 C1 A1 8C
 F3 BC 6F D6 7C 06 35 26 4F 79 48 31 82 F7 3B 2E
 29 A0 A4 E7 01 1F E2 BF 31 8A 40 D2 F9 8E 32 A1
 EE 4C E3 FD E7 AC 00 5F FF E2 CC 67 3F 5A 4D EB
 98 AD 0E 28 35 2D 1C AA 89 21 4A 8A D2 2A E5 AA
 50 17 61 83 65 0D 23 62 34 92 04 06 0A 29 3C 90
 F2 41 C3 9F 60 3F DE 68 CB 40 6E 89 E3 90 BB 52
 4A 4F 0C 15 AC 04 59 49 5C 91 FE 2A F1 AC 49 0E
 24 F3 E0 18 86 A0 C6 6F 81 14 8A 50 60 EE B6 E9
 6D 0F 31 D1 7C 55 BC 4A 1D 30 D6 CD 69 29 D4 64
 05 55 C3 3E 4D D5 EF 51 D0 2C 85 57 5C 68 54 16
 71 5E 84 C9 CB E4 30 36 0E CB 6C 38 FC 87 E9 24
 66 15 12 BE EE 36 79 79 25 83 15 A6 7D F4 CE 6A
 87 3C 4B E5 7D DD B3 AA 41 8A 06 07 27 A5 FF F4
 50 87 01 3D FE 8B AC C7 C2 CB 21 E1 BC 2D FC 30
 B5 07 9C 69 81 0B B6 A0 1A 66 23 6F 68 75 01 58
 09 30 FC EB E6 D4 29 AF D6 4F C4 09 4C 8C 8A 09
 94 8D 7A 40 03 50 0D 4A 93 09 72 F2 10 BE A6 66
 A9 F1 A5 25 A3 A0 86 43 12 2A E4 0B 71 81 E7 1A
 29 DC 5D 23 C0 0B AD A2 12 F1 A8 46 E7 DD 78 B7
 F0 B5 8F 76 03 D4 C7 C2 4C C4 3D 08 D1 77 55 6B
 DA 40 78 A0 A0 C9 01 AD 2C 85 D5 AD 2F AE 82 48
 B9 2B E3 73 90 BB A3 83 B6 34 38 54 28 F0 7F 22
 53 91 AF 64 EB 90 DE FF 8D FA 6E 06 BD 04 26 2F
 FF 19 1A 91 8C B5 44 E5 96 6C 05 20 40 55 AA BB
 9A F4 09 B0 73 D9 CE D7 97 46 82 EF 06 5C 1F E4
 F6 7F 02 F6 D5 81 1A 04 80 8E FB 04 CB 00 BB 64
 BC 7E 4A CB 74 53 6E 0F 18 E8 A0 2E D0 8A 98 40
 4C 5F 00 72 35 98 70 37 A6 25 CD 77 DE 99 12 E8
 74 86 E0 CD 18 06 08 95 F4 1E 47 00 4B 31 A1 85
 A8 BE 92 35 38 98 66 D7 1C 17 8D 0B FB 89 D5 C2
 02 BC 37 8F 14 B0 02 49 D3 A5 DB 9F 77 FB 60 87
 FC D7 94 87 30 59 98 11 16 05 AB 68 33 A7 D5 B8
 BA AD E9 A6 47 A3 93 27 35 8E 44 C0 64 35 48 68
 CE 93 74 F4 BE 5C DD 4C 3B 32 8B E1 78 E4 1E A6
 65 55 1B F8 31 B9 F0 54 5F CA E3 53 97 EB C9 58
 6E 5D 28 A2 EA 93 32 15 77 F1 49 DE 14 72 AA FE
 85 78 29 91 12 C8 66 71 7A 22 75 D3 60 50 EA 61
 43 4E 03 EA 2E EA CA 27 96 ED 25 8E A3 2B 5F 16
 D7 29 54 B6 1F 68 5A BC 32 91 CD F8 61 36 72 92
 5F B1 A3 49 29 32 DD 84 A8 62 92 A6 A2 CF DB 4A
 6B 71 6E 33 99 68 35 D4 FC E6 25 FB 72 B2 CF 1F
 03 E1 28 11 68 90 25 E9 9E A6 C8 ED 47 15 14 B6
 C9 AF FF CE 76 4C 5E 25 C3 92 FB C9 3A 39 D4 EE
 E4 BA 39 FD CF FA 8E 17 42 79 D3 1B 10 09 FF 3A
 56 59 E1 FF 18 26 27 23 AB 61 F1 B7 76 90 87 D8
 EB D9 E0 77 55 9E 2A 06 D7 FE 6B E0 C0 84 E2 27
 92 24 67 34 B4 6B B0 0C 15 78 01 44 EF 8A 68 82
 DC 65 47 AA 08 13 EB 9B 8A 86 65 6D 92 56 1E 14
 96 F9 BB 75 91 D6 DF 36 18 DD C7 F0 B8 E0 8B 3E
 96 48 2D 02 5C 75 3E 53 02 4D F7 A5 7C E2 35 76
 F0 62 9C 90 08 06 DD 4A EF EB 0A C2 02 9C E9 32
 41 92 71 44 B3 12 C4 C2 D1 16 9F 0D FC FE 77 E4
 0E 07 31 D0 D3 80 F5 35 C6 93 DB 93 6C CA AF A3
 3B 6F FA F6 FE B4 B6 EC F2 F5 98 5F BE 21 8F C1
 7C 80 F7 86 B1 66 DD 9D CA 4C 98 1A 91 4A 71 39
 89 9F 3F 16 6B 67 8A C2 58 6E 44 4A D4 C8 52 58
 52 0C 62 4F 0D 1F B7 13 4C 04 EB 49 A2 8E F2 AD
 93 B9 58 EB C6 44 29 E9 CD 9A BF F3 54 3D D4 3A
 5D A6 C6 84 6E 82 96 40 C6 00 BA 84 EE 71 0A 0B
 72 D0 D0 04 36 82 E5 9A DF 11 5A 1A B8 70 77 1D
 07 E7 B7 8E B0 F5 56 2C 04 67 23 15 7A 82 59 A7
 F3 3A 60 52 C8 8A 8D 00 32 51 F5 C6 D7 59 81 72
 C2 2D 6F B5 8E 4C E0 C7 EA 5E 9C 35 13 AA 61 F2
 54 74 09 46 FB 67 83 BC A3 C2 E3 32 AC FB DB 8A
 ED 88 63 DB 96 83 2E BF 16 34 39 FB 7B 71 97 FE
 D8 25 D3 54 58 A2 D6 B1 23 33 47 2E F6 5B E1 A5
 EA 98 00 7E F4 3B 56 37 84 AC CC 24 A0 B1 95 CF
 EC 54 B6 C6 EC 26 3A 06 A2 29 E3 C4 7B FB 59 33
 29 90 77 66 9E C7 42 BE 36 51 C3 99 71 AE 2F C9
 91 2D 74 1B 2D F6 FD E8 B7 A9 FC 58 1B AD C6 49
 D7 22 FB 6E 0B 57 C0 4C 3C 3B FC 9A 05 2D A5 0F
 50 7A 4D 2C 2B 7B 24 BE 96 3F 00 06 DE 6E 75 A6
 B8 4C B9 7A 84 D5 93 43 A8 E9 41 26 E5 AE 9D 40
 09 82 8D DE 41 F8 DC C0 6D 04 48 68 B4 F5 67 EC
 4B 64 08 C4 C1 7A 76 78 EA 34 36 09 38 28 16 46
 07 7B 66 91 3D 42 79 BC 37 86 E3 D0 22 29 8E A7
 5F 22 50 4B C3 D8 14 A0 8B 4F 3D 31 95 EB 98 C9
 32 A6 A5 76 1A 0E 74 85 86 4F 19 D1 EF 63 E6 2A
 DA DC A1 F3 42 20 09 DB 58 39 4F CA 25 62 7F 79
 DC 6F 6F 9C 22 79 53 56 F7 C9 E8 62 61 CD E3 8E
 46 3A 03 CF BF 58 8F B0 73 DD E4 16 67 A0 5B 83
 91 7D 74 5D 16 D9 57 A9 6E FD 90 36 52 4E 6C 25
 27 DA F4 DB F4 2D 4F C4 63 63 C0 A8 C8 11 42 36
 D7 A5 70 72 C3 82 89 87 66 4B 7E 3D C2 CF D1 AD
 EC 1C 0F C7 F5 22 71 C5 64 C5 4F 09 3D 54 C8 5C
 62 6B D0 38 DF E5 41 DA 62 12 49 88 67 37 44 D7
 4B 8C 55 55 EA 4B 11 AD 3E 39 1F 6D 10 CB B8 DB
 56 36 8E 10 77 A4 72 EC 07 42 D3 7D A1 13 F4 86
 E3 9C AD 6F 84 24 BB 9A 4B 1D F6 8E 92 E1 96 C9
 C6 D3 3B 0E F2 E8 BC 4D 1D F5 A6 61 4A DE 7D B8
 1A 15 D4 00 FC FD 30 24 D1 50 EE EE 99 93 A0 65
 EB 78 93 F7 F6 83 D5 BF 4A 69 67 17 61 08 61 A3
 F0 BF 85 2F 4C F8 60 D1 D6 4C 67 90 C5 B0 90 A3
 B8 77 F6 1D 93 43 10 0C 37 AE F4 DB 25 44 7B 7E
 76 6A 1F E1 30 FC 7D 1F EF 96 13 C7 51 95 4F ED
 0B E0 03 39 F7 57 9E 0D FA 36 08 7E F3 10 39 D0
 24 AC 23 32 C4 DE 6B 98 E9 85 87 D0 DA 76 0A 6E
 3D 76 B9 56 AD 4B BE F7 D1 85 FD 15 13 CE 37 E8
 53 3D DF ED 1D 18 90 52 FC 73 F4 C4 98 AD 55 BA
 87 71 84 1D 77 18 F6 9C 36 45 93 78 A5 5E DE DB
 EC DD 9C DE 4E 5E 74 FC 0E 42 2E EF C3 F3 9F 84
 41 EC 5F 6B B1 13 3E F1 B0 79 46 07 53 B3 11 B3
 F7 F0 B9 ED 65 8E DC BF 6F E9 73 C0 E1 E1 16 58
 68 9E E8 10 F6 BB 52 CF E8 DA 13 CE 69 76 2D 02
 3D E0 20 54 EA 74 91 F7 B9 6A 69 DF 06 23 4C 7D
 11 F7 EC 03 56 F3 AD 64 97 7C E7 05 D1 65 E1 2B
 09 9B 11 76 41 D7 10 66 F6 39 61 A5 5D 58 71 CB
 2A 0C 0D 97 6D 27 BB 26 FB 84 14 26 42 2A 98 9C
 A0 F7 C6 B1 15 14 FC BD 85 FA 9A 1E 30 A7 DD D6
 3B 78 70 BF 14 CB D5 01 B0 3C 9E 9B 9E 6B AD 2E
 B8 61 78 15 26 73 83 A8 E2 A3 6B 33 C4 AA 54 AD
 6D FD 99 FF 32 38 7C D3 CA FA 59 5C A4 4E 8B 5C
 E4 D1 EF BC DF 2C AF 23 AE 05 2F 36 93 65 82 04
 9D B5 15 AD D2 49 5F EC A8 99 75 E3 3D 09 9E 64
 A2 F7 A7 D7 38 5C 56 21 37 83 E8 6E 82 96 E4 47
 48 1C EE 48 43 35 A6 51 C7 A8 96 4B 17 F5 6D 0F
 76 EA 1C 23 F8 31 DB 84 DD 79 04 7C 31 5A 14 B0
 B4 E5 D8 B8 FB 26 8D 4A E9 1E F3 5E 21 5F A3 B2
 B4 E9 B5 83 FF 03 1B 5A A8 04 C4 FE 64 53 C4 1E
 3C 99 2C 5C F3 55 E7 7A 5F 99 B7 7E BB D8 5A 88
 F6 2E 05 49 C9 74 A3 0D 93 97 33 7A 67 33 D1 C7
 EC 9E 13 A6 DA C9 D6 6A 40 FC 7A 70 2E 4A CB 5E
 BD 27 BC 25 A5 F3 03 F8 17 80 46 FF 51 66 04 0F
 C6 E8 41 C1 FE 92 62 53 35 F2 29 89 19 34 01 A3
 E9 2E 0C A9 DE 50 62 71 07 26 2E E0 23 FD AD EB
 0C B9 B2 55 40 60 92 6A CE 04 B9 9D 35 B4 6A 06
 8D FE C7 C9 40 6F CE 1F 78 5C A7 45 36 79 81 1E
 DE 3C 9F 7F 10 92 1D C4 47 DA CE 62 8F 18 3C 20
 57 DE 66 44 AD C4 70 86 F1 17 00 66 96 35 AD D9
 46 77 4F D6 BE 9B E0 7D F1 61 BD 54 1E BC 64 BB
 49 13 63 83 22 EB 37 40 8B 6A D7 AD B2 92 63 34
 D6 A5 0D 12 0A 03 01 FC 5A BC 64 D7 A9 61 E6 7F
 41 5B 79 59 9C 26 F0 7D 35 EB A2 EF 39 47 36 79
 9A 3D 66 A9 ED F9 E5 85 67 F1 31 C9 D8 07 90 53
 74 FB C7 D0 4A 01 A6 49 B2 DC 23 6F 78 11 31 F4
 F1 01 57 18 6D 18 42 94 0C 1B EC A4 78 B1 7E 22
 65 95 9A 9F F4 4D D5 E9 5A 33 07 98 41 57 2A 84
 3E 07 0F 9A 7F 9F 28 87 D8 B5 97 7B 5E 96 4B 4D
 84 5B 19 38 E7 14 2B AC 23 EC 9E 38 5E 9B E8 B9
 A5 29 6F 64 EA 4C 93 8E 28 60 29 3B 07 A5 51 50
 C1 23 D5 FE 21 D3 2A D5 59 AF 60 C6 58 65 5A 8C
 D9 46 8F 60 08 2F 29 D6 D8 EF 40 FB CB 76 CE 1B
 5A E2 BD 25 06 FA F7 F1 AC 78 EF 92 7E 02 3D 17
 89 B7 D7 42 B1 BA A0 C1 FB EF 10 CD BC 6D AE 65
 B0 E2 57 C9 97 B4 A1 3D EF D0 60 4E 9E 42 D7 EE
 3A 37 FD D3 76 25 1C C6 A0 EF 98 53 76 4A 2F 10
 E5 1A AB FB 18 4B A5 91 C3 D3 EC 69 A5 23 F6 F2
 7D 6B 02 12 3F 4A 10 A1 7C CD 15 F8 A2 23 6C D9
 66 9B 0B 6D E3 04 41 68 46 38 85 A6 1F 59 21 2E
 32 52 5E B7 C5 E6 8E 36 43 9A BA 4B 00 0C 46 07
 6E 8F B4 CF F3 AF C6 D8 05 AA 50 8C 12 0C 7B 9F
 AE FE 88 83 C7 63 1D B7 0A 3D 4F A8 46 EA 02 C1
 2A C6 FF 38 03 7F F9 F4 B3 6B C8 FD 86 17 0B C8
 FC 72 0C 1A A8 BB 0A 01 6D 24 46 90 F9 A1 82 DE
 29 EF B8 CD 29 4D 7A F2 E8 6F 49 D9 3C 93 47 5C
 BA D3 D8 5F 86 83 83 72 B7 8D F0 86 9A 9C D6 AD
 A9 AD D8 50 32 0E FA 3E 71 E9 E2 70 6F 98 16 37
 C9 41 A2 09 B8 91 4D A6 C4 8B 19 6D 81 6D 0B 5A
 E2 DC C9 E1 A7 ED D2 1C 95 B0 81 5C 8E 45 CF E6
 DC 1D D0 20 6F 06 3B D9 45 3F 2A 6A 9C 2D CE 8C
 C2 16 02 47 0F 00 CC 80 1E BA BA 44 31 4B 9C BB
 53 01 01 08 A6 61 79 41 FD D9 97 02 0E A7 8F 53
 66 C3 3F 5E BD 14 5D 1D A4 B4 B2 A5 D3 55 DB 5F
 89 2E 19 77 52 AD AC F7 3C BF 78 FF C2 6A E3 01
 64 BD F7 C0 7F 0C A0 2F F4 D5 BB C3 1E 51 F4 AA
 B0 03 88 53 FE AA 9D 2B F6 36 A2 CC 5D 08 8E FD
 F8 4C B3 74 21 E6 04 1C E9 48 99 CE 46 DC 47 C5
 8D CB 70 B4 7A A3 1A 96 F8 C8 CA 19 E4 F2 2B 75
 AA AE 38 78 91 B8 41 C6 CB ED 06 51 55 F2 52 A1
 90 F1 43 EB 35 FD 01 42 17 A4 C5 24 6A 73 8E C7
 F0 ED D9 E1 2C CD 82 F4 D3 EE 20 88 FA 20 60 1A
 05 17 7C 97 65 C5 D6 D6 90 0B 63 0A C5 11 89 A7
 90 6C 1B 06 C6 68 5C 17 2E F9 D7 67 19 6F 1F CE
 5E D5 34 4A 23 88 47 70 F2 77 08 71 7C D5 DE 7B
 7B 64 99 2A BB 85 99 48 8B 14 A1 51 25 DE E3 4F
 28 36 BE 73 B4 16 AD 81 34 29 B7 A1 EA E4 DE B8
 BB 4D 8E 40 5F FA D6 E9 C9 24 AF 72 31 4C 01 F2
 BF 87 91 84 5F 33 2B 89 00 F9 E0 C7 CF 1E 5D B2
 7F 30 31 5C 6D E2 7F 75 32 66 EB 4D B5 37 7D 68
 9F 2E 9D 79 33 1E 92 C4 1E 61 F2 AD A1 85 A2 83
 54 BA CF A6 82 E1 E9 EA EE 1D 38 A5 C8 D4 21 11
 40 EE 17 2A 07 61 8B 66 00 81 A0 4F 3A 35 C7 59
 04 C8 08 20 9A 47 8E 39 E5 22 9A 64 C4 E7 AC 2D
 BA 36 14 64 2D 92 56 27 F1 D5 DB 0A 37 9A 65 EB
 14 E9 58 01 FB 51 50 F9 47 0D D0 1A F2 12 76 C5
 00 91 EF 96 70 18 EC 2A 93 00 DA 33 7A 22 D4 D9
 CB 38 F8 7F 44 47 07 F4 94 34 EC 93 28 74 3B FD
 34 7D 81 D0 29 34 6B 22 FD 35 5B 33 58 5C 43 BF
 AF A1 D4 11 79 16 15 C6 98 3A F4 A0 B3 5F 9B BD
 6D 01 78 0F 60 3F 16 90 C2 46 E4 3E 0C 98 D4 6D
 02 BD 23 72 7D C6 99 85 9F 15 45 25 1E D7 B5 CD
 01 A8 B7 F8 87 C6 09 C9 61 E7 E8 4C AC 5D C1 C9
 4D 58 58 06 D4 19 92 88 4E 38 41 07 A0 8F 7C 73
 89 7A 05 64 B5 AB 81 38 D9 17 86 81 D4 2E A2 11
 31 02 5F 3E A1 A6 87 7D 8B A1 59 D0 F9 D6 8E 8A
 A7 CE 69 EA F3 7F 11 88 20 E6 E6 66 DA 55 00 71
 68 F4 4C 7D C4 DD EF A9 C7 3B 52 07 3F F1 88 BB
 AC 69 8F 5B 89 43 3F 20 BB 2C 10 D7 38 D0 82 65
 13 66 F1 77 E7 FF FE 6A A8 76 09 9B C2 0C EC 9D
 38 D4 1C 27 70 C4 88 6A C7 6D 02 11 39 CC A5 08
 DA E5 5D B3 9E 7E 26 1A 59 CC 6F 16 D5 FF 4B 91
 AB 6D 20 BB 3A 92 17 A5 DA 0B D7 C8 D1 E7 F5 B6
 83 B5 25 AD 62 C8 5E 45 D5 FC 72 C9 A0 C9 D6 45
 F1 8D 84 2D CE A1 B0 CC D4 89 81 69 1A 53 42 EE
 10 1F 96 69 A9 94 A8 86 D1 13 01 27 94 51 B1 82
 89 3B 2D A3 64 E1 3A 2C F9 30 10 49 A9 C2 93 41
 25 F2 14 B2 A4 BE FC 44 53 40 33 E5 D9 AC E4 0A
 CB DD CA B6 3F AE D6 F9 6E DE 73 7B 41 15 8A 09
 FC AE 3F 15 AF 83 3F 9B B8 54 13 E1 8D 72 47 DA
 1F C2 40 DF 64 49 CB 63 AF EA 52 95 2C 51 12 34
 3C DE C4 86 0F 3D 13 D2 31 5F 6B 3F E8 FF 61 28
 4B 9E 23 14 46 E2 AE 56 1E BF 1D 3B CB C5 10 97
 33 6C 1A A1 2F DB 95 3E 20 39 40 14 A2 E6 41 59
 1E 70 E9 A7 26 B2 D3 7A 28 2E 1D 37 B3 34 7D 15
 A2 46 DA 2B F4 FD 1D DB 9B 56 11 B9 30 F0 7E 0A
 E3 1D 4E 03 94 26 78 22 B1 96 66 7A 70 84 1F E7
 E7 22 97 8E D3 E3 2F BF DF B6 78 2E 3E A3 2D 38
 62 A9 83 0F C3 46 A7 F4 E3 88 35 58 CB 32 92 EE
 76 84 F6 0E 44 9B 46 B2 B4 58 D9 FD 93 D7 11 F1
 BB 3B 77 15 0C 6A 48 AD 7A 6D AB C7 B7 F5 F8 4E
 2D 4B 55 03 78 AB 1F 37 64 8B 69 0F 0F 27 44 F6
 E8 AA BC 53 83 08 FE E9 BA 67 CF 30 3D 07 B6 DF
 B9 9E 4E 4D FE D7 41 7F 20 E9 AC 5C A6 E9 0D 78
 46 9A 43 55 62 32 45 DC 34 CF 01 5D DF 56 90 E4
 4C 4F 23 F8 58 DE BE 05 5E 8E 99 80 D7 F0 A9 9E
 64 5F C3 D9 DA A9 DD 6F 22 0F 57 F0 86 42 0C 18
 E5 92 93 A8 AE 4E 84 1A BF 53 BA 2A C5 05 0A DC
 9F 6C 4D A8 39 0E 5D 0A 6A 41 66 9E 78 3C 6C 58
 8A 50 2C D3 AD 56 A9 2F 3C 67 4B F5 D3 59 E9 21
 10 EC 42 F4 47 D5 15 BE 3C 40 A3 9E B3 97 F6 A8
 DE B7 26 CD 7E 6D 1C 58 2C 31 DF 48 7B C3 11 27
 17 B4 47 2D C6 3B 94 6A 02 D1 AF 15 71 52 C2 A3
 C1 E7 29 00 6B F2 28 71 5B 34 CA 10 B3 65 23 93
 F8 77 C6 9F 0E BB 15 29 70 96 50 0E 07 6B 02 15
 95 23 26 FF 0D 94 B0 E3 BB 2D 93 0D 20 10 B9 31
 09 37 EF F1 8E 51 74 A3 03 95 FD 4B B2 89 57 83
 B9 7C ED A9 AB E1 52 78 97 71 11 5B AD 71 5B 4F
 85 D7 F3 EE E1 F8 34 B5 CC 11 CF A3 C0 24 C9 12
 C7 66 FC 1A 79 3D BE 08 F6 37 BA FA 98 D3 6C 09
 0E 4C C8 F2 7E A6 AA 63 D8 E7 4F 5B FC 19 5B 96
 D0 C3 B5 05 BA 7B B9 02 5A 1D A6 C3 C6 A6 4F 18
 27 A4 E9 30 8D DF C8 50 CA F8 01 50 86 52 17 95
 DE 6F 59 2A 65 96 53 56 AB B9 A9 06 77 F6 8B 4C
 9E 93 1E D8 73 B9 B7 A7 1B FE D0 05 39 09 74 E2
 F1 36 C7 B2 91 C5 4B C8 96 C2 4C F1 52 76 33 EA
 D9 51 EB EF 0D C6 3E F0 6D 87 9A 54 68 79 22 DF
 D5 95 78 75 F4 1C 26 2C 3F 59 79 E4 C9 EB 64 DD
 25 53 BF E1 42 37 FC CB AC 10 52 E4 7E E1 A2 6E
 BE 05 17 3A BE 0A 60 07 DF 04 31 EE BF 51 8B EB
 AD 91 7F 7C CF 60 13 90 7A B9 FC EA 41 39 14 37
 38 3E F6 9F 8A F5 F6 BF 83 64 69 C8 29 77 18 F7
 E0 FC 65 70 78 6F 05 FE 47 2A F1 9D 67 05 24 19
 7E 54 FB 68 33 75 4B 8D 37 85 18 CE AA DC 78 39
 42 9A 0F 29 AC 14 CC 36 7B 4C 87 AB A7 42 C3 59
 15 6C 14 45 25 D5 D0 62 06 3E 4D 4D 63 AB 55 62
 A8 62 9F 50 6B 91 33 EC B1 5D EF 16 45 5E 38 77
 34 48 40 DE 01 DE DA 0E 20 82 77 8D 8D 53 47 96
 59 EE 23 20 53 D0 AE F7 94 D8 97 96 85 55 0D A6
 70 0B 68 51 5B 92 F9 BC 3A 77 ED 4F B4 62 F3 26
 0C 59 3E 36 C0 88 B6 6E D6 48 53 06 E0 0A AA 96
 07 C4 53 3A 9D D0 B0 2A C8 E7 65 2B C3 6B 21 8F
 7B B5 A1 5A 99 D5 0B 76 08 EB F3 AC 12 18 65 CF
 9C 45 93 53 76 AF 28 59 9F 28 EC 14 91 CD ED 73
 AD 24 AC D4 73 F8 F2 19 62 68 9D 71 2D A5 D8 76
 B1 18 94 09 EA 46 27 B8 E6 1A B0 5F 14 70 0A 3B
 C2 3C 50 96 06 89 AD 44 0C 4E F6 F2 70 AB ED 4B
 64 12 1F 1D 24 09 C5 DB FC 0F 59 09 E6 CA C6 F5
 77 D0 4A 12 9B B4 FA 2E D5 1A 37 49 23 03 95 10
 1A E8 A8 E4 E1 ED 37 E8 C1 75 1B 25 FD 9C 47 C9
 78 51 63 3D 0A 3C 4C 00 56 0E 75 83 C9 C3 4C BA
 C2 B9 02 D9 06 52 FC 17 90 3A D3 B3 F4 A0 BF AB
 60 05 1D 33 51 1C D6 CF 9A 82 62 9A 0E 1D 25 C5
 5E 47 25 52 69 2A D1 D0 F2 42 7E 9D B3 45 B2 8D
 D9 1F BA 92 03 2D 3E EF CE AB 44 F8 DE 8A E5 4F
 17 D4 E2 01 27 30 35 E1 B4 02 57 62 D1 1A 46 6C
 3A 80 00 FC C4 EB 25 8E D7 62 EC 07 B2 01 31 40
 64 0B F6 F9 E5 8A 38 ED CE 70 65 66 E2 5A CA 76
 ED 91 94 F4 01 B4 2F 01 CC 0D A0 D3 AF 12 5F 4F
 91 4A E2 70 53 4F 48 25 B0 88 AE 2B F9 70 EF E4
 AA 89 EF 3B 00 81 B1 AB 4F A7 89 7C CF E1 B4 20
 C2 F9 C8 91 8C 21 0A 27 9A EE 98 7B E5 18 8A 0B
 75 B8 F2 D5 95 F4 C5 D2 21 91 FD 22 B5 D5 9B A6
 CA 88 FB 37 F2 86 B3 F8 99 17 13 A1 0F 53 6C E1
 66 A9 69 1B 57 9A 9F 7E 71 CC 1C 10 7A BA 48 AB
 0E 2D 2D 9D 1E D5 A8 79 77 16 BA DE D6 C7 01 DA
 40 60 BD 19 2A 58 44 7C CC CA C0 E6 74 60 2D 8A
 64 6E CA C3 BF 7C CF 78 73 FD A3 5E AD 39 2F 03
 94 AE 1B 89 A2 79 6B 51 9E 8E 57 2B 4D B5 78 56
 52 C1 1B C3 EA 9F 46 01 9E 80 61 78 AE B2 E8 B4
 66 9E 90 0F 3D A8 09 77 6E A7 59 22 85 29 86 D8
 07 64 7B 90 3B 4B C2 5D B9 03 3B 90 F9 1F FA 90
 85 7C 69 B2 53 B6 21 0E E6 BC 35 84 A4 07 0F D6
 96 C2 EE B6 B9 9A F4 78 4F E8 08 79 9C 48 ED 50
 C7 84 E0 A9 2D BB F0 DE AC 8F FA 7A 34 8B 83 83
 C8 19 B0 4D A0 E3 56 A5 11 28 DE E6 AF CA 9F 37
 20 8A EE E7 06 06 23 4D 57 E9 EA A8 38 27 63 67
 E6 CF D3 9E A6 14 C6 FD 5E 91 69 BF 2D 38 91 1D
 58 EA 7C C1 24 5E E6 98 56 58 4A A9 91 79 6D 0A
 34 40 14 4D C0 F5 93 46 28 C4 8B F1 EC C3 E4 0C
 E8 E6 08 9D 53 73 6B 2F AE F8 68 53 2B AA 21 B3
 8D 99 86 06 E9 23 86 63 C3 ED 8F 0A AB 96 9D 9A
 0D B9 2C D5 7C 9E A8 82 B2 85 01 46 F7 20 74 58
 0C 9A 8C 0B 96 21 4B 5F C4 86 38 23 6E 3B BE 0E
 F5 D4 C8 5D B7 FF 83 6D 21 E8 F9 06 3D 09 04 B2
 FE 42 14 C8 FE 50 A7 7E C7 61 D4 93 3C CF 74 6F
 6A 18 B8 03 BE C6 4C D3 DA 1D A1 31 E3 5E 38 87
 88 72 B6 A3 A5 7E B4 5A 33 5A BB 08 B3 0E 51 FA
 4B DA CF 22 D4 A6 DE EB 42 D8 C7 FF 63 C2 D7 A2
 85 2F 6B 0F 72 45 6A 3F 5D 61 BF BE 55 AB BE 2D
 60 04 9C EE CC AF 8D AB 0B 12 AC 5A 75 93 76 B0
 06 59 90 D7 DF 8E 28 61 2C 11 DF BD 69 3C 69 A4
 7C E8 32 98 33 34 A3 10 A5 12 D4 AF 16 61 EC 5D
 84 55 FC 04 A7 4A EB FA E6 A5 5D AB 2F 98 1E 02
 5A 90 BA 21 3F 96 2E 5B 43 29 11 EC F2 47 69 55
 07 DC 79 6F FC 2A A4 4E ED 33 94 4C EC 64 F2 E1
 B5 90 D2 02 81 5A C2 15 32 82 25 3E 2A C5 A1 39
 2A 3B 5E EF 59 DC B9 FF 7F 61 E2 CC E1 8F 47 7B
 55 38 40 9B DB 6B 55 7E B8 1F C5 32 93 09 4B A1
 9C 2A 07 B2 94 26 58 35 70 24 86 9D 05 28 92 17
 D5 1D 51 1B B9 C6 8B ED 10 F9 0A AB 1E 7D 9A DA
 32 15 60 1C 45 80 49 DA 41 7C B1 24 08 8D CF 13
 56 9D B8 38 62 82 04 46 E9 55 C2 77 4B 79 B7 79
 B3 FA D1 96 D0 52 1D 68 B5 F8 D1 28 D5 2C 14 94
 DB 0D 90 94 8F 32 B2 77 73 0E BD 08 56 E5 23 4E
 06 08 2D F1 87 2F D0 CB 95 E8 F4 53 D8 15 61 DA
 FD AB 33 D2 7E DC 1E F5 3F 92 71 83 9A C3 6F 84
 A6 52 B3 BB 4A 6D 3D 1D FF 4D CB E6 55 96 B4 ED
 60 24 B2 A8 11 CE 94 5F 0C 10 87 F9 8E 9A B9 78
 0E 7B 84 68 65 19 9E 80 CB 6B E9 B3 56 6B 90 E8
 42 0A 30 12 E1 DC BE 73 10 B2 E1 C3 66 8D DD 72
 C8 2E A1 F0 46 53 3B 00 4E 24 C4 4A F3 1F 2B CE
 F0 E6 04 F3 43 24 92 43 6A 7F 1C 89 E7 F6 F9 93
 F9 F2 79 ED 7F 0D 5F 6D 62 D4 83 3B 4B B9 76 59
 79 DB 42 EB BC A4 93 3B CF 48 FF 6D F2 2D 42 61
 23 90 FD 1A 2A F5 65 CE 68 8A 68 32 FB AF 8D 5D
 0E 5D 86 FE 15 5F C0 07 8B D9 33 62 30 27 BD 4C
 7F A1 D3 14 AC E6 DD C2 0A 39 E9 E3 8F 69 82 66
 67 5E 41 79 A7 1F D2 EA 1E CF AD 47 56 B3 26 A2
 BF 52 82 9F 7B A8 58 1D E4 7A 98 24 49 0F 11 03
 A8 D7 A7 96 25 4D 37 38 63 61 83 7E 52 3D 36 24
 BD B5 7B C8 14 D0 A5 CF CD 2E 55 CA 88 8B 2E 68
 9E DE F0 0F 0E D5 BB B7 E3 A1 B4 98 B8 36 92 E0
 26 EC 63 FB 9D C4 E9 39 F8 3E D2 DE F2 3E 4E 01
 64 82 37 4A 42 AD AB EB 37 51 5B 16 A1 5E 38 36
 50 13 32 91 B4 7A 00 B7 FC B1 66 0C 8F DD 5B 6D
 76 20 83 4D 34 6B 88 3B E5 02 9A 08 0B AC 08 F4
 54 5A 66 82 7A 9E 95 A0 8D DC 9B A3 62 75 E9 09
 67 31 3D 90 24 21 F7 75 36 DF C7 38 EC 61 E8 24
 4E 45 E7 95 5E A1 A3 4C 0F 44 EC 76 94 2B C1 BF
 BC 42 85 7E E8 C6 82 51 8C EE 4A B7 94 93 B5 86
 58 9E FD 04 D2 74 C7 AF 21 95 F1 3D 14 82 D5 57
 B1 10 82 BE B1 B1 A5 F7 A1 5A 17 C2 59 8D CB B4
 3F 48 46 11 80 F4 F6 80 55 1B 7A 69 72 20 BC 05
 55 A0 C2 81 B2 F0 B2 F4 0C 2C FB 47 45 5E 4D 42
 1A 58 BC 1A F4 06 F4 F4 6E 2D B3 F5 D9 F7 86 F7
 A6 E5 B7 C3 BC AE 20 79 ED 7A 5D E3 32 35 5D B5
 4A 42 93 40 09 37 17 52 BD 2C 2D 7B F3 3C 41 48
 27 54 36 5B 8B F8 EC A6 E9 55 C9 DB 28 95 17 69
 78 F9 D3 9D 35 5D CB 15 60 A8 D1 5C 45 FB 52 44
 31 D6 BF 82 E2 78 58 DB A2 AC 9C E3 44 6B 37 A2
 54 64 C6 89 6B 74 82 A6 C2 A6 49 63 F2 2F 1A 9B
 A7 FB B2 53 01 FB 48 57 29 5A 8E AE 35 63 22 C4
 47 3E ED BC FD 19 6C E9 11 C7 95 CE E6 85 90 96
 FA 2A F9 D8 46 BB F5 1B A1 27 8B CF 5E D1 E1 17
 37 79 F7 41 69 B6 07 D9 D6 12 40 FD 81 30 86 03
 AE F3 28 B2 FF 44 F6 35 20 12 FF CA 83 2A 2F F8
 53 65 DE 61 97 51 C7 76 CA 48 44 C1 D2 68 6F 03
 53 CA 01 B5 BC 7D BA 9A A5 D8 75 E1 01 3F 88 2E
 24 2F 05 98 47 1C 75 E4 EC F8 ED 0A BD 5D 1C 74
 FD A0 05 46 EC AA 5A 98 66 AC C4 64 F8 93 C8 2A
 C0 DB 45 E0 D6 3F 06 0A F4 20 F4 49 37 88 B6 63
 B5 9D 2E D2 8F A5 A5 81 23 55 6B 87 B5 65 DB 32
 51 DC 8E 30 BA 41 F1 72 BF 2E C8 C5 26 4D C3 F7
 22 9A D7 05 CC A0 24 58 CD 33 56 47 80 FB 8C 0C
 5B 9C ED AA 28 3D 5A 6E 8C 25 12 5C 77 8F 29 E2
 CA DD 8B 11 F1 47 58 B0 97 7C 0E 32 FB F6 56 3B
 84 D6 27 CB 57 60 0C 17 6A 51 DB 23 03 C9 34 F6
 B6 FF 74 73 07 E2 75 72 B5 A0 17 9B 07 7A 6B FC
 42 8A 46 3E B7 E8 27 50 0B 87 49 26 36 32 53 5F
 86 AD CD 13 1F B7 A7 AD 85 A5 81 B0 11 E7 65 EB
 2A C1 BF B2 AA B4 25 7A FF A0 EB 8E 72 CA 3F C9
 3E 4D 3E 49 11 1D FF 31 A4 D8 18 D6 5A 96 E1 4B
 BF 74 FC BC F3 BF BD 01 18 69 93 30 E6 B9 9A 79
 3D 05 94 ED 2F BF 0F C8 42 1C B7 AF 62 AC 64 5C
 B0 41 4F 42 7B 3F 88 ED 90 28 BC 8F CD B5 60 DB
 26 25 28 BA 82 70 05 32 FC 9F CD 6E ED B0 B1 52
 86 EF A1 B5 14 4E CB 1F EC B9 D2 D7 F0 81 03 37
 90 99 90 70 C2 3A 02 15 FB 9B F0 6F E3 D8 CD CD
 FC E7 56 BE DF A0 3A 0B 6A DA 3D 9D 12 A9 92 6F
 A5 AB 13 9C 71 81 40 72 E8 FB 45 83 8B 7E 44 10
 B7 27 FA F8 A7 48 EC ED B8 CE 5A 1F 9C 62 AB B7
 C3 46 3E DC 14 87 49 98 1A D0 7D 15 34 FD CE 66
 39 8E BB 8B 4D C3 DB 87 28 3C E6 45 27 E3 4A 87
 C4 37 44 F4 3F 42 21 44 FC 7C 72 0B 3C 09 EE 7E
 0E E4 DF 1D 9B 53 B2 29 4C 13 E9 E4 B6 73 23 2C
 17 C6 E5 DB 39 2F 55 12 BB DB E5 6A 1E C5 CB 65
 02 8F 03 2E 50 48 7F 35 1B 06 06 1F BA 6E 5D 9B
 E9 35 7C 66 9A 00 E1 16 B5 20 64 1C E9 00 27 AE
 8E 57 15 5F 4C 4A 64 AC F1 92 5E F8 FC BC CC 57
 27 16 93 BC F7 79 18 9F 4A 63 6D 99 5D 29 1E 6A
 02 E3 FF 9B 8E AF 68 20 A6 A9 92 68 C6 C8 2F 0D
 AB 05 EA 24 92 A5 98 B3 BA 51 AF D5 7C C8 5F BD
 D2 0F AA 9A BF D0 6A 84 95 8F B8 6C F4 36 C6 3B
 C2 3F EF 37 19 0D 14 CD EE B4 BE D8 3E D5 4A 99
 FD 49 B5 E3 78 43 6C 13 1A 3F 8E 23 7B D0 1D 0E
 A6 45 75 BA 19 3B F8 13 57 7B 05 E1 B1 5B A6 70
 37 C1 46 F2 45 3F 45 EC EB 01 7A BC 27 C8 68 44
 DA AB B2 C6 94 B7 3F C3 52 F3 E3 0B 34 DE EA 17
 B5 4D F9 7C 0A 24 E2 62 90 3C 54 FB 76 19 03 A9
 AF F0 08 CE 74 05 A2 C8 B7 00 4C 8D 1C 16 AF 2B
 41 A2 E8 EB 45 DF F0 8D C7 6D EF CF B1 DF 2A A5
 30 1A 0C 40 B1 F3 29 00 B2 A4 EF AD A7 0A 61 B5
 E9 E2 9F 6A 37 5D C9 73 69 4E BE 8E 93 05 4F 7D
 9B FF 86 A6 57 3A 6B 9C 18 78 8F 72 82 D5 09 2E
 C5 30 DF 29 8E 5C 61 AB 3E A8 11 2F AA D4 C8 11
 80 F9 C2 6A 83 DC 94 4D 84 16 88 10 23 D9 D8 89
 3D B8 F8 27 68 4C DB 1E D0 15 0E 2A CA 61 CF 24
 DB 20 4C 16 D6 30 87 5A 33 34 10 64 BC 82 22 D5
 82 71 48 8A 74 7A D9 8A B8 A3 A9 C2 CD 4D E7 12
 B0 65 E9 03 D0 CF 08 02 E4 35 9C 6F CF 0F C5 D7
 73 36 F6 4B 2B 27 74 7A FA 8D F6 1F D1 95 77 EE
 19 2A 96 2E D8 A7 20 7F 66 87 69 88 7D 82 35 1A
 8D E9 5E 16 93 BA CE 72 1B 2E AF 1A D2 AA EE 74
 ED DA 4C 21 C3 FA 39 ED 38 B9 A0 EE B2 CD 66 0B
 FB 28 BF 56 AF 6A 3B 6E F0 FE B3 77 BF 56 37 22
 6F C8 46 A4 B8 C8 19 53 E9 58 00 A4 CD 3E 2A 16
 8D 21 06 88 E4 BC 80 11 F6 55 CB 34 FD A4 CE DF
 D7 81 2C 6D 7F 25 E7 44 DD 46 AC 16 6A 1F 1F FF
 A8 94 19 AC 0A EA 4E D1 47 5F 63 2D 76 41 CE EC
 CE B9 7D E4 94 14 1B 75 45 0C 51 D6 F1 80 4C 4E
 38 3B A5 6F 43 81 A3 43 56 F8 A9 8C C9 CE BE 26
 18 A5 89 B7 E4 DA 75 CB CF 48 8E FB 02 7C 83 8B
 12 F5 E7 1F 58 4C 66 C8 21 F0 BF 0D 73 EF 06 53
 66 EA 91 5D 1F 18 06 89 95 78 9C 79 DE DC 38 EB
 59 CB 45 27 F9 11 4B 04 BD BF 91 B9 AC 54 39 ED
 07 D3 5F 07 F3 F0 5C CE D2 6A 67 0E 8D 04 D3 01
 71 AC EE 50 40 11 F6 1A 38 2D 2A 91 72 8E BA 9F
 4B A7 93 EA 71 B4 E9 63 B0 1F DB F0 2E F5 39 76
 99 CA 0B 0D E5 5C 19 43 90 83 4C 68 C5 3F 21 90
 9D 1D A7 2C BD 8F A3 D1 ED BD 14 63 D3 1E FC 14
 CD 2D 72 59 85 B8 AF CF 1F 61 0A 14 A4 F6 B9 E5
 4F 64 EC 20 B6 22 D3 45 7B 2C F9 6D 9C 5C 98 99
 0D 70 D3 9C 9E 84 BE A0 B7 71 32 68 12 81 49 E6
 4A CE BD 80 0F 2C AC 5E D7 D3 3B 2D F8 EC 6F 22
 A9 4A 93 8E B4 05 B5 EB 65 0D 81 C4 D9 20 B3 EC
 D8 0A 7D 42 74 A6 CD B2 B3 7D 03 49 BE 08 CC A8
 22 C7 FB BA AE DE 07 73 2B D7 20 3D 43 DD 8E BD
 D8 8A 27 F7 06 52 75 98 4B F5 5D A8 B6 0D 25 BB
 10 C2 6D 81 8A E3 59 D9 7E 25 0C 49 D0 97 62 72
 E3 2A 02 FF B6 ED 2B 8A 16 F6 98 FC 28 CA A6 E1
 BD E8 98 63 19 12 F1 54 76 38 16 4E 23 CA 84 C8
 D4 FD E7 54 31 45 66 F7 37 AD 0E 42 D1 B6 67 CC
 C5 F6 65 26 6C 59 E7 91 C5 1F FF DC D0 B4 A6 FB
 DB B5 A1 6F C9 14 E1 78 B5 98 01 24 9F 96 11 05
 B0 E3 0D 2F 57 C7 E8 14 23 C6 4C 32 65 F0 87 C3
 59 8E 83 65 58 10 7D 48 7E 53 DB 51 C2 19 22 D4
 D3 3A D9 BF 87 30 D7 8F A8 60 9C 3C DD BC 9D 77
 6B 23 84 30 FB 78 DC AF B2 3B AF 09 01 0F 14 E6
 52 5C EF 7B 0A 17 40 EC F8 5A A0 56 46 D7 97 9E
 07 02 71 55 69 13 76 55 63 17 10 6B EC 08 B0 A0
 FB D1 E4 63 01 41 C5 8E DC 39 34 F0 FF 73 6F 95
 65 B2 AE DC 30 0F 86 E9 54 9D FB A4 EC 7F D7 C7
 B8 07 88 5C EC DC AC 38 C6 78 E8 8F C6 7F 5D 1F
 6A 5E 6D B7 42 EA 4D 97 94 57 4A C1 6B 8A DB 8D
 7B 0D 10 6D 36 95 3A CC 8E F5 9E DF AA 00 00 EB
 09 E9 32 32 84 7D 6F 89 19 B8 55 E7 68 0F B0 23
 70 61 45 86 FF CF CD F0 4D 84 61 7F 7D B3 0B 9B
 40 0E 98 07 10 3D C6 3D EE 06 2E F9 12 18 A3 2E
 C8 4B 7F 22 8F 37 F4 AC F3 76 52 E1 EE 72 9F 05
 0D D0 F3 86 48 2A 3C B4 7E 3D 1D E4 B0 8A 52 B5
 8D 39 A5 9B 4A 3A 61 45 64 49 5D FC CA 92 54 DD
 69 BB 85 AD DC D1 64 6E C4 7B D3 ED 53 F1 12 51
 65 C4 18 B2 D9 68 15 43 48 34 9C EB A0 EA 7A EE
 3B 2C 39 9D 18 ED 8C 8D 3F EF 16 7C 61 95 84 3C
 F8 B7 56 3B CE A2 36 34 B2 01 22 38 34 31 02 BF
 6D C7 8A C5 69 88 B5 89 C6 E0 44 84 79 DE 52 D9
 53 70 BC 76 1D 35 68 2A 76 70 AC 7F C5 B7 76 2B
 20 BC 6F 12 24 64 F8 DA 6A 5E E2 31 76 2F 54 82
 D2 43 2E 92 00 9F EE F5 8A E3 7C 84 FA 93 C3 E9
 CC 10 37 E5 4C A8 93 86 73 21 8C 7F F9 4E 1D 3C
 0C 57 F3 43 C6 C1 70 15 C3 3A 75 9A 44 C2 90 72
 44 50 16 C3 DE CD FE CA 22 8E F4 63 EA B2 7B 28
 8F 94 91 4C 6A 78 91 B8 BA 06 FD 61 E1 F8 86 A4
 AB 93 A5 E6 E0 BC 0C 6E 12 9E 22 8C 43 EE 42 AD
 88 AB 00 66 AB E6 67 E4 97 51 20 71 33 FE 11 72
 B8 78 C5 98 D9 AD 1B 4E 7E 81 75 18 A1 0A F7 35
 DF 0D 1F B5 34 61 C3 7D FA 42 0D D9 3C A2 44 A5
 69 6B B3 65 CE BB 02 A5 41 4F 61 76 D7 F4 19 B7
 4C B6 05 D1 03 1F C5 10 B8 D7 D8 C6 2F 0F E0 9C
 DD D0 3E 38 49 51 3D 50 4E 9E 04 5F 93 12 14 A5
 0D CD EB 63 D4 52 E6 5E 8D 5F B2 2F CB B2 0B 32
 F1 10 6A B8 8B 89 72 54 97 64 8F E1 E7 52 40 9D
 24 CC D0 AA 8B BF FC 00 F5 8F 10 BD FE 52 AA 55
 49 7A C9 1C 97 CB C8 02 8F 29 8C 23 05 7D 08 9C
 7E 71 0E 58 0A EF 9A 19 DE C5 FC BB 29 17 66 6B
 51 E4 97 2E 05 14 B7 FA 6E 18 CA 09 DF B7 60 4F
 1B DE 31 B1 E1 F0 87 99 E3 D1 11 00 72 60 9C BE
 CD 7C A2 0F 97 FA EB E2 4B 1B 4E 96 E8 F2 42 36
 F6 72 F7 62 27 E2 44 2B BE 29 DE 6A 88 C0 C7 E4
 DC D5 DA 48 7B 72 5B 89 C4 B3 8F CE 09 1C 17 67
 02 75 31 67 49 EC FF 76 D8 DE 32 78 39 AA 6A BB
 51 DE CA 4E 55 5E 03 86 B3 B8 93 FA 1C 95 8E 06
 FF 63 22 83 E9 86 73 C9 45 36 C1 53 C8 CC 4A 7C
 6D C5 00 CE 75 4D F7 96 7E 05 FE 33 DC 22 41 C2
 AF 2E 9F 74 77 9B F8 AB 51 CD 8F 81 25 6E 4C 56
 13 DE 35 1C EF B6 F5 E7 25 07 92 B2 3B 6E 86 2D
 40 67 63 53 D6 0B 8A 6C 0C 3D C1 EF 36 57 60 34
 66 E9 30 61 D3 57 17 44 37 10 27 A5 FA F9 17 25
 A4 C2 FD 56 9F 56 F4 FA 3F BB F3 D0 10 DA FB 23
 BF 56 A8 A5 0C D9 EB 10 09 46 6A 34 40 FE 27 A0
 F0 45 61 29 9C E8 0C D7 BA 3F DA A5 B9 2C CD 38
 92 1E 0A 69 F6 4E 9C 0A E2 22 0A 35 55 23 13 2C
 B7 AD A6 54 27 03 21 88 B6 9E F3 54 98 55 D4 42
 2E 54 C1 D5 72 95 48 61 72 64 C4 5C 8F 62 E0 EF
 B4 C2 9C 7A 2C F1 02 59 E6 E0 DF 5B BE BD 8A 39
 24 1B 12 31 2F AC 61 BD E9 23 A9 A1 0F CD FB A6
 19 54 78 B5 59 CF F1 78 34 E4 E4 28 F9 89 88 FA
 C0 F3 2A CC 5C 00 8F 89 C5 3E 96 8D 50 C5 61 56
 B6 2B CA 3E D5 89 16 6C 51 06 F7 D0 2F 3B E1 5E
 E4 2B C9 44 20 63 F2 BE 16 45 8D 7A 29 6B 4F 08
 49 92 9F 29 43 82 08 7E 5A 38 D4 FF AB 41 E3 71
 23 9E 31 97 0E 74 1E D1 14 37 1F 57 44 A5 AC D2
 34 4E F6 FD BA AD 71 E1 DB 83 D0 91 4B 87 58 FB
 04 87 E9 A6 03 E0 3A A8 B9 72 27 B7 B3 3C 6B 09
 73 2D 82 5A 6D 1A 78 F7 77 95 B0 DA 12 AF EC 20
 30 CD 6E 16 9B F4 24 98 9A 51 2C 0E 22 72 4F 74
 A2 50 A0 D3 B8 01 82 B0 D6 25 E2 CB 07 37 3D 16
 38 6F 52 B4 F6 EE C1 6C 47 67 30 68 0E 5F A2 AB
 59 78 FC EE 55 56 C7 78 85 04 9E 22 C1 4F 19 3F
 E8 AB 04 FE 2F 57 2D D3 B6 A3 D0 F4 57 E2 B0 73
 3B 44 4B 6C 5E 1F EF 8D A8 4B FB 39 91 9D 73 28
 5F 05 E9 63 81 CE 38 9E 87 0E FA B8 EB 90 D4 FC
 EF 09 28 60 34 F2 EC FB 19 D3 B5 D1 74 FB DA 9F
 DC FF FB 40 73 08 70 59 1F B7 BB 09 74 71 CF DB
 A8 C2 2E 49 A8 48 62 14 8E DC FD 5E 71 8C D2 C5
 BF 62 75 11 15 20 2E C3 C4 43 C3 EC C4 94 0A 13
 A4 03 53 B6 60 FE 93 35 83 C7 B1 33 20 3C 55 3F
 40 A8 D6 60 F6 27 CD D3 AE 1B 68 9C 6F 7C 3D 49
 4B 20 05 CA A0 0B 55 60 F5 D3 14 4A 17 2A 4F 22
 39 E6 39 F7 C9 6C 9E A0 66 D7 DA 00 56 CE 97 D2
 0D 11 9D A2 06 62 57 46 35 75 66 10 C6 00 56 C3
 7D 89 82 3B C1 80 14 4F C0 42 75 B3 90 48 EB D8
 14 7B 78 4A 7F D9 B1 51 B4 F6 36 BF DE CD 8D EC
 69 72 12 79 AA E6 64 E9 FD E1 8E 32 77 5B B7 88
 7D C5 3F 2B 92 72 28 6B 10 7F D0 35 BB A3 BB BF
 A7 AA 10 7C 4D 56 69 96 2D D0 A9 97 06 0C E4 BB
 03 54 32 55 9F B8 3C E2 F4 9A 52 66 C6 47 EE EC
 05 1B 3A 19 80 61 38 26 5B 0E 29 BE 13 11 39 94
 D1 EE 4C 98 29 51 23 32 85 93 9C C0 99 7B 7A 09
 FF B8 F3 0F 85 C9 8B 0C BD B9 DC 6C 21 9B 1F 30
 F0 64 83 5D EA 74 B5 3D 94 C3 24 00 33 C0 32 DF
 E9 D0 24 66 D1 61 BD 23 8C 3A B8 12 50 B3 AC 00
 8D 87 CF 0C 18 91 2E 0F B3 AA 90 80 DC FD 22 DA
 7E 08 4F 7F A4 46 78 98 3E 51 9F 18 15 39 BB FE
 14 56 A4 44 DA 58 D3 E3 42 86 13 FE F0 AA 3D 44
 A4 10 6B 73 90 05 FA 55 66 07 B0 0E 92 93 8B C7
 49 96 42 8E 6A 46 1C 4C 92 E6 25 A3 30 11 2A AA
 BD BD 3A E4 D9 32 03 CD 92 27 5D 9E C6 4D 93 0F
 28 0A A2 B6 9C D8 42 2E 4B 50 F8 84 EF 56 2A FD
 D4 FA 40 02 C0 5A 24 2D 8B F5 91 23 E3 04 CC BD
 B2 17 70 E6 C1 28 C0 F1 6E DC B8 AA B7 30 25 26
 40 34 BA EA 75 53 6E 88 A9 72 38 35 FF 36 4C F5
 B9 4E 6A 73 1F 6B D6 A8 1F F9 0B 91 AD BC CF 66
 F8 04 9B 42 33 C2 91 E0 03 EF B8 8B C4 F9 AE 19
 4F 43 15 83 A0 2C F6 39 B5 76 37 51 EA 61 0B 53
 85 0E D9 03 3D F0 21 20 41 0C 07 F4 90 DA FA 46
 F5 B2 0A 4F 94 AB EC 2D C8 07 0A F4 B1 4C 9F E5
 3C 68 F1 30 4A 05 06 DC EF 84 C5 61 75 E4 D2 A3
 A7 F4 2D 64 A5 7A 7D 9C 58 30 32 AF 95 BF 97 B3
 19 AC EF 1E 3B CF 8F 1E 8D 27 9C D7 BE F6 5C AB
 B6 90 5C 25 6B 41 1E 6A 00 36 33 88 05 BA 53 D6
 E4 3C EA BB E8 FB AD F2 84 3B 47 B1 3B B7 B2 89
 72 88 17 BC 1C 6D 17 86 19 C2 A2 A8 FA F7 84 61
 A1 3B E5 7B D3 50 FB D0 DB 3C 62 83 46 0F 4E 75
 C8 93 E2 87 83 A6 F7 66 78 B1 95 A9 89 22 D8 99
 C9 FD 5E 75 B5 F2 B7 D3 97 E4 8F 01 76 F0 D2 D0
 B0 61 67 D4 28 D3 45 7A EF 20 2C 77 1E 12 07 50
 63 BF C0 71 A3 07 95 43 51 42 25 1D BF 6E D4 E1
 84 1B 45 55 80 0C FF 77 C9 1A 6C 02 14 9A D2 FA
 68 F8 74 FA 45 75 D3 54 2B C9 69 BC 5F 6B AF 7C
 8A 24 51 1A F2 E0 77 B4 B5 EB 86 89 21 37 34 D9
 EA 06 B3 96 02 CE 85 66 01 D4 CA 3D 9F E9 3B 20
 1C 84 52 9F 73 D8 7A 87 25 85 16 3C F7 96 AC E5
 79 B2 AC 7D 6E E7 45 82 3A 0A 77 A7 74 9B B1 94
 B9 91 9D A2 62 56 32 AD 91 F8 6B 75 74 8B 7E 87
 1D 12 B2 14 70 5D 9C B2 1F C7 10 05 9F 1F FC 18
 33 F5 67 DA 5A 3F 8E 08 3B AC C4 E4 13 D4 65 EA
 03 E1 21 97 45 11 5D 1F 6D 11 C1 F1 33 38 FB FB
 18 EB 1B 7F 4B 12 5C 69 53 5E 24 7B 57 88 8D AA
 2E 3C 1C DC F7 9E D2 47 37 08 42 F0 5A C0 BD 19
 C4 5A C4 0C E2 28 C4 8B 66 3E DC E2 53 CB 08 85
 86 02 4A 0D DC AA AC 23 56 3C 7E 63 08 0E 41 46
 5F 7B 7E 5E 00 8D F6 48 67 AE E4 83 05 0D DB C0
 A7 2D B2 4F 05 A5 99 13 02 98 3F B5 C8 75 68 3E
 F5 97 9D 4D 24 B6 F0 78 30 84 A8 E5 7A 04 C7 22
 45 B1 7E AB 24 E4 AB 6F 13 88 FE E4 F9 E1 C1 E2
 A7 56 0E 46 80 F4 F9 8E F9 BC ED 56 B0 A6 A3 9E
 AF E6 3D 65 D0 20 C7 DE 71 D3 71 08 6F B3 26 F4
 5F 61 C1 88 AC ED 3B 31 64 48 FE 31 DB 41 12 22
 2F 9B 64 A7 B9 17 21 0C 5C 62 03 2C 3D 7B 19 27
 CA 2F 1F 95 89 02 D1 7B 0B 11 EE EE 3F 06 21 C1
 F7 3C B6 68 11 8B BE 71 01 DB 44 E6 16 5F B5 33
 80 19 8E 71 8F 61 AC 4A 78 0C 17 A4 34 ED CE AB
 56 66 E0 25 4C 04 0F 08 C6 C5 65 9D 97 28 47 70
 FD 3A 32 06 29 AD 08 4D 05 99 CC 25 72 39 D7 EA
 39 95 FB 73 B4 BB A2 F9 6B F1 85 7E 83 4B C7 27
 B3 E3 A0 2F 22 17 E7 9C 6D 64 70 78 17 05 B9 66
 B9 02 DF 06 76 EB 09 DC 2B CF 8A 04 AE E7 BE 39
 12 76 E3 DC 79 8A 60 77 69 4E 45 08 73 25 42 FE
 7C 30 C8 2F E8 F4 00 85 4A A4 C0 88 68 1F 40 B1
 90 E0 86 78 56 B7 70 33 2C A3 EE 41 5A BE FE A2
 78 D5 BC A6 7E 2A 37 63 EB A6 44 E4 AC FF 01 0D
 09 94 D6 70 DC A7 6C F9 62 78 D3 DD 4A 7E F0 E0
 14 88 5C 25 59 35 A2 FC 11 A6 73 B6 AA BC 05 86
 9C 20 36 ED 26 22 93 9A 1D FE DE 8E 70 B9 AE 81
 C0 0D E4 15 E1 78 1C 89 1B DA 28 40 6C 44 93 30
 9D A3 FB E2 86 B6 D5 DF 9C 7F 7A E2 EB CC 3B B7
 48 22 52 6F F7 F9 A3 C0 B5 25 87 37 F7 76 4D DE
 A0 2E C5 E3 5C 27 6D A1 07 C7 74 AB 2F A0 A9 A6
 FE 27 7D 8D 24 01 96 5E 0A 9E 3A 00 72 A6 2C 0C
 84 B4 C4 F3 BB 2C 64 86 57 D4 D5 8E 8B 7B 25 F5
 93 A3 38 7D 53 5D 72 90 FB E0 D7 28 F9 B5 4E 60
 26 85 02 29 E6 29 09 39 79 AB 9F 50 2A 60 3C E0
 E5 B9 73 79 C4 E9 2B FE B4 84 8A D2 B5 53 B2 84
 D5 07 78 0A 41 25 C0 62 53 F3 BF E3 3D 96 85 9E
 7B 74 1D 8B 5A 8A 25 31 21 7F B0 B0 19 DC 8E E8
 EB D8 A4 FE 41 15 B6 B5 E2 50 35 F5 C2 8E C4 F9
 68 11 AA 72 2A 0A 87 43 7E 63 F0 B5 04 1B 6D 77
 62 8A E5 03 6F BB B7 3A 42 CB C2 25 69 A9 86 62
 8F B5 DC C3 65 10 38 86 9F 89 A8 8E 18 A4 E3 EB
 25 63 F8 53 80 A4 18 08 A3 B5 28 1C 97 29 EE 63
 D2 67 D6 2B 3C 5D 5F 3E B2 E8 96 49 10 A4 7A C0
 EC F5 08 D5 71 36 F5 82 29 D1 F8 9B 32 04 FB 09
 CB FF 8D A0 37 6A B9 95 60 21 80 14 C0 2B 41 35
 2F F6 14 21 32 D3 ED 05 B7 7C FC 42 88 ED 5B 88
 33 A2 64 00 13 07 A6 27 C7 CA EA 07 13 26 C8 07
 73 FA 99 86 B9 18 D0 35 D7 9D D2 A6 E2 9B 54 BF
 F5 8E D1 41 AA 8C 73 26 EC AE F1 C7 53 FC 2C A7
 FF 0E 75 9F A2 3B 7A 27 EE 47 3D 8F B5 CD CF 8C
 3D A2 4D 7B 99 8F D6 48 33 7B 97 BC C6 A2 82 C4
 3F F1 3D D3 1F 4D FD A0 12 3E 95 66 48 13 6B 56
 00 47 CD BF C8 7E A5 2C 70 91 A9 E6 3D A2 05 C7
 9A 4C 67 AC 27 54 06 E6 36 1E 65 1B FE D8 78 44
 DC 42 17 47 27 03 0A EF 71 EA 12 2D C4 47 73 E5
 2E FD 38 21 19 40 76 78 19 CF 7C 93 EE 07 FE 84
 31 6B 4F EC 6A 73 22 E9 64 BA C1 D5 6A 8A 39 01
 F5 C4 D4 A2 63 71 80 CF 23 E8 37 19 F7 6F 45 CD
 9A 1C 55 BF 5B 06 34 39 C9 5F 53 86 2A 6F 12 75
 E3 54 4D 63 87 D1 C5 BC 9D 53 AA E1 52 B9 D4 22
 2F 7E 27 E1 F1 51 87 8D A0 6B 7C B7 F4 1D FC 7E
 A2 5F 3E 36 4F 7E 62 E3 78 98 F4 FA 55 8C 13 6E
 9E 19 EE BE 42 0D FA CA F2 7F 6B 24 8D 14 51 D1
 D5 7D 66 D1 84 6E EC 33 72 75 AF D3 52 23 15 14
 09 B1 85 C1 82 8F F3 51 04 C5 2F FA 77 BE BD BA
 F6 36 A6 36 AB E8 B6 95 AB F7 DE 5B 53 83 53 89
 06 C8 29 D4 FF AA 00 E8 C0 EB F5 46 88 59 BF 25
 F5 83 EE A5 9D BB 74 B7 93 3E 8D E7 1B 7D DC 8A
 C0 45 BA C2 47 99 31 1B EC FF C1 A5 5C 07 CA D2
 78 00 00 05 6A FD 1D 18 B1 FB 44 E6 47 C1 92 44
 38 F7 43 FE 97 43 0D B5 DD 94 53 DF 8C BD 8E F1
 3F 72 87 0C 26 24 DF E6 7C 3B 5D 53 BC 21 20 C3
 4B 74 C6 F8 0E 64 92 8A 96 EF 6B AA 03 6D E9 20
 17 1C B1 A2 9F E8 C1 6A 9A 1B 6F E8 35 DB FF 64
 C8 FD F6 9B 09 AF 4A 37 3B 2D 1E 46 37 FD 16 B5
 EC 18 5E 49 07 87 FD D5 7E 27 98 02 C1 99 C8 88
 BE 82 38 1E 53 E7 2D 23 54 31 FB 85 CA 71 27 A0
 A5 A6 B1 9F 5B CE DC 42 49 AF C1 32 85 13 B5 20
 91 DC AF 9A 94 AF ED 5A 59 B2 9B 4C 50 62 F1 77
 95 0C EE 9E 41 B9 E5 41 E8 26 FD 63 4A 90 45 DD
 66 DC F7 72 0A 42 BF 16 41 57 AE 27 28 60 6A E8
 33 FC 21 A9 53 2D 15 7F DD 59 ED 83 D8 91 B9 4A
 46 37 49 06 6E 7A FA D7 C1 A2 0F 15 90 F8 33 80
 3F 4D 96 6C 3E 90 59 2A 8A 04 A4 89 6A DC 0F 80
 A5 D7 A1 7C E2 CA 46 32 D7 03 06 E1 1A 0D 68 B2
 78 4D 18 C4 7F 4D 7A 58 84 91 65 A2 34 76 D1 44
 61 15 55 1D BF 4C CE A6 4E 73 5D B0 6E 1B B2 C8
 6C 6A A2 9B E7 85 45 02 1B 74 23 E9 83 19 A8 FA
 48 53 C2 5D FC B0 62 45 29 77 AE 2B 59 E6 5D 71
 CA E6 3C B5 EC C4 E7 9A EB 36 48 1F A3 E0 C2 10
 BD C3 C9 76 B2 49 DE 9C B5 EC 5F FD 0D B1 14 98
 F3 FB 21 D9 01 2F AA 0C 2B 72 A9 ED C2 37 51 1E
 E0 C6 5C B0 F0 25 B2 67 C6 24 3A 6C 4D 42 B0 8F
 C7 49 4E 46 5F BC A0 F2 13 9F 0E A7 30 CB E0 60
 32 F8 91 F7 8A 9C 0F 32 29 F9 6D 9E 0A 65 06 FD
 D8 71 6D 5D 12 8E 2F 94 6A 91 41 09 64 D1 93 99
 17 B3 8E A4 94 37 F7 D3 BA 81 FB 75 46 82 23 CD
 3E D4 6E 79 0C 2C 47 40 70 E3 8B F4 9E 5A DA FB
 ED 40 FA 6A DC 3F B9 CB F8 E7 29 79 C4 97 F7 89
 08 23 EB 7E 07 E5 47 0B 4C 36 F5 93 CF D6 50 FF
 72 74 98 49 7A 0F C7 C1 8F AD 43 8C 7E A8 A1 AA
 BB AF 75 6D D8 79 0F D3 6E DD FD 5C 6D 08 C1 36
 EE 7C 77 53 7A 07 CC 24 BC 32 82 C9 4C AE 86 45
 FE 95 56 48 80 9B 1B 2B 3B 44 94 FE 36 10 97 C3
 33 46 AC F8 90 B4 5E 71 69 62 75 34 24 1E 33 70
 27 E8 97 5F 91 60 9F 61 AB 00 EB BF EC 8B E2 0E
 B9 19 54 16 2E 38 E7 69 67 57 71 9D 07 5C 0F 37
 55 94 3D B4 B1 55 CE BA CC BD A8 7B 22 BD DE 01
 4A 8B BF 5E 67 0D A7 2C B6 E2 A9 7F 37 C8 49 3F
 47 DC 7F A2 F2 51 7E 28 71 52 52 27 CE BE D7 8E
 08 C9 72 4E C6 69 08 80 54 01 46 C5 63 1D 47 48
 58 87 0F 83 0E 92 F4 09 73 6D FE EB CB 0F 18 1D
 C6 A7 A4 31 E2 19 21 6A 9D 56 F7 B1 DB 21 6E A8
 F4 1A 66 51 6C 4D 94 29 86 3D F5 71 D2 07 10 1A
 78 B6 7B 07 63 8E 0B FC B8 28 EB C1 07 99 A5 4F
 60 49 10 A1 59 4D 13 8A 45 74 AD C0 AB BB DC 55
 F8 05 B8 6B E1 67 4F AC 03 3A 48 D6 CE 1D 76 43
 B1 2D F4 70 94 38 78 A9 CC 38 48 E5 99 8F 12 FE
 EC 1C 96 9D 74 AC C6 33 91 92 02 56 57 05 72 38
 B2 1C 1D 6D 91 4D 49 74 F2 96 C1 E4 5B 20 5A 05
 12 AA 5E 7E AF 6E 59 5C DF 6B 1C A7 6E F6 36 E9
 B3 10 D2 17 16 FC D1 F9 8F 74 C7 0C 6C 61 2C DB
 A0 22 F0 5F 02 84 A8 BF 08 CD 4B 5E E2 BE 3B B1
 48 BE 45 44 B6 4D 1F DE C4 0F EB C0 4B 00 AE 01
 C6 8F 3E EE F2 8E FF 3B 87 78 03 09 D4 0D C3 29
 5D 90 44 0B 40 0B 7D 5C F1 9A 6F 91 A0 8D A2 CD
 A2 21 10 FD A2 A9 D6 96 D9 A4 EB AC 48 00 AF E1
 5C AF 5F 1B 0C CF CF 10 A9 20 08 88 17 A3 6A ED
 61 82 73 89 C6 5D 75 DA 91 D3 A1 CD BE 1A CA 26
 6F 4A 3A C5 FF 47 44 11 61 13 58 62 4A A5 BB E6
 E4 ED 5F 44 EF B5 B5 54 20 84 9E ED F3 87 72 9D
 03 59 03 39 08 1A EF F5 26 CE A0 98 5D A3 21 A5
 4C B3 A3 10 BC 6E 67 3A 25 79 F8 B2 90 99 F4 CE
 D3 D3 39 15 CB FD D6 2A 5D 51 F2 50 9E AE C5 E9
 7C 93 0B 1C 85 80 15 9B 71 21 5A 63 72 56 F8 49
 60 7A A3 D7 3C 1E 48 C6 EF 13 91 86 C2 AB 1F 9E
 56 62 20 FD D6 15 BB 2E DF 26 10 EF 62 D2 E5 3A
 36 41 4B CB E7 82 DB 50 F9 5A 1C 4A 26 5F 89 81
 4F EC 2A 79 04 BD 7F D2 6A A3 03 7B 21 D4 48 B5
 D8 09 53 00 66 EC 4B A1 A8 B4 3F 8E 45 7B EF 74
 A8 0D E5 87 86 37 CF A9 D0 FA 3A 98 4E 68 8F 65
 37 9C 98 C5 AE 86 0B 1C E8 BA 88 E3 A5 BA 91 DB
 CC 58 BF 06 24 E9 E8 A2 22 2C 22 7B 03 1D 74 93
 54 7C 0E 6A AE 5B 43 D2 51 F2 59 C2 F5 B2 98 8C
 2C 1C E9 81 D8 47 BB EB 96 03 D8 A9 B8 F1 1C E8
 8B 2C 9F 99 BD AE B6 03 84 E4 2E 08 62 F2 8C C3
 65 F0 3D 4C B0 97 18 10 0F 33 1F E0 92 AD EF 45
 66 7F 74 CB 77 01 08 59 B7 44 C2 62 9D 7F 02 5C
 A6 58 4A B8 19 71 CE 61 4A 63 B2 85 8E 3A 98 24
 C1 71 A2 ED 16 51 94 8F 52 E7 9D 15 DC 11 62 22
 2C DE 7B 20 1A 72 2D 13 F9 AE A9 94 F8 ED 6F 27
 42 60 E2 45 04 AE 8F 6E 87 62 91 3B 7E 15 F8 0C
 24 A9 A3 57 85 5E 35 24 5C 06 7C CE 79 5F 3F EC
 DF 90 CE 88 A9 3A 49 F6 50 CB 18 DC 34 2C B2 91
 99 59 13 2C C1 D7 D6 BE DE BE 16 D3 A0 C8 33 76
 F5 E3 7F BD C9 0B 90 EA 27 01 8B 7D 40 92 A6 12
 4F C6 13 DF 8E 5D 02 FB 13 35 C5 25 38 9E F6 BD
 1B C1 64 36 D2 40 32 19 C8 0E 85 10 02 63 A4 0C
 D1 99 56 07 B5 DC F3 1F A9 C2 01 D0 2F AD 14 9A
 57 81 7A E7 73 9A 41 76 E9 49 49 41 A1 4C AD 50
 7B 2D A3 83 B4 EA D9 EA AF 93 BF 17 2B 1A F6 A4
 D1 65 83 8D E6 23 D4 BC 86 BF 0F FD 55 7C FA 4C
 D0 F1 86 5C FC 65 32 9A 2A 28 05 F5 59 95 07 F2
 BD 7E 7B D6 F5 70 A6 02 89 0D F3 CA F8 CC 2C 4B
 C1 E2 72 0C D3 EF 9D D2 A3 C8 1B 26 A1 87 10 65
 F8 4C 3C D7 10 FF AD 0D 8C 1D 12 86 06 64 0C B9
 C9 29 E7 A3 A1 5B 55 32 D7 F6 74 38 E2 38 77 D9
 17 CD C8 93 66 BF B6 5A E7 4E 75 0F 3A 4A F7 7C
 0F 6F 55 96 E5 CF 00 D3 7B FC 73 46 9B 7B 5D 8B
 56 14 45 79 1F 9E 2A 36 38 57 2D 9B C1 7E 8E 62
 0C A7 28 72 7D 81 BB 2A F1 1C EF 01 24 BC 39 73
 78 56 C7 1D C6 E4 69 92 90 12 52 97 E6 0E E6 96
 27 D4 FA A0 64 55 DF 16 60 19 16 E9 E8 1B 3E 67
 2A 2B 64 E6 A1 47 1F 7D 1B E1 25 30 0B 70 33 1F
 E4 7B 3D 7B D8 C4 CF D0 D1 11 B0 E6 20 BD 71 C6
 0A D1 2C 21 4D B1 9E AA E1 C2 93 82 E9 1F 25 72
 AE 4D 97 F7 3E 79 49 7D 3F 66 D9 59 52 9D 36 79
 C7 A1 DE ED 68 A4 AD AB B0 D0 DC 0D 19 B9 BA 53
 30 B8 C5 5B 72 69 28 98 E1 78 A8 48 61 84 14 27
 6C 60 41 63 B8 84 3D 86 8A AE 57 2F 10 8C 22 B8
 D2 F2 CE D1 BF 62 62 FA 4F 1F 4E C0 A8 1F C8 CA
 8F 32 ED 75 EC FE 6A 9E DD 33 8F 3A 66 57 80 FD
 FD 7F 58 6B 70 E0 A2 62 DC 98 82 46 16 3C 5D 0E
 08 E1 96 B2 84 3B 16 18 83 05 AC D0 1D 85 A8 DB
 B4 8D E4 BA 29 D7 A8 B8 67 C0 7B 47 C6 AE ED 22
 A2 05 81 56 D7 5C 13 27 DB 0B C2 2E 0B 23 CB 5F
 88 A9 A9 CE 10 00 11 CE 7E B9 5F 27 0A 72 B2 E1
 13 84 85 F5 6D 6D 5E D9 68 6C 34 0C BB 00 13 3C
 5B 2E 71 A9 1A 63 EA F2 D5 D8 5F BD 0B 80 B6 49
 73 2B E7 79 08 F2 AE FE CF C2 01 B8 2C 44 46 03
 17 9C FE EF 34 77 16 B4 70 51 4B C5 72 F9 71 89
 45 55 6D 17 20 F2 CA 51 9E EE 9E 7C AD 8A 61 93
 07 3E 1A 01 91 42 E0 63 9D 46 8F 65 07 F2 DB 1E
 BD 56 04 21 3F 5F 3E F8 F8 8B EF 79 2A 93 2B 85
 40 8A 66 A0 23 26 3E 27 6D 04 D4 65 FD 05 1C 1B
 31 8D D0 D2 14 CC D3 F1 AC 62 B3 A3 AB 62 8B 03
 FF 51 E1 DD C6 99 DA 8B 79 06 39 63 6A 97 F8 D7
 53 CE 25 20 13 FA 41 53 3F BB 19 46 94 D9 B4 D9
 78 BE BF 89 0F C4 0B 26 6D 31 ED B4 D0 C7 B0 18
 3A AC FB B9 DC 23 1A 4B 63 B9 E0 57 FF 31 69 C4
 77 07 E2 47 F6 61 12 C7 55 29 67 6F 13 DE 92 91
 D0 A6 30 92 14 A2 76 10 60 DB A1 D1 BF 89 92 60
 CC 18 0E F1 A6 56 61 F5 4A E3 9D 4F 38 CC 65 D3
 4A 1F CF F5 31 C0 1E 4A BE D5 B0 F6 1D C8 0D 94
 B9 14 87 EA 98 A5 97 D5 75 1D 3F 3E 97 EF 6A D8
 8C 37 E4 4C EC 15 07 C8 E3 CD 0A 56 19 18 25 3C
 87 DB 35 54 A5 BA 75 DA 84 6C 8E 51 20 5C BA BB
 01 8B 5C 89 A5 A3 A3 91 8B 7E 94 DA 6C B6 F1 F1
 97 18 2E A4 A0 D4 EA 03 D0 60 91 42 3B 76 E0 89
 DA 9C AD 03 AB 1D 64 CC 01 33 82 F7 58 B5 B3 71
 C7 98 53 0B CB 1F 02 57 AB 7F DE 90 E8 48 31 D7
 65 08 A7 DF 43 B4 D4 7B 98 36 F2 78 E7 89 AB 13
 32 1E F7 6A 70 FC 94 A1 43 2A D2 38 DE F7 7D DA
 94 80 7C 99 59 E7 E8 ED CC D5 23 08 AA CF B1 D4
 60 B5 CA 78 A9 88 E6 42 4A 07 6C 52 B7 7A ED 8A
 6E 39 BB A0 5F 7C 45 0F 75 9B 56 56 5F 01 67 68
 8A A1 9C 56 9D 08 A4 7E 6D 81 8B D5 E6 61 E9 1B
 70 75 D5 0E 8B 9C 32 3A 62 33 B1 48 14 F8 F2 79
 8E B1 EA 6B 34 0D 57 6A 2B 6F 60 A9 16 47 A5 31
 0A EB 8D 6B 74 6B CF C2 3D C1 0A 50 1A DC 1B B4
 45 BE 83 B9 B7 83 50 83 C1 69 14 F4 D0 00 71 20
 62 6D D1 1F 89 B5 B3 6C 5F 7B 90 55 C3 1A 8F E5
 4F 1B 08 79 E3 2C C2 43 8C E1 CB 97 EB 34 85 00
 5A 32 37 57 A9 D0 2F F5 50 44 FB 53 B3 1A 5C 0D
 EF A6 34 D8 B9 C6 14 FF 4D 61 7D 00 7C 39 A0 5C
 9A 31 19 95 07 50 86 DC 90 A3 99 83 6B DD DE 80
 C9 76 86 66 58 2C 50 76 7E 1F 24 AB CA 58 7E 1F
 34 B1 6A 68 46 66 51 F1 25 EB 0F 30 E7 8E A2 14
 43 83 1F D6 6B 06 5C 88 FF 6E CC D8 4D FF B4 0D
 AC 27 1A A4 75 4D BA BC 6F 7C 51 E3 13 AD B6 D6
 E2 CF 17 B6 E3 B4 9F 46 AB AB 0F 77 9F AC B6 02
 B9 61 37 74 79 A3 CD 4C E7 DB 36 B8 FB 30 7D 5B
 77 2B 6D 8D 34 0C 17 41 26 3C 51 B5 C2 4D 4F 49
 AD D8 1C E0 C0 67 E7 B7 56 B0 CE 64 25 5B AA 1C
 FA 80 8E 7D D7 78 7F 06 1B 5E 48 50 2F 07 B6 A9
 1F 86 0E 88 09 F5 77 A7 29 84 DC B5 39 4D 4F D6
 E6 A1 A0 E3 96 2A 4F DD BA FB C4 A0 97 0A 99 EB
 1C E5 79 02 EC 96 4C 3C 84 FF 55 B0 05 A2 B2 BA
 96 12 EA 04 54 91 FB DD E7 16 49 CE 32 B3 0D 3F
 45 A4 6A 49 85 BC 4F DC 48 CA 1B F8 1D F7 8F B6
 84 20 98 1F C5 FC BA 12 77 F1 1E 51 8B E3 C6 22
 51 3E F0 83 81 DD C8 2A 7F DB 9B 82 78 13 93 4F
 62 A2 33 A5 C3 14 86 88 E5 EB 29 94 E0 D9 4F FB
 9B 28 46 BC FA AF 1B 05 4A 78 9A EF 1C 72 5A 7D
 95 57 27 9D 8F 38 A8 38 9E 21 2D 0D 92 9A 44 05
 C0 FB 8D 02 41 F8 40 28 A8 74 CB 83 31 0C A2 B3
 53 08 1D E7 F8 4A 94 B5 2E 99 A1 D8 55 C3 BE 92
 7D E9 7C 97 4D 03 59 A3 8B 43 6A 7E EA 1B 63 7A
 C9 3B 81 E5 49 68 83 3F 3F ED 47 DF 06 1E 7F 91
 8B C9 28 97 39 B0 79 10 B2 4A 54 55 98 F8 5D 39
 8A 7D 08 43 A8 21 8C AF 5A E6 1C 42 DB 6A BD 7A
 A6 56 2A D9 30 B2 C9 B9 E9 D9 2D 8A 69 17 B8 CA
 76 9B 5D CC F3 08 AB 11 48 8E 1A 0A 12 BF 4F 76
 3C 2B 61 7A 09 D9 D3 F7 03 7A 48 68 78 D0 DD 44
 7D 67 3C 12 BD EF 95 CC E6 70 CA CF 40 8F F2 7F
 BA C1 04 64 29 32 FE 7F 19 60 59 A7 1E 18 07 BF
 B3 93 5B 51 19 10 98 72 AA 6D 28 44 FF EC 9F E1
 47 F6 51 33 79 0B 82 EB 2D DE E5 DD CF 25 31 65
 62 21 FE 1D 5B 26 66 D8 F0 EB F2 E0 C0 8A 00 9F
 C2 D1 A4 4B CC 8B D4 56 03 CF A2 D6 D2 90 3E 72
 32 7E 56 B5 66 EB 21 FB B4 B6 97 2E AB FE 84 BC
 3E A3 9A 19 C0 8A 8E 00 36 28 39 85 3B 6E D1 F6
 3F 74 8B 36 BE BD 0D A2 37 B1 17 D5 83 E4 0B B1
 78 6F 58 F4 D2 50 0E 4F 22 F6 02 E0 F5 52 B8 A6
 4C 0B B7 98 3A 2A 61 9A BA 64 8F 3B ED B6 36 79
 25 0C 74 7A 5C 10 EE 6D E9 11 2B AB BA 4A BF EF
 78 77 5D 25 BF F0 89 67 57 89 59 89 9F DB D8 6C
 A8 8C 86 26 51 CE D5 00 E4 BA D0 3E 38 E5 E9 0D
 F8 03 99 4E 1B 79 6F 32 24 6D 43 92 67 F2 F1 32
 1A 76 A3 3C 5D 5C 33 77 04 6F 2C 76 73 27 4D 9E
 67 EF E5 CF 8D 43 75 ED 85 D1 08 37 62 92 77 C7
 4F 3D E8 7B D1 8E 12 09 02 E5 D5 95 37 85 AA 89
 82 FB 9A AF 59 EF E5 74 B3 C6 EE CF A6 00 F6 DB
 DC A4 89 22 8D F2 A8 45 43 CA 80 8A B4 06 EE 0A
 0A 67 19 8D 3D 1D 78 BF E0 1E 9F 59 00 D0 42 99
 93 71 05 6D 91 3F 1A A7 F6 DD D4 2E 5A 02 1A FE
 0C 9C 1E 1A EA 14 80 8D DD 31 A1 C6 3C 3C C1 3C
 76 37 07 D3 49 82 26 20 08 3D DB 5F BD 46 89 26
 CD F9 77 9F 28 0C 39 19 10 A0 4C D3 6A 8A 7B BF
 82 7A 8A A7 03 5E C5 87 3A 38 F2 6B 88 D8 DA AF
 4D 7C 77 EA 42 12 70 A4 1A 03 01 9D 22 51 7D E0
 86 F2 AC DC AD 0F 27 4C 49 BB 44 DE 3F D2 11 EF
 BD 97 A9 70 47 3C 5B 2C 35 98 92 A9 D0 50 AC F6
 80 9C 94 F3 E9 41 06 A4 C2 8C 4E AE F2 90 F5 37
 EA B2 4A A2 FB 98 17 AC BF E6 02 71 B5 B3 F1 88
 24 02 80 6D 42 5A 4F 4C F8 DC 25 B2 C8 04 81 46
 56 60 17 0F 03 3D A3 D9 9F 69 F9 A2 13 3C 2A A2
 63 E7 C6 6B E2 D6 EC B9 DE EF 70 B5 A3 48 9E E4
 F6 32 AD E6 51 E6 A1 81 AC 67 99 B3 0F B5 AE FA
 9C 1C D7 A9 91 1C DC 11 5C DE 5F EE 4C C2 48 1C
 A5 F1 8E 60 52 63 E2 DA 25 F6 64 6D 0A 61 51 84
 7D 39 54 CC 38 2F E4 0A 43 A9 AC 87 DA A9 FA 2D
 13 A0 09 41 21 CB CD 31 AE 8A D6 F4 71 0F 0D F3
 A9 E1 14 15 81 73 28 82 B4 FB 71 69 1E 7D 30 42
 C7 3F 51 2B 65 5F 06 53 EA 18 36 92 4D AD B4 BB
 AB 7E CC 62 F4 CE 87 BB E2 05 F4 5A C1 41 9B D5
 36 55 88 D0 46 BD 19 AE 4D 46 70 44 5D 8D 0B 27
 33 11 13 98 67 F5 25 76 DD 58 FE 46 CA F2 33 0C
 20 B1 ED 43 DD 2E 81 B3 D8 15 FC 50 87 29 9D 61
 48 96 6C 2F 31 15 15 7C F5 D7 C5 C0 39 FC 60 29
 AA FD 58 F3 C5 C3 3B 9F CB 50 4B D4 B3 86 C8 24
 AC E9 F4 59 1E 24 AB D7 D9 98 91 05 90 74 CD F2
 CA E3 21 53 DE 40 75 3E D5 87 89 B7 29 E7 05 1E
 3A C7 4D C0 58 A9 A4 BB 13 D0 77 CC 6F 3C 6F E6
 13 3B 59 1B 4C D8 7A 8B CE C3 10 12 2D 9C C2 74
 E7 6B 6C FF 26 38 4D E8 AF 19 0E 9A CC D5 DC BE
 2E B9 23 09 45 1D C6 F0 25 D9 3B EF 13 8A 00 6C
 1B 27 9B 5F 18 A0 35 19 A8 1E 3C F1 5E EF 80 D4
 1A 1D 5D B4 79 32 D4 01 4E D6 16 DE A2 B0 F0 43
 56 50 AB 86 FC 39 8C AC DE 68 A1 1C C5 1C B4 F8
 D4 37 4C 1A 0C 30 A6 AA 08 96 FA 7A F1 60 60 0B
 7C 25 4E 3A 1D 9E BE B1 7B BD C7 41 A4 62 EE 6D
 71 12 81 F4 E1 77 52 1A 2B 4D 5B 48 D9 94 23 7C
 73 24 A1 A4 DE 4D FD A4 A2 8E 8E FB 61 55 E8 29
 33 8C 6C C0 E3 14 27 91 C6 2E 8B 73 11 7E D7 92
 A6 67 A2 C0 54 84 28 3C A4 6F CF 05 7D CF E1 55
 44 09 F2 80 D7 F9 44 77 3D 76 EE 25 3D 4C D9 9D
 61 4A 57 F1 85 5E F5 4E E3 B5 E4 D2 5C 91 09 47
 D8 25 8C B5 1E 6D 57 23 C6 8A AE B4 70 85 D0 48
 0E E5 72 BE 11 03 52 47 BD 92 A9 B5 BC 1D 91 F2
 15 BA EC C0 05 6E CE 76 A2 14 F8 3B CE 29 37 C3
 4C 72 28 2A 36 4C C4 F3 19 37 71 61 22 99 E1 23
 0D C5 60 B6 A3 4A FF 3E C2 E6 79 EE 32 8C E9 E4
 12 88 39 F8 4C 86 ED 7F 45 10 B0 05 66 36 31 84
 66 1D 2B B8 51 A9 E8 A4 84 B8 88 92 77 CA 61 3D
 DF F7 AA 35 4A FB 91 76 B0 19 56 DB AA A8 B2 48
 B5 1E 71 9F 21 AB 40 CD C2 BE C4 FE E9 91 DB 7A
 B7 F0 C7 E5 61 7E 97 98 BC EF C7 E3 34 04 25 CE
 C6 F8 4E F8 C4 CF 0D 09 23 4B 83 C6 40 C8 1B 42
 DC CD E8 68 86 02 09 CC 91 DB 21 AE A1 BC 3C 22
 72 3C E1 58 A3 7A DF 5F E3 67 EB CD 35 47 FB CD
 9E 40 81 E4 42 53 43 53 70 BF 54 8E CB C1 3E 33
 C7 44 F8 7B BC 51 74 0C FE 2A CF C0 3F 49 0E 8E
 BF 9C 47 26 A4 3D 67 CD 06 37 66 89 10 58 BD 5E
 8C 29 53 6E 7A 26 C9 4D 32 F5 B0 B0 AB 6F 0E 44
 94 2A 11 BC A6 77 A8 FC 2A C1 D0 F9 EF 35 6D 3C
 5B BA C1 AA A2 38 85 C2 C2 23 75 FC BE 87 DA 2A
 82 34 3D 6F 4F 01 E9 68 2B 17 66 6A F6 7A C0 0D
 2A C6 2A 5F FA ED DE CD 60 F3 E3 41 3A 76 51 0F
 2C 42 97 0A 91 50 B9 01 DF E2 85 EF 84 A0 EF 69
 6A 8A 84 38 D4 96 0B 1D AB DA B9 D8 95 35 7B AA
 3D 87 EB 24 23 1F DF 93 3C 20 95 5C EC 06 CC 6F
 43 4F 14 CD AF 3C 62 43 D6 F9 7F 82 95 99 37 08
 E8 34 61 AB B3 5A 68 10 53 5D 32 13 E4 71 02 2F
 13 13 7E 9B C5 7B D6 DC 54 9E BB D9 E6 FA 0F 8F
 2C D1 4A BA 27 0F F3 E9 63 0B 79 77 8B B3 52 31
 05 61 B0 C3 B1 A4 96 0E 35 7E 78 93 A4 B6 C9 A1
 66 F7 9B 41 54 F3 18 20 F8 27 C5 23 FF 44 68 FF
 18 74 7C CB 0E 74 91 84 1C 80 D8 0A B2 79 C7 C9
 5F 1E 5C 6D 8A 90 25 E8 A8 7E AC A6 46 AE A7 5F
 7E 20 8D CA 7B 08 11 D9 61 DE B8 73 9A 2C 70 B8
 BC 24 C7 C5 16 6B 01 19 B2 94 E9 4B 1B D4 5A 47
 54 8B 25 2E 70 1F 08 31 67 49 2B FA 1C 69 33 B7
 8C 12 1C C7 81 CD E8 6C 7A 1F 4F 99 0A 89 D7 A9
 72 77 EE C8 63 50 C3 E7 1D 39 07 75 17 7D 2A 4D
 A7 E4 4C 05 77 5F C3 8D C6 15 A5 49 9D 10 4A 63
 FD 19 02 D3 4A D5 9B A0 DF 31 55 D6 FD 05 96 D1
 B5 78 4F 73 9A 3B 90 24 86 EB 50 AE 36 85 7C B4
 F6 4D D8 48 E2 34 EB 0C F6 02 78 6C F2 32 E0 8A
 5D 09 F2 22 10 38 30 78 0B 59 00 BA 5D 98 97 DA
 95 C1 10 19 80 0A 1A CA 61 A6 D2 03 8E 83 A8 A1
 2B 48 A2 77 77 7D 3D EB 27 60 C4 D5 8C 25 EE 51
 3D 0B 73 BB CF A9 EC AF 09 0F FE 2A 6E A7 91 47
 02 81 DC 24 EB 6A 72 D1 91 BD 0A 05 8F 1B 94 EE
 28 84 94 1A 09 E8 9C 2D 9C EE 1F 3A 07 01 2E DD
 31 C6 EC 69 39 50 66 4B 0C 77 DB 06 0C 94 7E 43
 DB 89 0C BD E2 74 5C D2 73 EC 60 D6 42 4A E2 29
 15 DD F2 DD D2 F8 13 E9 B1 A6 C9 B3 95 CB 5C 9D
 D1 B1 C7 31 FA 14 AF D6 75 FD BF E8 CB 4E 7E 23
 EE F2 89 1B 09 B0 F6 20 B6 53 6A C6 A8 08 9B 8C
 91 B2 62 29 64 F9 26 83 F0 E8 BC 26 FA C6 26 33
 0C FC 72 7B B4 5F 6E C2 C9 49 05 91 7D F8 87 E2
 F9 58 15 E6 1A E0 BC 8E 6A 1C A6 4E 3D 46 9A 20
 66 38 48 92 EF C3 9C 87 2E 5D 68 BF 75 63 5B 43
 67 6A 2C EA DB E5 04 00 C6 D6 63 3D 7C 34 57 C1
 68 D6 DB C8 DB 04 71 DC DD 0C 0C 4B 31 05 12 7B
 5B 80 93 75 81 85 B3 4F 7C CE 5F 5D 11 BA D3 E6
 CB BB EC 9A F2 90 24 F6 4B D4 E0 19 58 80 37 F0
 67 87 A7 CB A3 06 1F D9 EF D9 C6 37 CB EB 20 9E
 08 50 D9 06 B1 24 89 B1 F1 E5 65 07 E7 ED 6D E3
 AE 32 DB AE C6 83 A7 4B A7 89 80 BB 53 BF EC 4E
 F1 A2 73 E3 95 DE 08 AB A0 8D BC 12 8D A6 D2 E5
 2F 48 D3 77 73 02 5C 29 82 44 CB B4 94 12 95 14
 A5 72 1A F0 16 60 34 9B FB 0C 0C EB 81 60 AE 5F
 D4 81 BA 9B F3 13 FE 84 96 33 BF 98 72 C2 57 6B
 3C CA F9 9E E6 43 10 7F 73 A0 39 E9 BE AB B7 9A
 29 66 3E 11 D7 7B DE B5 45 07 E1 B5 82 BC 18 B5
 AE C4 9B 98 10 21 E8 AC D7 88 F1 FC 6F AE 36 A0
 C2 AF 40 5B CA 03 4A EB DD 5A 86 FA C0 29 F6 FF
 C1 2B 64 60 F1 1B C6 77 52 62 E7 7A 87 5D 69 6E
 95 0B 15 5B 4D F1 A9 E1 E6 DC 37 F0 61 3C 7F 8C
 95 97 30 BD A7 92 1F 45 F7 20 9F C8 2C F1 5B 3C
 E4 81 3F D9 8E 49 A1 04 EE CC 31 C3 11 69 EB 04
 2D 53 5A EE 74 F6 D0 E3 29 5D 08 99 CB 86 F3 81
 C3 81 3F 9C 7C A1 DC 0F C3 38 DC 33 FC FF 13 3E
 29 80 BF EE 24 D1 18 81 48 DF 58 90 1A 10 90 94
 2D BE 73 58 58 41 F1 55 57 91 75 2B C6 C5 7F F9
 23 C1 14 3F B3 B0 9C 25 E7 FD C5 63 71 D5 D9 2E
 41 3B 1F 45 B4 0D 1D 74 3D 75 3D 3B 71 72 E0 5F
 CE 70 38 19 DC DB 08 02 BC 46 5B A9 26 04 E9 7B
 4D 28 D4 7B 75 15 B8 A8 22 FA F6 3A FD 95 75 CC
 53 DF 82 EF 9C 93 C9 72 10 7B C1 61 38 C2 40 57
 76 74 40 74 C2 AB DC 0E 05 96 23 41 7C E3 91 DE
 46 AA 07 67 59 41 E1 87 EB 08 A1 8E C5 8E 43 70
 68 B4 B9 01 2F 44 84 26 71 E4 50 87 96 60 F2 98
 D4 52 4A C6 24 96 89 75 DE B7 58 1C 97 C3 1E E3
 1C 33 1D 2A 75 3C D3 79 19 2C 13 89 48 C3 2A 2B
 EC D3 1D 97 06 43 F7 18 D7 67 F0 5C C3 B5 F4 3F
 F6 0A 96 9A 82 2D 11 4E CF 42 6D 98 15 4D 69 47
 4D CA AF 99 9A 30 BE C5 C2 A4 A6 84 9A 5A E1 74
 D7 91 0D 63 40 17 6B 3D 90 E8 34 12 46 35 D6 25
 10 E6 F8 F2 AE 76 C8 62 5C 3F 1B 46 88 9E D2 0F
 92 2D 53 4C 35 D2 78 C4 01 BB 4E F3 FA 23 1E 46
 B7 E5 A2 AB 79 7D 75 6E 8D BC 50 33 8B 84 85 1B
 FB 90 73 D5 C6 EE 99 CB BD 14 7C C6 17 D8 BD F1
 29 5A 3F FA 1A 2B 57 DF EC 35 06 78 BE 96 45 7A
 E6 09 B2 82 14 E4 AA FC 83 BE 28 89 CB 62 0E 55
 9A 3C A4 F8 02 12 4B AB 4D 3C 11 37 BD B9 5A 17
 CD 48 30 EF D1 9C 03 EE 93 6E 57 C8 6D 1D C1 5D
 6A 1D 44 8E 4F C7 FB 3D B3 8C 71 A3 68 90 78 9E
 A6 92 2A 31 51 B9 05 D2 B2 74 3E B1 DE 62 10 13
 C2 4B EB F3 B5 B6 47 9C 3D CB 0D 14 96 22 6A A6
 6B 27 4C BD 1D 44 99 5E E2 6A 43 79 61 AC 67 B0
 8C A4 70 5C E7 D7 67 1F D6 E6 B9 A7 F7 14 EC A7
 C9 D9 44 72 EF 82 45 65 C3 FB D9 F4 40 DF A0 32
 36 1F 6A C6 66 7B E9 3E 6C 4F 19 55 BE B6 0B 73
 C8 7A 87 C6 9C 0B BF 49 C9 05 CA 0B 32 BF 27 04
 21 F2 31 9E 55 67 93 A2 6E 01 B5 AD F0 B9 DD A6
 CC 07 A7 4C 7A 4C 61 35 3B D9 57 CF 16 27 26 5E
 37 11 A5 DA 3C B1 9C 3C 07 49 92 F4 B6 E8 15 3A
 49 95 A4 3F C5 51 BB 3F 43 FD 32 6A A9 15 EC 43
 26 CD 73 46 42 EE 56 08 7B 72 0F 6F DC 7F 6A 92
 18 E5 3C CA D0 A0 02 70 93 F8 AF CA 58 17 10 1D
 2C 42 CE 1F F1 F8 43 36 83 AE C8 6F A6 90 9E 9C
 C4 7B 8B 70 C0 99 89 88 D4 DC 62 DC EC 56 06 CE
 26 FA F8 41 5B 95 79 C9 92 10 70 B0 E8 C1 17 AA
 19 DE CC D3 E9 6E 48 D5 17 BB D8 4D D8 73 FC 6F
 9E 4D 63 96 B8 93 E9 26 5F FC 1D C3 27 F0 20 9D
 28 23 A3 0C B9 6B F7 EA 66 E9 18 3F C7 A6 62 C1
 69 9B CC A9 39 88 B3 73 22 E7 98 C9 2F 87 4D 34
 54 A1 20 12 49 3C 72 C4 91 EF 51 9E 13 66 3A FD
 62 33 B8 C7 93 B6 AF 7B B9 72 B0 BB 71 91 B4 7F
 7C 4B 82 72 4D 8A 37 70 A1 63 31 8C 0F A5 81 F5
 42 A5 AC AA 4F 47 92 8F D7 CD 0E 0E 07 BA 9D 82
 B2 74 6C F6 B8 A1 7F 0C 68 DA 6A A6 14 AF 04 69
 EB 81 F5 96 1D E1 DD AC 45 E9 5E 35 E5 12 BA C3
 EF 53 F1 A0 95 AA 88 67 E2 77 E6 21 30 F4 0E 6A
 67 F8 CA 0D CE F3 AD C1 E9 E6 48 A6 07 69 43 42
 B7 83 F1 6F 70 7F 5F 17 C6 CC 8D 87 E4 C0 83 22
 23 11 88 53 E8 E2 79 F6 FA A4 79 BE 48 B1 B1 38
 5D 00 96 E9 AE 5B 08 61 2E 46 46 E0 61 F7 E9 15
 17 6F DF 2C E0 FD A5 FE 3C 79 E5 F7 A0 72 41 01
 DB 5F C4 06 D3 23 86 9B E5 CE CE 5A 3B 9D DF 9F
 D3 5B CC 0C FF B8 EF 8F C9 98 7A 61 2B C8 01 39
 D7 19 39 B9 3D A2 FA DA DF DD 48 E4 83 F3 D3 40
 EB 16 D8 E3 9F BA FC 48 4B 01 C1 54 66 5D EF 33
 0F 01 EF B8 F9 E4 86 67 74 2C B0 AA A8 A6 A3 2E
 FA 0C E7 BC FC 11 6C DC 2B F2 ED 41 8F 22 11 95
 60 E7 35 9E 69 4B AB 79 7F B4 F3 C8 A7 54 D0 45
 9A 74 33 D8 CA C6 B7 9E AD 7B 40 3C 12 FC 26 C2
 18 BA 81 24 73 32 6E A4 A3 71 FE C4 9B 02 30 4F
 EE 5A 4B 3B C1 67 15 B6 69 63 A3 6B 9B FD 61 E9
 A5 70 38 5B D3 97 AB D8 B8 72 D8 51 6E 3F FD 2E
 5B 86 6D BF 5B EB 71 4E 21 FA 79 81 25 C4 10 1E
 1E 37 40 F1 E6 D8 EF 32 B8 F9 02 8A 4A D5 23 BB
 F1 5E 7F 4C F5 1A 60 08 C3 93 BF 4D 38 42 30 96
 01 DA 3E 26 41 D0 8E CC 1E 0B 0D 86 8B C1 8F 34
 18 7C E4 6C 3C BF 39 65 03 BC 9B 2A C4 C5 C5 77
 B4 C4 1F D5 80 33 82 B0 37 2E 5C 1D AF 61 0B 13
 C2 D3 87 8B 46 B7 DC 36 B4 4E E3 41 13 10 06 A0
 35 F6 7C F1 F0 82 8C 50 06 59 3A 0A 74 5C 25 54
 8B 8B 60 43 CD A6 75 AB DC 9D 40 F2 91 A5 52 AF
 05 F0 D7 9F 1B 55 26 E9 EE 7F 30 6E 54 B8 78 DB
 F1 C2 3E EE 7A AE 8B 29 C2 1E 37 28 93 CE F5 4F
 BD 80 49 D4 26 3C 10 66 AC 27 CF 46 D5 03 A0 E1
 43 6A 9F B3 D5 12 5B A2 34 1A 78 40 02 2C C4 0F
 1A C0 E1 D4 14 9D 76 2A 4D 41 1B CD 35 94 E9 86
 1C C3 CD 9C 84 05 15 B0 1A 2A 06 87 D5 5C 17 0F
 62 5D 5B 57 21 BC 4B 4B 64 5D 7C 11 37 E4 78 FD
 ED 05 7D 8A 31 DF 8F 69 24 D0 CD 1C 43 3E A9 3D
 3D 8E 35 58 3E E5 7C 86 24 EF D3 20 0C E9 7F AD
 E9 77 E6 D9 ED 93 7E D8 10 E0 D3 60 7F 05 90 E9
 CF 69 8C E8 E5 AB D8 E6 CA 9C 60 0C 39 AD F4 0E
 C5 40 FF AE E8 F2 03 98 3C 32 73 30 C5 FE 92 76
 AB B5 C8 FD 92 04 24 76 FA B7 09 78 5F B5 4B C6
 BA 33 C1 AB BA EF 74 21 4C E9 40 5B 06 CE 55 82
 86 3D 93 64 1A 51 AA C8 72 CD 5C D3 75 41 3A 33
 FB EC 04 46 C1 C6 6F 29 6D BD DC 78 46 FD 60 FD
 7F 0D 9F 3F 61 B9 7F 27 1A CB 6F EC 19 29 D4 82
 2D 72 30 EB B6 24 51 F7 EC 08 04 0A B7 5D 56 E2
 55 60 BA 10 8F 06 C7 7A 62 1B 23 05 A3 C4 C1 59
 EB 07 F0 A7 2C 04 38 00 E7 73 AC 69 64 AF D6 49
 F3 F0 64 FD AD F6 EC A9 33 DE 1F 33 95 90 07 16
 FE 20 14 B3 68 1E 0E 0C A0 70 6B BB AD 10 A4 41
 9E C3 B9 A1 AF E9 55 2B 17 40 49 26 45 61 5D 86
 2E 08 BF C8 5E 65 61 18 A7 46 E0 53 6C 7D 4D 94
 A9 F3 C8 5A 21 27 F6 CD 0B AA 69 94 1F 69 74 8E
 15 3B 17 16 67 F5 FE CC 6D 09 D5 A6 47 55 20 27
 41 38 31 21 75 AA E7 19 68 F7 60 CE 48 38 F5 9B
 EE 16 BE 02 BC 74 64 21 5A 53 75 9F 21 88 5A 4A
 00 45 E4 64 5E B3 A2 73 B9 B0 DC 14 31 07 B6 B5
 ED 50 17 66 B2 94 E0 53 47 31 85 DE FD A0 7E 28
 FD BC 5E 37 45 A2 68 6F E9 82 33 92 A7 B6 3B DD
 93 39 73 39 87 78 F0 22 AC F9 A4 CA 2E E8 38 08
 68 DC 7C 97 E8 A2 83 E7 25 2E CB 60 82 82 3E 60
 28 28 6F 46 F1 21 2C E7 B5 43 A5 31 D1 DC AC BB
 C3 9D B3 74 93 EC 5B F4 1B 47 77 13 FC 2B 35 CF
 C8 BF CE E2 46 7A CF B9 5C F7 5A A7 55 15 6B 19
 42 8B BF 63 73 F3 36 17 7B D6 C4 A9 3D 97 EA 2D
 31 A1 9F B8 A8 A0 D9 19 53 D3 F4 42 56 91 15 95
 6C EF 14 1C 0B DD E3 97 DC 1F 32 35 43 2C 96 DE
 17 5E 27 16 61 BF B6 47 29 48 FC 4D 42 04 A1 48
 8E 7A AB A7 57 8A B3 8A DB C9 4F 8B 1E 61 0B 95
 01 F8 0D AD E4 F7 BA 94 1B F9 51 E3 C8 48 55 16
 43 26 EC 77 3A 1C 08 E0 24 94 25 39 37 E8 B4 45
 98 8C B4 4D 63 00 B9 A1 58 FA 84 6D F0 2A 02 D6
 E4 6A 6A 73 E0 F8 2A E0 E2 47 6B B3 B8 CE ED 77
 B7 1B 12 BA BB 70 4F E4 84 A8 6B 15 47 F2 7B 2A
 B0 51 AB 45 DC 11 BE B0 8D 3B A1 46 DB 27 50 CB
 C7 D1 3F 76 D0 C7 FD D3 C6 79 16 5F 21 8F 45 C5
 19 F9 3B 7B 97 6F 11 4B 0A C6 13 75 21 55 A1 37
 14 A6 BE A8 F6 9D 5E 70 40 78 58 0C 19 68 61 A9
 3C C8 80 20 02 1B BB 4F 58 E9 78 A4 8D 2D 09 3F
 D7 2E 69 BD 09 04 7A 1C 6F 2A 89 99 08 B2 2E 12
 F3 46 DD 27 D5 9E B0 A7 B3 32 FF F2 DF 4A C3 74
 BB 72 BE F1 97 97 B5 D8 B9 9C 0C EB 91 9A 37 A1
 A3 6E 64 BE 75 F9 08 41 0C 41 D3 A8 8D 4F 3E 22
 A8 AD E9 08 B1 02 09 ED AF 3B A1 7E 4E 40 50 F3
 F6 26 66 0E 5D 1E D1 A7 7E F6 72 83 4C 57 11 BB
 ED CD C6 32 2A 10 92 BB 05 3B 54 21 E0 9E D8 FB
 E0 1C A9 16 A2 7D BA 70 6F DB BD 16 6C 7F EC FB
 C5 B9 E4 6D A1 26 9F F2 D4 B0 4A 1C 4F D4 F6 44
 36 54 AD 5F 0C 26 45 2F AA 5E 34 AC 30 48 84 00
 5B 24 6C 7E 47 45 FB 25 3E 09 51 D2 B9 30 99 9A
 7D 28 2A D1 34 0B 7C 1D A9 1E 4F 82 7F 83 FE E7
 0D 73 B6 00 E6 61 5B 42 39 4A DD 5A 74 85 52 62
 53 0D 79 16 C0 67 12 62 68 C2 84 CA 86 CA 03 BE
 FD F5 A1 00 54 0E F5 6B 3B AE C5 5F 22 77 BD 23
 44 6B 5D AC CF E2 01 EB 51 D0 19 BA 86 AB A9 67
 A5 63 95 16 2A 38 A1 D8 75 0F 7E 1D 6F 59 D9 8E
 4D F6 2E FF 7A 02 29 D2 F4 61 99 BC 10 42 9D FD
 9C CF 93 F0 0B F4 1F 58 DA E3 CC E5 FD 80 A5 26
 17 D3 6B 79 1B 68 C1 CE 84 CC D3 5E 6F 2A 77 30
 1C FB D8 B1 F5 0A 35 19 FB 38 A8 14 56 BD BD E4
 4E A4 24 7E 73 09 FA 9F 76 A3 F5 5E CD 9D 2C EF
 17 D0 CF 3D D7 F7 37 E3 AA 34 0F 90 2C 5E D0 97
 0E 67 85 4C 77 BA FD D6 E8 CF 6B 14 36 53 21 0A
 8C 0A 62 2C AB EE 24 56 44 60 38 85 EB 88 05 B5
 A6 70 6C 08 2B AD 20 14 B4 49 16 1E B1 E3 85 49
 AE 87 32 E4 07 F9 FF 19 BB 64 20 92 4F 69 4F 71
 88 B1 9F 8D 18 8A DB 4E B4 D6 E2 C4 1E A3 85 45
 71 40 F8 5C 7A FB 95 2F 32 B0 9A 2A 64 10 49 03
 E3 A2 A8 06 0F E0 F3 6B CD 76 52 3F A2 FE 3C 1D
 D0 33 80 AC 75 CF BC A5 E9 56 69 73 84 FB 38 DF
 6B C3 27 B1 4E 1F 00 21 E3 BC 32 EA 35 96 45 A7
 BA 32 F8 B5 11 B1 79 5C BB 78 61 7B C3 10 14 6E
 49 EB 42 D1 A5 5B D1 D7 84 38 48 44 6A B8 3C 72
 86 BC C8 D4 6A 59 E5 A9 FA 8F 6D 90 A1 B0 D4 6B
 4F 9A D7 93 7C 74 90 3D B8 F5 44 5C 6A 56 FE BC
 02 F8 FA C3 F1 C3 46 83 59 46 4F 61 0F 93 00 67
 19 C4 5E 0F A2 8B C8 D0 85 CA 21 27 39 54 1E 52
 5B 6B 86 1F 82 F0 5E DB FA 98 C2 4C 78 BB A0 BA
 EC 29 5E E7 05 4E 75 CD 18 E0 37 66 01 4C F4 7B
 60 92 77 01 A4 A0 46 28 95 40 92 87 02 3E AB 27
 BD 2B E3 C6 DD D1 58 F1 B3 CB 68 87 7F B2 21 23
 DC FC 8B C1 16 39 13 FF A3 40 14 52 A8 B9 C9 05
 08 60 B4 ED 4E 66 B1 56 D7 31 D2 11 3F 0F 90 46
 4F 08 97 FA B5 08 9E 97 13 85 E0 38 6E 81 38 60
 80 9E BE 08 06 F6 1F 30 BF 99 34 95 8D 4C AA F9
 1D F1 2A DE 2F E1 CC 09 47 70 3D 30 B6 FD 46 3B
 F6 3B 53 65 2A 8E 80 BE 6C AB 41 1C 27 F0 73 D0
 32 EF 35 DF B7 86 10 D2 FA 78 3D F5 BE BC 8E 4B
 B6 7B 26 43 0D 0D CD 0F 03 48 E3 59 B0 F7 49 19
 A8 EA AF C0 66 9C 45 E2 1B 54 86 6D 41 45 8C D7
 83 04 20 06 98 60 41 D6 DD 4D 49 E6 6B 20 3C E4
 46 5B F0 E4 2B 88 39 E8 7B 2F 21 E9 1A 78 D1 47
 70 38 DB 46 0F 39 3B 37 7E 17 C8 D7 D0 D6 7B 70
 45 C8 C1 61 6B EB 44 D3 71 79 ED E9 C4 1D 11 EC
 CC 24 04 4E 27 67 56 66 2D 75 8C 64 65 59 7F FA
 D0 B5 11 CF 65 3A 79 FB 7C F6 B3 85 6D C7 D5 A6
 10 60 A4 52 3B 64 B6 72 95 2D 78 5F F4 54 76 72
 53 36 CB B4 E9 07 D4 6C F7 9A 12 0C FE B7 C1 8D
 E1 CA 51 65 C2 0B 95 83 E2 42 10 69 0C AC 58 B6
 EC 1D FC FE 3C F7 D5 FC 51 43 D9 03 18 AF 91 BF
 5D 02 CA 74 3A E9 68 91 CB 94 DC E3 F5 C6 18 3E
 E5 D0 51 2C 93 11 48 52 E5 7B 24 41 22 F0 47 35
 8F 6E 9F CB 35 35 B2 88 AE 13 E9 CA 3A 20 E7 71
 B1 CF 09 2D 08 CD 58 97 53 0D 5A 5A DB 61 55 F6
 DC 0D 88 5A 35 E6 13 6D 3E 37 DD C7 0B BA 2E 96
 C8 58 DA 8D 61 60 03 57 D5 A4 67 45 94 99 01 63
 96 28 31 86 2A CE 07 28 C9 10 D9 DF 14 20 0C 06
 68 4D C3 B4 F6 46 A6 D7 7F D4 40 E0 94 75 73 13
 4D 16 5E 93 EC 5E F2 15 DD 94 91 7F 48 17 DE B3
 ED BC F8 59 27 40 25 72 89 47 3E 13 5A 21 A1 15
 4F 40 A4 00 CE 9F C3 CE 9A BD 8A F4 EE 3B ED 90
 FB B3 1B D6 8D F1 4C FF E4 D4 E6 21 8D 18 6F BC
 CE 6A EE F6 22 A5 0E D4 9D B6 10 53 B4 F2 CB 37
 38 79 C5 58 15 A5 D3 7D AF 71 10 5E C2 AF 54 03
 85 2F 52 4A C2 E4 13 FA AE D0 03 C0 40 3C B5 42
 A6 E4 89 AC 28 92 21 F0 11 EA BE 2B 95 E5 16 F7
 6D 66 26 59 13 70 58 1B 96 2C B3 4E 93 B0 C1 17
 A6 AA 84 CA 0F 5C 0F 02 BF D2 14 53 33 63 C7 55
 21 8E AF 2F CF D1 91 68 8C 7D 6E 8C 9B 8C 85 D3
 DF 81 90 3E 84 71 69 2A 72 72 B0 A7 D6 E2 36 DC
 B5 83 73 FA 2D CA 71 E3 10 CA 3B E7 DE A8 88 ED
 64 BF 3F 94 0B 55 76 FB 0D DB 72 5E 9D 8E 7F 81
 59 D4 6B 0F D5 AD 90 62 43 84 3C E9 A9 B0 6A E9
 D8 DA D4 B9 F6 46 CE 6B 4A E9 2C DB 9C 73 99 9B
 9B D2 8D 4E 36 0B 37 67 AA 3E 48 EE EF E1 4E B7
 0D 5E 64 DE BA 5E 76 B2 0D 22 50 05 C2 97 BE 20
 4A 21 96 C7 65 2F 2B 5A 09 F2 E1 9A 62 56 4A 40
 92 51 7E 3B 30 1D 64 A0 B4 78 E4 05 01 4C 39 1A
 34 1D ED 6B 32 47 A2 BF 82 74 C4 3F 96 61 67 1F
 4B 28 AA CC 59 BE AF E2 9E 1B 50 2F BA A0 09 A6
 96 2A 86 1D 41 ED B6 E0 9F 22 E5 61 F6 F7 58 7D
 A9 44 57 64 60 9A 45 C6 89 8D 5B D4 3E 81 7B 03
 9F F7 77 8B 37 DF 26 22 80 2A 3B 7C 89 12 ED D4
 76 BC 79 C5 0F A1 E4 70 0F 6C 42 35 64 B0 73 57
 64 E4 82 2F ED 8C 5C EB D6 B4 B0 10 E7 6B CC 44
 BB 19 54 03 EF 58 57 81 FD 63 16 DE 37 AF 61 89
 EB EB 60 94 C8 C6 DE 66 28 B4 8C FA BE E9 8C 2D
 8D 32 C6 28 BA F8 48 DA 8D BF B1 E0 2A 95 B9 15
 CE 37 6E A6 5A A3 BA 57 C8 2F A9 87 6D 54 07 A3
 BA 2C 00 83 9A 50 F4 07 6D 8D AD BD 25 AB 23 41
 51 F9 70 12 8A D2 39 52 CA 59 18 C4 E9 B5 DB CC
 C3 9F 77 E9 17 45 F6 24 3B 93 8D 57 68 C6 FB A7
 46 16 13 A5 F9 53 EA AB C9 17 B8 71 F4 BE 8C 3F
 CB 35 FE 13 4D 86 98 15 BF CF 92 2D 5E D6 E3 F5
 40 EB 95 26 E0 BE 86 57 7A 53 D8 3B 45 70 F6 01
 3F 7B A1 19 78 2F 46 D5 E7 84 1D E1 D3 09 82 1B
 DC 6B 5A D9 DA D0 37 32 5B 0F CF 5E 4C AC 5B 9E
 A6 24 D2 71 AD DB B0 0B 3B 26 4B 5A BE 1F 3A 6C
 55 A6 D1 80 68 6F 2A E4 E6 DC 9B 9E 12 1C 4F 20
 1F C9 B4 36 AF 43 99 CA 8E 1C C0 65 DD 4B 56 77
 84 43 1D 4F B3 29 30 62 A4 C4 5E AB 40 1B 2A 0C
 A1 64 2A 7B 6A 79 5B BC F4 E3 2B 0E DD 55 54 4E
 E3 F0 B8 CA 75 DA 4C C3 60 0A 67 86 D5 57 E5 4C
 A1 01 12 44 34 F4 BD 60 C3 77 CC 1A 8E FB 38 7C
 66 F2 7B 36 BE 18 B7 56 EC 0F DB 14 66 40 9D D7
 C7 D6 2E 89 C7 C7 40 EE DB 81 39 48 22 E6 A4 1D
 46 D3 00 07 01 F2 AA 0D 0F D8 93 D1 DB F2 11 7D
 9B E7 E1 D3 69 C0 32 EF 63 EC 35 25 24 31 92 8F
 EE CD AA 4B E9 81 F7 86 61 C8 39 FD 41 4D E9 A3
 89 11 13 77 A3 E4 B0 DA 9E DC A8 C2 5C 90 B9 BE
 24 47 45 81 CA 43 9A A4 BE 81 46 D9 DB DC 9C F3
 E0 7C A1 E9 6E 23 27 16 CB DC 0C DB B3 9A E4 C0
 13 47 07 88 F0 78 59 92 48 6B D4 54 8A 55 FF 63
 5C 55 33 72 33 E7 A5 F2 CD 92 43 B0 42 A7 74 25
 A7 87 5D 04 9E 24 04 67 56 E2 FD 0E A4 2C FF DC
 45 9A 37 F3 C1 C3 59 5B F0 2D 74 54 E8 E7 CF 57
 E3 6D 58 B8 37 8E 45 C5 FE 61 BC DF E1 8C 9F 7C
 A7 B5 03 CC B3 7B 87 F8 3A 7B 63 9F 8F A6 B2 D9
 69 9E 64 0F BB F9 BA AD F3 4E EE 89 4C 27 81 11
 94 0F 4C 99 67 A4 02 89 9C BC 0C 1E B1 34 02 DC
 22 AA 02 BD EE 79 D6 6D 19 E2 18 E9 48 C5 0A 3D
 F2 63 3A 3A 68 2A 86 A2 DD 52 4B 27 BA 5C BE 6B
 0A B0 3F 79 9C 39 E9 BD 71 57 A7 7B 12 BF 7C 5A
 42 A2 D2 2B 9E 71 D6 E8 03 01 CF F3 8A B7 7D B0
 2F 40 55 6B C6 72 6F C2 18 BA 27 A8 0F 30 43 37
 7C 6D 30 31 DD 13 6F 26 FE 6B 76 35 57 F7 FC 56
 5E DE A0 5B 81 A2 81 4C 96 BD ED 98 F4 96 D9 65
 55 4B 7F AC 63 87 74 2B D0 DA A7 AD 3D 0E 2E 3C
 BA B1 3A 74 23 EB 9E 50 8B 3F B3 09 1B 27 A1 5C
 6C 1E 4D EB 54 90 CE 2C 8E E9 77 26 0D DD 96 A2
 97 D6 26 E8 00 FD F2 26 AB EA AE 4E 74 6D 61 B6
 D8 E1 5D A1 6F 41 6B 59 E0 0F 26 43 A3 BA FC 93
 96 09 85 C9 82 08 73 6C 2F F7 45 61 0D D8 EB D0
 7E C7 96 5D 66 6C C9 1C 81 63 78 E1 24 DD 13 40
 3F B6 52 2D 72 1A 09 96 40 B5 C7 BF FE 79 AC C4
 A8 7D 8B 20 F7 16 5E B0 59 F4 1E D5 36 A6 7C CB
 68 24 43 9B 67 20 97 0D C3 66 01 E5 7C DD FB 06
 BC BD 76 41 BF BC FA CB FE AE 23 2A A1 BA 5F 12
 05 EC 84 FD D5 D0 FD B6 9C 66 19 5B 95 7F 97 DC
 AB 51 E1 F1 C5 FD 50 0F 05 C7 CF 16 8F F5 DA C9
 E3 81 CF C3 1F 70 2C 4D C9 4E AE DB 01 5C 92 D1
 65 71 BB F6 FA EA 3D 8C D1 6C 35 5A BC 2E 8E E3
 AD 29 05 57 9B 8C 10 E7 FF E7 DC DA 77 77 87 E1
 6B DB 8E CD 72 C8 84 25 5E BA FE D9 99 14 85 1F
 28 A5 3C 92 54 09 AF CC 0C 14 38 57 5C D8 6C E6
 F0 E5 70 4D A9 68 95 4B EA B2 21 16 53 CC 0D 17
 D2 67 5F 33 0C 5A 4E 14 B6 39 5E BD 87 0E F3 0C
 C1 85 98 84 66 2B 6D AD FB 83 35 9E 33 78 22 A8
 3C F5 BD 3D 05 7F 3C 67 97 BC 99 3D 67 32 45 60
 CA 30 73 38 7E 35 20 1D ED 07 77 CD D6 EF C2 EA
 9E ED 06 27 A6 61 48 68 7C 8B A7 57 DD 12 C9 4D
 D7 03 F1 54 0A DC D9 25 B1 CD 9A 27 F0 EC 4D D0
 EB AD 66 F8 C4 D2 B2 5C E4 61 FB D1 BD 0F 41 41
 F7 70 22 78 B1 BE 19 B3 6F 63 B6 AD 4D F9 63 98
 7D DE DE 91 D6 57 27 7E 21 CB 36 87 43 A6 8C 27
 50 40 70 07 3D 4A E6 3F 06 D3 49 94 D2 B6 A4 3D
 89 1C F4 9F E4 3F D5 1A 9E EB CC BB AC CB 12 03
 CF 79 5B 0D 2D A3 29 5B 31 87 BC 0B 73 57 88 B2
 46 82 01 6E 3F 90 3A 4B 87 3D E6 12 C9 4F 48 0D
 66 E6 DD FF 33 BA 74 FE C5 0A E3 C6 E6 BF C6 8C
 84 C0 AC C1 56 EF 18 68 66 87 EB 1A 2E 7A 66 94
 6A 71 0C FA F0 F8 90 AE CB 42 85 F4 88 D1 8C D4
 4C 6A 02 8B 63 AA C5 FB 41 87 ED 38 6D 7F C3 DE
 AB 66 82 8F 77 CA 33 45 55 C6 46 DD 44 FC 11 C4
 06 37 1F E1 D6 58 FE EB 44 A6 A1 8E 50 09 9E C3
 BF DD E1 8B B2 72 7A B4 C8 83 6F FA 52 68 60 F7
 9D 89 F5 A6 1C BD D6 41 7A 34 1E 8F 61 10 49 F3
 36 35 C7 F4 9F 84 A2 41 5C DD D1 45 F5 A6 7F 4A
 82 46 15 3D E0 0D E5 F2 36 2E 43 F2 50 76 D0 28
 08 34 9F 40 2A CF E7 60 76 28 66 75 10 F7 D0 41
 E6 5F 65 50 59 C4 08 0B 9B 97 96 E1 8A 81 97 A8
 69 9B C7 B7 58 2E A2 AD B2 C3 51 04 70 DF 39 C7
 5E F1 1C 95 79 8D 6B 9F 36 EE 23 73 7E 9E AB 29
 6C 49 D5 6D EE 75 D3 C2 E3 DB FB DC 0F 95 0C E9
 E8 C2 D7 0C E3 BA 39 31 B7 C6 C8 F5 39 D1 81 74
 3F CC 89 6D BB CC F1 59 31 7E CF 0D 77 06 9C BA
 AC B0 BF DD 88 61 18 F7 09 56 D3 8B 79 DC 6D 9E
 C8 A7 77 93 9A C2 0B 10 E7 B2 BB 62 1E F7 0B 60
 3F 8B 3F 4B E4 AC 33 6D 56 2E 9A 6A 6F A7 B7 E6
 8C 88 A4 5B E4 B0 F2 AC D2 E6 D7 4B DE 0E F4 7B
 5C 12 0B 9B 6F 3A C6 2F 28 B0 49 AF 55 03 50 4A
 DF BA 68 5A B0 94 DB 5B 9E 7D C7 FD F6 1F E5 E2
 13 9A 6E DC 0D 92 6D 7F 6A D2 14 77 EE EC C2 70
 F6 27 BB EE 09 7D 30 E4 26 60 EB 4B F5 DE 39 20
 0E 54 AD 95 1C 97 93 AC 05 F1 22 A3 8E A3 FA CC
 BA F0 EB 2A CC 82 68 C0 85 12 24 54 6A 38 BE 9C
 12 1B 1D 06 8B 6C E9 E1 E3 04 52 78 50 D7 8A AB
 CC 82 23 1D A9 54 80 65 86 85 73 FB D9 31 35 F9
 3F 33 34 C2 0C E6 63 A1 ED B2 2A 4C E4 8F AE AD
 E0 9B 48 27 B2 89 F3 B5 EB 8F 9C 2A 41 35 F6 5E
 A9 42 65 3A 2A 90 BF 50 78 F5 A1 63 57 96 02 8E
 3F BA 28 71 CA 89 CA 5F C0 8A 4B 02 7A F4 E4 75
 E6 16 30 C1 55 89 B5 2F C4 09 22 39 72 DD F7 91
 CB 5E 47 FB CF 15 C9 4B 37 F6 9A 1C BB F5 49 83
 F1 62 33 62 C2 EE 01 23 78 AA 03 81 0A C1 76 D2
 63 9C 20 46 9E AF BC 35 27 1A FF 3C 9C AA 1E 70
 BB C0 82 A2 3C A3 12 BA 9B BD EE E4 25 C9 3A 96
 F2 66 E3 B7 50 B3 31 72 86 61 A6 CD 27 7C 3C 1D
 D1 8D 90 21 98 96 27 D4 E9 22 48 46 6A BC 57 4A
 1D 90 99 B2 64 86 AA 87 2A E3 D5 27 B9 6B EE CC
 65 D4 F7 19 76 9A 0C EC D2 87 5A BD 39 93 18 7B
 55 D0 14 A4 BC C5 9A 9F 56 F5 D9 CB 3B 28 12 AF
 8D 1B 0F D0 B1 06 94 3B CE BC 00 37 62 2A F1 20
 68 97 F9 B0 DD 76 2D D3 B8 4D 2C 2B 06 66 EA C6
 A2 57 FD 47 4B 93 42 05 77 38 A8 66 F1 F6 FB EA
 A1 C9 B1 CE 25 C6 6A 4D F1 34 79 A2 33 BC A5 39
 EE 84 7E 06 5D 98 93 9D D1 31 D8 65 0B 8B 77 53
 AF 6F 18 12 51 05 A0 46 BE 0B 48 99 97 60 63 DB
 01 A4 EF 45 60 C4 35 98 71 3B 09 30 AA 26 FB 99
 34 E6 DB C1 3F CE B9 AD 70 84 4D C1 C5 9F D8 21
 78 0B E6 65 46 0D C8 AD AC DA BF 2D 5E E4 85 6B
 29 8C 54 07 65 79 A8 FA 2F 0A FF D2 5C 28 85 E1
 F9 FB E8 8D 9E D9 38 16 96 84 D8 13 21 D1 FE 5F
 D7 DC 21 D3 98 BD 92 70 27 52 A5 7F C0 1A 5B 94
 AA 14 13 F3 E1 86 75 8F C1 1C 14 52 C6 21 2F 3F
 8B 26 96 AA 17 5D F8 3C 51 11 4B 97 20 44 5E D1
 99 2C 46 23 C7 9B 64 5B 1A F7 37 7E D6 FC AF EF
 F3 54 F9 2E 81 7A 5C C1 34 FF F5 AB 08 E0 54 4C
 D1 D1 46 A4 B9 CF 66 34 D5 73 0D 41 73 A8 F8 3F
 40 59 A9 7D 51 9D 84 41 07 26 52 15 D1 44 DB AC
 89 15 56 8D 9E 0F 4A 60 6A 64 16 15 A3 F8 7E 2A
 00 1E 00 5A BD 31 0B 1A 46 A8 5C 8C F2 4D B8 84
 3C 3E 60 AA B9 56 31 0D 5F 2D 33 81 90 D7 D6 35
 4B 21 6A E9 ED 47 CA 42 B2 19 B5 14 FE F5 95 0B
 25 46 1D CE DA 31 2F FC 79 7D 4C 55 D3 01 3B FA
 8E C2 30 65 6A 07 8A C5 A0 0D 24 19 B0 F5 B5 DE
 0E A7 C2 26 59 01 A4 CA 71 20 AA A5 A3 E4 7E 0E
 1C B7 F7 41 8A 66 11 F7 3C A4 BD 5F 34 1F A7 C4
 EC 13 AD DE 9D 99 7C 2F 86 B3 78 F5 91 DA E1 D5
 09 46 46 CB E2 BB 23 F0 88 FA E7 1C 7C 29 35 D4
 EF C3 B5 40 10 F9 5E BD 46 B5 F8 53 79 0E 83 1B
 B6 F9 A4 2F 42 8A 67 29 80 7F AA 9F BA 14 C9 4A
 B3 C1 80 35 86 D2 D8 C5 82 15 63 0A 09 5F 88 A4
 C8 BD 90 FC D3 62 B8 99 06 FB A3 99 40 DE 90 8F
 8A BC 61 E7 6F 3C BE D1 33 FE C8 DB 66 FC 1B D8
 B2 EC 5D F2 08 3A FB FD D0 76 A2 18 FE F1 3F A6
 06 82 4B A8 0E AF FE 46 E0 83 67 71 F9 49 F6 92
 14 A4 F8 20 97 C7 E8 70 9A A5 AC 65 D0 F8 00 99
 BA 4C FD 86 28 32 86 12 9C A8 23 32 F0 BB CE 2E
 52 62 1D A2 0E 2D 48 97 22 A1 59 83 D7 DB 9F B4
 3B EA 1A 2A 71 71 70 7B C1 C3 A5 5C 7A 89 F6 43
 45 69 80 DC 3C 6F DB E1 3C 0E DA 92 A0 23 8A 82
 92 85 54 45 E1 45 38 1A 10 94 C1 84 66 AC 20 DB
 C0 91 B2 65 45 82 0D E8 D3 39 21 65 AC 6F F2 55
 BF A0 6D F2 FC BE 1F 17 D8 89 6A 4E CC 6A E7 61
 BA A5 53 97 2B 43 31 D1 EB 2E 9F D2 6B C8 00 8D
 2C 25 1F 6E E0 2D 76 F7 31 07 83 81 CC DE 06 FA
 F9 6B B6 E8 84 B3 D5 6C E9 D4 4B EB BE 95 84 8B
 BC E1 FA D1 22 AD 34 61 28 6E 09 41 1D 3C 42 E4
 4B 6D 1E 80 43 E9 00 BF D2 98 FF 95 0B 56 79 B3
 38 72 9D 11 DC 00 4B 99 0F 34 66 F2 40 28 0C 36
 70 C5 9F 80 BC 2D 01 9D 58 A0 79 E2 6F 4B 34 5B
 6E 58 EB 90 CE 45 77 48 EB 1D DA 0E 0A 61 BA 99
 38 F8 C1 CB B1 02 C0 5E 4A 62 20 08 1C 03 42 87
 F8 09 0B 8B 1D A5 0B FE 04 9C 42 6B 38 69 62 7D
 8E A1 07 33 15 11 B2 F9 00 89 BE AC 95 2E 4D 0D
 4A 8C F5 C6 8E 42 FB CE FB 38 D1 F6 34 05 9D 2F
 9A 57 77 7E F0 F0 BF 73 02 0D EE 8B 66 4C 3D B4
 AE D5 EC AF 36 42 23 FE 63 75 9B F3 62 FB 5B 0D
 6B 54 B1 E9 8D CD 4D 5D 4D 2D 75 7E 47 49 91 BD
 B2 EC 0D AE 18 1B 16 5B 7C FE CF 9D FE 81 BF 51
 C8 76 1D 9D 07 D6 EE 07 4A 61 44 D7 FA 67 08 BC
 8A 2B D7 A4 58 55 28 F7 B8 B5 CB CC 66 CA A5 B0
 8A E1 B4 EE B6 AB B2 E8 BA D4 31 05 B4 EB D7 F6
 48 EF 6E 9D 0B CA 59 3E 69 28 7F A1 E7 B0 B9 47
 C2 D4 35 3D 07 E8 A0 0D 45 6D 41 35 84 B3 E1 A5
 89 19 2F A6 26 EA D1 C4 3E 0F E8 63 11 4A D4 9C
 E8 25 05 B3 ED 2D E1 4B 21 B9 24 30 CD BB 0F 13
 F3 B9 93 AE 38 82 70 5C D8 9E 92 A9 92 2E 6A 5E
 3E 90 79 2E 62 F5 D5 36 2F EB A4 56 83 A3 90 4C
 2D 6D F3 8E CB 52 CD BA B2 D3 B4 45 01 8E 51 CA
 1C 9A A2 E6 65 FB 6F 06 5B EB B8 D3 DA 73 E3 D3
 1E 37 0C 38 1D 99 4E 22 3A 80 A6 78 94 DF 8F 9A
 D6 0B B9 3E 02 6C F9 3D 22 79 96 80 98 1A 43 7E
 34 C9 C7 3E DE 73 E7 C2 15 98 F1 DD B3 C8 DD 3B
 AE C2 55 C4 D4 DF DC 4D 88 62 3F FE 9C 82 0F 0F
 31 AC 76 A4 3D FC 1F 34 DC AB 7E EC DC 07 41 6B
 CD 70 65 5B 02 74 52 12 81 6E 06 51 2B 30 43 AE
 B4 19 13 31 A5 DC B5 9E C3 B3 53 D9 40 D7 84 AE
 29 0B 6A 48 9B F1 20 A6 08 5B F8 DD 6C 32 3E FC
 E8 03 46 BB BE DD B9 C7 27 6A A7 77 DE 01 48 AE
 81 A4 EA DF 0C EF 99 A6 07 1B C3 70 BB 3D B6 48
 3B 3E 88 9D C1 B0 98 AE 0C 1D 5F 27 C3 42 C7 19
 2C EF 2C 37 73 B5 58 61 13 C0 54 43 FC 1B 57 BF
 EC 0B C2 3A B1 B6 70 7B AB 73 68 97 36 C1 5C 72
 E6 DE 43 96 F3 D8 53 5F 62 24 AA 84 EF 26 0C 32
 F6 B9 E5 46 C5 6C 5A F8 DF B6 A2 77 13 A9 E8 1F
 47 2B E5 D1 F8 86 94 34 D3 52 BF DE 7A CB 00 22
 B7 C0 78 C3 D6 94 51 E0 4A 3A D5 95 AD 35 E6 79
 15 64 ED AC 14 42 7B 53 5D 6B D7 96 03 71 FC AD
 21 3D BB 0D 10 AC 45 FA 77 D8 54 C1 4B 87 F6 A0
 AC C9 DC 0F 44 41 DD 8F 61 2D C0 CE F5 C4 7C 50
 18 85 43 89 77 5B 93 EF AE 01 22 95 79 68 82 25
 63 33 68 3E 87 04 25 2F CE 71 9E E8 C9 F3 CA FC
 96 E6 93 41 A0 8E FF BD A6 71 6C 3B 7C 89 D2 50
 F5 20 7A 8D 47 DA 39 5B C7 06 9A FD 58 1C AF AF
 66 FC C6 C2 FE 15 47 14 3D C6 85 29 3F 70 00 A8
 8B FC 60 94 24 48 62 7E A9 F6 F6 C2 DB B3 CD C2
 DB D7 B4 06 EE E6 2F 04 4F A0 66 D9 F8 15 B9 13
 E8 04 0E 8E 6D 36 3D 74 CA D9 07 48 05 3E A6 DB
 A3 3C 63 86 24 63 22 67 48 19 A6 40 B5 BF 49 D0
 54 FD 52 36 93 4F BD 7D 94 6F AB EC 96 F9 FA 22
 8A FD 51 C5 18 28 81 3A CE 0C 93 F6 86 55 BF F9
 FF 24 D3 D7 65 41 70 0B F4 36 09 B5 82 8D 67 4A
 33 2C 76 02 C9 DA 23 09 DC 28 CB 52 87 63 4C 4F
 9B 0B 8E FA 30 9D 3F 7A B4 39 8C 95 71 C4 45 E3
 E4 C4 FC 7D 40 17 18 16 6A 26 A6 7D 52 32 02 63
 2E 10 59 79 AE D5 C8 27 2C 46 C7 D0 31 B7 15 7D
 69 A9 A9 3C EC 48 A0 E8 4B AF BC F5 C6 E9 F5 0F
 45 81 5A 4F 2B 2E 10 8A 49 92 14 E2 C9 09 21 F5
 8E D4 2B DA 76 36 81 B8 A8 B4 2E B2 4E A6 CE C3
 43 58 17 A6 24 AA 39 CC EB 8A 61 F2 51 D9 1D FF
 3F A9 79 65 52 81 A2 AE 8A CD 3E 35 7A 92 20 B8
 E2 D8 33 66 68 D4 3E 1C AF 08 B5 D6 17 F1 B9 76
 07 27 69 2C 66 FD 72 F9 45 43 3E CB 00 A8 49 E6
 DC D4 FD F8 1E 25 F2 F2 0B D9 F1 A3 FD 88 51 B6
 23 78 D2 C0 65 2B 13 93 D6 03 3E 46 C0 50 D3 3E
 43 70 3D 15 8C 41 40 AA C7 9A 44 F5 86 B4 DE D6
 50 3C 20 C1 E3 84 DC A6 F0 56 7F 32 91 FA 1D 26
 F2 F7 CC E9 D1 17 F4 E9 3B C5 F2 B7 D5 B9 36 B4
 02 53 D8 C2 E3 04 60 18 80 4B F4 62 3E 61 61 F1
 B7 8C A1 58 22 B0 C7 9B 62 48 D2 EE 86 8B 95 12
 E2 22 9A C9 CD A8 74 69 5F 4D F3 10 89 9F 38 34
 3C 02 AA F0 88 9F 10 08 D6 E1 64 65 54 71 1A 6D
 17 B2 60 95 2B 59 69 87 F9 D2 D5 7A FD 33 E2 4C
 CD 06 76 07 A1 67 78 D6 C8 6A 09 79 3D 5F 61 10
 7A 76 07 97 BA 52 10 CD 3D A6 67 34 61 C8 CE 54
 26 F6 4B D1 F3 F0 E4 D4 E5 59 63 A5 1B EC 4C 29
 F4 79 1F F9 6A 23 13 48 28 72 28 1D C4 6F C8 3F
 11 60 4B 88 BA 48 BB C7 F0 6D 67 EE 05 D0 04 F3
 7F DD 02 C4 A0 F3 E9 2E 19 87 3C 8A E6 9E 28 4D
 41 62 EF 3B 26 1C 1F 2C 4C 90 FE 60 B5 08 6B 51
 C8 B1 0C DA 72 83 8E 86 A6 AF D0 A8 FE 10 CD 2E
 C4 90 DB DB AC 05 46 9D 68 C6 7E C2 11 CB 7B 29
 FD 43 1F BD 39 11 24 9F E8 90 4A FB 60 ED 09 EE
 8A D3 ED 6C FA 52 CD 7E B6 86 30 37 8E DE 1B D8
 74 51 08 0B 51 AB 18 21 91 25 53 8C 3B FF 8D 7E
 48 7F 98 74 CD 21 F3 97 03 B9 A8 EE 1A D2 42 87
 22 C3 43 C8 ED B8 47 0B 3A 30 62 23 AC AF F2 F5
 61 F3 86 36 2B 60 08 64 5B F9 13 B6 1C 73 86 3F
 1B CC D6 29 C1 CF EF 7D FC CD 63 C0 1B 86 53 A9
 93 BC 7C AF 6C F8 89 0E 81 6D 8C 98 1D 37 78 98
 57 92 54 8F E9 C8 6A 9C 39 B2 C1 21 AC 08 4D 0E
 98 F1 05 4E 8C 60 D1 3D AB 4E 32 9D A8 B7 0E A5
 00 7B BF 66 51 DC 45 20 74 00 35 39 A4 05 BB 30
 AA 21 16 B8 4C 96 B1 05 83 34 4F C8 FC 30 0A DA
 72 B6 72 66 12 04 DF 44 8F 40 B4 29 B0 A5 85 A3
 CD 03 07 2F 5C CF 84 6E DC 56 EE 8F E5 31 A3 A3
 3A CD 80 7B 1D AD 8F 7A 43 7A C0 C2 1C E6 E9 77
 E9 8F 89 16 7E 82 7A 19 54 DE 8C A2 59 1B 5F 13
 D5 45 D4 59 43 27 82 53 AC 56 4E 7B 85 55 04 1E
 B5 91 79 D1 9A F9 F2 1C 8E C6 8E 2E 0E 19 23 66
 1C E2 D0 BA 10 31 32 43 D4 CA E0 C3 BB F1 E2 A9
 8C 0E 57 75 3C 7B 3C AF 97 09 0E 29 85 78 95 EE
 F7 32 A1 5F 1F 60 25 55 5D 18 50 AF FE 1E F0 F2
 E8 40 6C 45 E0 37 39 F3 3F CA 3F 55 D6 F0 B2 1E
 C9 AC DC 63 25 6A CE 28 17 3E DF 49 F1 E5 76 E1
 79 69 82 3B 4C 88 FD B0 3A AA E9 E0 02 6C 7D 6C
 B7 AA B2 51 23 9F A4 7B 31 53 79 DA B1 E5 2A C9
 22 80 61 28 1C BC 06 C9 F5 CA 6D 3D 91 94 68 23
 24 30 5F 88 20 67 10 D9 99 95 B7 CF AB D5 FF A7
 D9 E8 35 36 21 4C 90 21 05 BD 9C 7F 14 29 2F 39
 1E 06 BD 14 44 B2 F3 82 D9 47 7B 57 25 97 EA 9D
 F0 DC D4 0E 50 7F 52 2C 6E FA EF 25 67 2F 93 45
 A6 E2 C7 3C 96 5A 33 FE B8 25 33 FB ED 05 D5 FA
 9F A9 FE AF AB F4 7F F9 61 6E 87 D6 CE 18 AF 60
 A6 CA 87 E5 8F A1 80 6C 4A 20 87 DE E5 42 1E 24
 0D 7B 6A 82 3C 9F 50 46 EB 41 04 7E C9 F8 2A EC
 0F A4 45 A5 87 02 F2 11 DC 74 19 37 09 AA 5D 5C
 40 A2 E8 A5 80 5D 9C 89 0C BE 58 BD 7A 85 69 81
 AE 67 51 1C BB BD 14 B0 DB CD 6D D4 AC B7 6E F4
 61 C6 33 2F D0 B6 3F 59 12 31 EB AB 05 F1 40 17
 66 CF 3F 8B 3B 60 DE 79 EB 71 AC 3B 39 6E 6A C5
 A2 27 65 42 20 90 A5 8F 87 2C 0B 0B AD F8 24 27
 D7 29 CD 9C 75 87 09 89 73 1F 96 63 AF DF DB 8E
 91 BB 1D 5F C2 50 CD BF 8E 4D F3 F6 E8 83 FB 00
 35 08 14 92 9F EF 67 A5 CD A5 21 8F C5 16 F9 B2
 CA 7E 4D 5E 58 DD 59 2F 80 C3 06 56 8F A6 70 1D
 5F FA DE E8 91 40 59 9C 2A 53 DB 47 0B A2 E4 74
 F3 C5 DB 1A 8B 53 F1 96 0B A2 74 2C C5 AA 64 96
 E9 C0 18 79 74 04 38 B5 58 F5 4B E7 00 1F 6D 44
 90 83 B9 EA 93 9E 65 2A 81 E1 51 18 BA 97 FE 2F
 A1 B8 6B F7 CF 2C DA B8 17 BF E3 86 66 DD BC D9
 7E 97 2B 3C A8 3D FC B5 2F 35 F8 9F A2 34 53 0D
 1F BD 18 C6 C0 20 39 53 E6 50 A5 27 18 7C 33 ED
 F2 72 64 FD B9 D6 03 7C 51 EF F3 53 4E F6 93 E0
 4F A9 17 66 CC EA C7 2E 15 FF 48 9E 50 21 CE C0
 EA 52 BF BE A4 F6 0E CA F1 5B FB 53 70 E4 4C 24
 45 19 2A 98 39 83 62 92 F2 1A FD ED AF 90 AB 62
 6A AC 09 E4 0A DA ED CD A6 B4 38 A7 C5 0D A7 F2
 13 1A F4 91 57 8B C0 0E 09 6B 43 BA E0 54 F0 EC
 F4 67 3C E2 7C 00 FD 7E 01 AC 5A C4 B2 F1 29 F6
 F7 4A 50 F8 CA 96 B6 7A E6 AE 13 F9 8D 15 ED A0
 89 31 73 CB 0D 10 3E 1A 5A 1C 7C 6D 0B A0 96 29
 97 FD EE BB 41 8F 75 71 4C B8 96 E7 FD 0D 93 9E
 B1 F4 BD 20 A4 96 09 42 BC 33 12 7F 19 96 F4 C5
 FE 99 50 35 6E 85 55 B6 9C BD D6 53 FD 73 C8 09
 BB 58 2D C3 16 79 04 AE 20 C1 1E 40 9E 27 7F A0
 F4 6C B8 EF BA A4 BD 88 06 1F 90 34 5F D7 B1 08
 1A 31 6C 6F D0 8B 63 03 F2 AD C7 E0 6C CC 08 91
 FB 45 BF 4E 90 8D FF 58 D8 5F C4 3D B6 DC 59 0D
 7D 5A D4 88 F9 C9 B3 E1 EC BF 12 4F BD 16 67 4F
 07 BE 4C 7D 63 74 AF EB E5 CC 2E 21 8E 85 35 46
 F9 26 5C F1 E3 10 D0 08 A3 EE 6C 0F 5D 8A F7 85
 8D 14 C0 C3 D0 EC 33 37 26 E1 14 25 95 7E 0F 34
 5F 2B 37 A6 65 57 6C F3 A6 2D CF 8E C5 7C D4 5F
 0A C8 FD 0B F6 38 93 32 1C C5 AB 31 19 55 6C 7E
 66 35 01 93 19 AF 9F EF B3 54 2F E7 E3 3E A5 BA
 8B EF 61 DF 5B BA B7 70 9A 47 F0 76 78 B1 46 2D
 E4 21 01 BF 3C 31 1F F0 2E BA D6 41 D7 EB 87 1C
 86 AA 8D 9A CE F6 82 8E 18 81 5B 34 0D F0 33 45
 B8 F0 31 11 45 0A 4A AE 54 CA 1C 8B B3 4A A7 B9
 7E 69 CB 47 36 E0 8D 88 C6 B8 D0 CD 46 8D 2B 42
 0F 69 65 CD C8 62 BB D8 9D D7 09 01 30 D0 A7 03
 58 4A 44 34 ED 1B C8 91 37 A2 2C F4 0B 38 AB ED
 24 9C 05 7D 53 71 09 7C 86 56 94 EC C4 2D FD 04
 69 95 15 1E CF A0 01 D3 EB 29 24 0B 3D 13 3C E3
 80 58 29 FD 5E 09 64 90 6A BC 6F 9B AA 8F 4B 86
 90 C0 5A C7 C3 AE 4E B7 51 F2 A5 FE 7B 37 D2 30
 07 78 91 8B 80 B0 57 14 13 6B 04 AE A2 38 C2 F2
 68 D9 98 31 5C 26 E3 C9 74 0B 59 BA 70 98 EA 59
 D7 2D B6 C0 74 E8 4D 9D 89 A1 44 44 03 55 C5 6D
 B3 16 82 75 8E F3 AC 7F DC 07 5D BD 75 8E 1F F7
 83 61 C1 68 EA E2 2F 16 12 47 2A B2 FC 4C B0 4C
 C3 0C E6 BF AB 43 BD BA D8 90 AF D1 B0 85 AB CE
 8D D1 02 32 D4 17 9C 81 E1 02 9A DC 2A 23 DD 6D
 1D 06 37 12 93 66 59 43 3F 26 D3 AC 38 6A 56 AA
 65 82 51 92 93 9B 69 25 8F 33 45 84 B4 6D 67 F3
 DB CF D8 DD E2 1E 79 B2 F8 71 A4 68 E9 63 FA 3F
 74 CC C3 73 2C 6C 75 00 9C 5F 71 8E 15 68 24 D1
 08 28 D2 A7 0C AA 8A 41 4B 64 DA B3 94 52 98 68
 5F 80 88 14 28 23 D0 C9 DC B0 FC B8 C9 97 38 A0
 B7 BB E6 DB 6A 7B EA 3B 98 1E DA F3 C8 EB 9C A6
 5D 42 85 45 16 30 F0 7A 24 F1 0B 30 5E 29 D6 4C
 79 7B 36 FE 99 B9 46 6E E4 1F E3 5C 44 A8 63 EA
 86 E3 D8 89 FF 1E E7 C1 A9 F8 B3 FD ED F1 25 D7
 BC 4B E5 79 0B DF 4B 5A 5E 05 C4 F2 08 0B 21 52
 3F 38 B1 E7 08 CB 62 17 F6 D8 24 61 47 D2 15 AE
 68 81 D7 BB 80 6B 7F 63 2F BD 5C F8 44 AD 6B A2
 73 B0 D8 F2 4F C3 58 E7 C8 32 C2 29 C1 9E 78 34
 74 97 27 C5 95 59 8F B8 99 B1 D7 3D C4 0F A1 EF
 CC BB 06 23 DB 2D 07 81 80 66 63 A4 FF 16 5B 2F
 4D 22 13 F5 C3 20 0A E6 54 B4 3A 34 6C B8 4A 8F
 27 91 41 F3 FB 8A 4B 79 80 0E 53 9B 76 87 63 D4
 C4 B7 CC 3C C1 09 A9 6C 54 EB CA C9 98 72 66 36
 FD F8 AF AF 32 35 11 EC E6 5D 38 6E B4 38 36 BE
 6D 14 51 CC 50 73 C7 E0 C7 FB 74 C3 BB B2 D0 DF
 3D 6A 87 F0 C6 C3 03 9A 9A 8E 06 0E C9 CC 89 12
 85 E1 FE C1 C8 30 03 40 5B A0 32 D6 86 D2 CE 8A
 84 0B F5 EF C0 D7 45 FE 0C AA D9 6A A0 9C D6 D4
 6C 7A A9 EC A8 04 03 54 A1 B1 69 9F D3 0C 6B 3D
 0B 8D EA B5 C7 C1 00 20 8E E8 2E 70 38 91 50 0E
 41 05 FE B4 99 51 C2 C2 0D 0A 14 E6 80 B3 A1 42
 C4 F1 24 28 C7 83 63 8E 50 07 F1 DE 33 D5 E1 73
 CF 42 5F B8 F1 36 12 D6 15 FF 2C 97 22 52 C3 F4
 E1 2D A9 8B F0 A9 85 6A E4 57 7D B3 15 5A B4 5B
 96 68 68 F8 2E D0 03 5E 70 62 37 7C 42 41 48 97
 DD 6A FC 34 FA 2A C3 E6 60 A9 32 C3 92 85 01 4A
 E6 E8 8C 65 9E D5 09 F1 53 D2 D7 D4 1A D3 CC 8E
 60 F9 CA 2C 64 0B F4 3F 71 37 51 8F FA EB 62 23
 D1 9F D0 96 C6 B3 A2 40 F2 EE 83 0F 74 F0 0A 4E
 60 05 F4 A5 C3 DC AF 06 8B B3 F4 86 A8 85 1B F6
 96 AA 51 78 70 E3 6A A4 04 4A 7C FC 02 32 D3 0C
 B5 06 DE 54 26 45 FD DA 30 DF B5 AE D8 06 67 15
 68 AD F5 39 EF 89 F4 C4 CB B6 CD 15 16 90 16 D0
 62 66 7F 46 52 0E 69 02 69 31 D6 15 46 32 A3 32
 6C 2A 63 7B 1F 74 72 BA D5 01 4D 36 69 1D 77 C2
 54 11 BA 30 11 84 5F 5B 1A BF 00 99 7E 62 79 AE
 7A 14 C2 51 01 B0 AB F3 33 1B 34 87 02 98 9B BB
 BB 44 63 83 F6 31 F2 EB 03 81 8F A4 73 CF 24 40
 3B 0F 09 C7 5F 7C 6F EA AE 88 70 B2 38 03 A1 6C
 79 32 38 ED 0D B1 66 3B 65 18 16 91 89 01 FA DC
 53 D0 FE 11 F6 B3 A0 EC 93 28 6D 67 DE F9 07 5E
 CB F4 7B C1 8B E3 7A 3B A0 B6 C1 F1 FA 20 F8 E5
 26 B4 55 5D 10 47 16 37 30 1B DE 3F 59 98 B0 B6
 EF 0E D5 85 94 45 E6 48 CC 85 D3 84 8F 73 DB 50
 65 75 D7 32 4B D8 F3 5F F8 FA 8C ED 44 09 0F 66
 B6 C1 5A 8F 30 40 21 25 2A BC B4 7B 05 24 34 D8
 82 28 66 35 A2 68 74 40 46 C1 50 28 2F 42 C8 49
 C1 0E EE 26 F6 10 C2 01 16 2C 74 A8 D6 0F 52 A5
 D1 41 D1 4B 6D B6 1F 61 11 12 C9 D4 A1 7F D0 D3
 D0 E4 D3 DE 5E 8D EF 47 D1 FC BF 3E 30 85 D0 1C
 CD 87 44 0B 15 81 DA CD D4 09 03 46 C8 99 25 F3
 1E A9 49 83 9B 99 7A 1B 89 67 A3 04 5A C7 4D DE
 BA 9A A9 52 85 AE A9 52 02 3D FD 6F 05 28 9B BA
 2C 2A E8 95 BD F3 97 49 E7 C2 02 D2 3E 3A 23 A2
 CF 23 57 3A D8 D2 99 BA 9D 57 2D C3 26 31 9E E2
 98 CF 0B 9B 3C 8E 7E 28 AA B9 A5 47 52 31 49 F3
 E2 62 D3 B3 1A F8 44 EC FF D6 B9 8E E8 4A E2 80
 56 BF F5 E9 76 F4 6B 7E E6 96 18 18 0E AC 27 E5
 05 8F 8C D7 44 35 46 BA 6D 69 5C 4B 5B 4C 8A 15
 2F 81 50 66 B8 CD B8 07 D2 D7 48 D6 D0 F7 D9 47
 89 35 E1 84 B7 A9 DF 2E 15 9A 8B 1E 5B 06 14 67
 D3 6E 36 13 16 50 C5 37 AD 3F 1A 27 DA C9 6A 1E
 8F EB 4E E6 B7 55 A2 7D 89 C1 0F 03 C8 03 FA 23
 65 C1 FD 0B 42 74 8E C8 98 FE 37 70 1C EC 15 6A
 DA C9 18 03 21 C1 66 B1 49 61 B5 FF 8B 5D 09 DD
 A1 23 87 F1 80 92 89 3A 13 7B A6 DB 32 CE 45 06
 39 6A C1 83 EC D1 8F 8A 3A F2 DC 5A 7F F2 73 63
 B6 34 BF 26 DA 81 81 C5 2C 40 B8 CD 63 88 51 AF
 9D 46 2F B2 E2 32 58 95 5D DC 69 8A 7E 62 64 8C
 08 2A E0 F5 19 74 20 47 59 24 E1 7F B9 9B F5 50
 64 25 57 E2 6A 9D 9C CC FE 5B 79 F8 DA A1 2D A6
 67 47 6C DF A9 F2 43 12 6A 9A 60 71 F6 09 A1 96
 E4 AB 6D AE E6 A1 FD DD 5E 1B 51 C4 02 9C DB E4
 08 F2 91 F7 22 B6 4D 76 E2 1E 91 4A A2 6B 7A 2B
 37 67 95 A5 C1 70 CE 9C D7 CA 59 73 83 6F 5C F9
 02 F4 AB 18 05 33 7B 4D C0 28 6A D9 70 36 B5 DF
 54 60 A2 21 39 AA CA 92 46 08 09 88 4C F3 93 08
 FA 5C 8D EB F5 94 ED D4 AB D6 AC 35 6D 92 37 2E
 FE C6 17 92 07 FE B8 31 F7 2A CA D7 47 3F 74 11
 8A 06 E6 FA 39 99 8F 6A 24 FA CD 82 A4 A0 42 00
 28 E7 A7 61 86 68 D4 48 47 D9 4C 4E 32 22 42 48
 CD E1 56 7C FC 20 02 BC D9 1C 5D 54 1C ED D4 23
 20 68 6B DC 62 17 B6 62 8F 13 E6 21 7D C3 6E 8E
 4D B7 D4 EC 2E 81 E5 A6 FC E8 62 BB A6 05 D6 4C
 4B C1 56 BB 7C 0D 7D 77 51 9F 0E C5 59 D9 EE 53
 7B 19 AE 4A 03 7E E3 6A 1B 3C 98 92 0A FD D3 66
 64 90 74 5F A2 BD BF C5 24 2B 8A D8 24 65 FF 5D
 E1 6B EA 66 3B E2 B8 22 CE 4E 58 2B 3F 1A F6 5F
 46 5F 7A 02 D0 E9 8D 49 46 57 88 4F B8 B2 CA 0C
 AE D4 DA CE FB 55 AC 7F DD 01 40 90 CD 79 8C DF
 E8 5E 58 90 C3 42 3B 31 30 28 AC 3F D2 F5 B5 2C
 11 55 39 CB FD 12 70 00 C9 5B ED FE 67 CB 95 63
 11 87 A2 5B 90 6C B9 45 8C 2D 4B B2 24 39 0F 23
 48 0B A9 C9 25 58 11 D2 E7 BC 3C 8C 5F 5C 7D B7
 05 F9 B8 2D D5 DD 79 E1 6C 57 63 77 F3 81 07 D8
 6D D2 FC B9 7D 5C 0D 43 EF FF F2 81 07 04 37 3D
 7B 4A 52 DD 97 D6 C3 E1 CF 9E 78 39 39 6F 6E D1
 0A 8B 0A AF F3 BC 8A 61 C3 5C 0F DE 30 B8 66 1A
 69 D1 C1 37 15 9A 72 8E F3 F4 B1 41 2C DA CD 60
 99 9A 1D A5 93 DC 83 90 B4 C9 39 23 7F 79 4D DC
 FA 3E E0 F5 F1 06 46 FC FB 0B 4E A6 C2 55 13 1B
 0A 7D 2F 0B E9 9B 2E 13 A7 FC DF 34 5F 4B DD 32
 D0 41 81 ED B8 B3 97 6D 8D 48 FE 03 B7 2D 3C 80
 E2 86 AF 42 C0 CC D8 40 1A 1E 5C CD B6 1C 18 F9
 F5 1A EF 37 A6 F1 79 FC 5C 0F EE 7A B8 E0 85 65
 DC 15 08 9D 47 F2 6A 80 B5 12 E1 FA 54 10 D1 15
 A0 79 24 6D 91 F7 2E E0 B2 D8 0D 5F CD 89 40 2B
 3B D6 B9 34 33 0D 19 70 2F 0E 54 A6 65 07 EC F4
 9F EB AA A8 77 15 69 89 EE B4 0A A7 87 E0 4C 93
 1E 93 D2 1D B0 74 0C 12 4B 39 39 71 5D 91 ED 80
 52 99 A1 85 60 B5 48 7B D4 68 11 8F F0 F4 AF 25
 6A D6 B1 A9 DC E2 7E 00 6C B2 E9 FD 21 B0 F4 5C
 8F EA C8 84 00 13 F5 46 9B 7F 22 FB 30 24 F7 87
 F6 5F AD A2 C5 16 2B EA 4A 01 CD 37 22 F6 36 A4
 14 84 76 8A C9 EB FB 44 0B 61 CC E6 0A 74 A5 E1
 12 65 6D 19 DD 12 C1 3D 15 BF 18 98 91 D0 0F 84
 8B 9D 51 C2 44 4E 7E 82 F6 23 00 FF 9C 80 DE 1D
 62 FF 47 30 8A 9B 27 54 7B 98 C3 BB 34 2F 1D 9D
 B3 28 FF 2C 8F C2 92 9A A1 9D 00 A2 BC D6 4F 10
 31 60 4A 78 1E 45 EA 81 09 1C B4 A6 0F 4A 6B B5
 95 06 09 83 08 44 E6 1C 6A 03 B0 C4 B9 CF C9 C7
 E8 78 9A 49 70 3F 7F 3A 50 6E D4 60 B8 6C E8 FC
 8C D8 41 42 51 31 36 6F 11 12 16 C1 A0 98 ED E4
 56 6B 6A 2A 7D 21 69 F2 3E 29 FB 66 1F 3C 3D 4F
 F0 2D FD 57 F3 9F 0C 97 0D BB 05 2D C9 27 4B 6C
 C2 AC DA C2 9E 93 B7 84 DC 74 08 A8 49 5D 3F 94
 FD 6E 07 63 5C CC 21 EF 65 AF 93 ED 4E 60 50 00
 26 79 2D 1A CA 5C 99 BC 38 88 72 61 F2 8D F1 CE
 2C F9 29 BE FB 88 A9 73 C4 18 00 5C C4 4B 4B EC
 E7 3E C8 31 E8 0A 55 9A 99 B7 43 68 42 19 85 B0
 04 7E 93 22 FD 37 17 D7 76 E0 3C 16 CA 71 EE E5
 EC A9 98 22 A4 D7 6F 78 6A 06 B1 20 96 D7 0C 55
 BE 8E D9 44 8D 33 35 FB 82 AD A6 5F EA 54 7D 11
 4C CF 89 53 CB 02 93 FD 45 17 1C 13 59 7B 63 2F
 42 C6 09 4B 9B 86 06 88 34 57 B8 66 84 F8 71 F4
 0C 46 DB BE CA A3 C3 DB A4 8D 8A 47 6D 65 AA B4
 7F D2 60 40 61 63 86 AA 1D 6D EC 70 CB 44 71 33
 F3 B0 92 1D 43 63 A4 15 AF 72 06 99 E8 36 FB 0A
 97 27 6D 97 F4 AC D5 16 7B 32 67 F0 8A A9 0D E7
 38 37 97 F2 A4 A0 63 40 DB 8C 9A F9 47 D4 6F E1
 1F 43 E9 CD E5 B2 52 BD BD AC 87 B8 CE 45 B4 7B
 AC 77 11 F6 96 9E A2 0D B0 9F 19 04 32 4D 18 2F
 E9 91 40 18 93 77 CD A4 2B 2E D6 1A 03 8C FF B5
 C1 B7 83 D0 B6 59 3C 76 9D 4B 8B 4D A1 40 59 88
 70 B8 27 34 79 79 95 B0 4B 41 09 A4 48 BB 65 22
 C2 E5 3F 3D F0 8F 2F 46 FC 4A 6C 81 61 27 0F C2
 51 56 14 EE CB F8 70 9F 5D 1A 15 6C F8 82 9E 38
 D2 94 66 D4 87 3E 5E 96 19 B5 09 8B 97 B6 E1 5F
 C6 AA 8C 06 39 63 A6 D1 15 B0 0B FC AF 96 46 54
 F6 9F 1C BC 78 76 ED 7E C5 5F E1 A1 F7 D0 86 51
 80 00 DD 72 5E 8C 07 47 A5 83 02 A7 89 AE 02 0B
 50 EE D0 13 98 CD 22 6D 52 43 CD BB 8B D0 0F 9E
 A6 CB 89 02 C8 A6 FA E1 69 56 CB 51 A4 87 8E 3D
 A8 AA 69 63 33 CF 00 3E 12 7C 7B 7D DF 45 86 F1
 1E 24 5D B2 5D AD C8 FD 9E 95 F5 B6 58 4B 88 4F
 C2 42 1B 71 70 91 73 8B EA F1 1A 9C B0 B6 30 92
 76 CB FB 31 53 89 6D 08 D4 CB 84 65 A0 4C F9 B0
 A8 0A 7F 6D 8E 09 2F 98 90 A4 05 65 9D C8 AB 45
 7D 16 AD 83 DA 6F FD 2C 7B 87 5D 8C 8A 13 DC DB
 A1 AE 6B 19 4A D7 82 09 38 96 CC 8D C2 A0 6B 3B
 F5 24 D0 90 01 4F E4 23 C9 94 73 E5 BE C7 A0 9F
 90 94 A8 72 A7 47 B6 8D 6C F6 FA FE 86 FA 39 10
 21 C4 29 40 6F 0D 63 C6 78 12 2C BE A1 51 B6 43
 3E A2 6A F7 9B 51 AC C7 17 A7 41 6C 98 76 B5 31
 CA 28 E1 22 30 FD EF 73 69 1D 95 4D B9 A4 F9 A3
 E0 13 9A CE 44 8B 6B B8 A0 CF 3B AC 4D 0E 42 0D
 6A 4E 56 46 B0 D8 16 87 3A F0 3B 9A F7 A8 FC F2
 E5 CB 83 02 19 21 E5 B4 E7 07 91 E3 D3 1E 5C A2
 A8 B2 7C 80 FA 23 75 BD 92 50 BF EF 89 25 1F EB
 6E 04 22 11 02 69 6E 64 53 6A D4 FD 7B AF E6 DA
 BC B1 73 77 6D F1 5A 4B 2B 87 72 14 00 8A F6 AC
 AB 3F 1E 27 D8 C7 0E B4 FF B4 45 9F C0 1F AD 42
 22 A2 AD 55 EB 3F 15 B6 A3 C8 14 C5 C4 35 41 4C
 ED B8 A2 EC A6 FD DB 7F 65 20 31 FD 62 2D 4B 79
 4D 63 3C 8B AB 05 93 68 97 E8 9A 3D D6 D1 54 91
 B0 95 83 D5 5F FA E7 81 C9 0C 0B 95 C7 CD ED F9
 2E 7C 1E 4B B1 A4 86 93 5A 18 9F 19 6C D2 09 77
 8D 24 94 75 98 D8 AE DB B2 10 88 24 1E FB 29 27
 82 8B A2 57 92 F8 98 B1 9F 76 C0 27 6A 3B D5 B1
 6A F0 FE DE 11 4B 52 4F 86 D4 E0 1C F4 D9 67 C9
 D1 41 9A A6 F6 D3 B7 09 1E 6C 39 9E 8E F6 D6 BB
 35 8E 98 62 E9 F8 19 64 9F 41 78 57 FA 12 0C C7
 D5 FD 1F 2D 69 F8 81 C4 2E 20 33 45 5E FB A7 FC
 1A 9B 58 8D C2 20 54 6F 5F 1B A1 E1 E4 22 D5 6F
 83 BB 0B C7 D2 C7 9C 18 9D 1F F8 C5 32 1C B0 31
 54 DB 7E 76 23 7C B6 E8 6F 03 D4 DB 88 2F 80 81
 D1 49 2E CF F5 C9 B6 8E F9 A2 63 52 23 82 38 13
 C2 44 91 25 BE D0 81 26 35 83 93 AF CB 08 10 9F
 1B 75 1C 7F 1D F4 52 E9 19 16 AB E2 4C AD 3D 00
 DF D6 05 F4 9C 93 07 F3 A6 BD 8E 2F 9E FA ED 41
 9C 82 12 9D A6 90 22 8A 7D 68 4B 25 3F 88 5C 49
 6B B5 96 6C E8 3D 07 67 11 AE 0D 03 3A 08 D6 F6
 C2 53 A4 63 D1 04 C0 D5 53 92 F1 12 0A 2D 0B 89
 79 E6 E6 A4 21 88 51 B6 E9 FB 30 F0 6E E6 44 B6
 1F 1A B9 57 57 84 7A 9C 23 6D 74 98 9B E3 7B 5F
 B2 A1 19 7F 2E F6 0B 1C 61 43 F3 CB 6B 60 8C 85
 1E BD FA 45 7B CE D9 CF 5C 08 26 84 91 E6 08 7A
 0A F0 2F 18 6E F3 D6 CC 25 D4 43 41 DB CF 33 77
 0A E5 16 AA 74 99 51 4C 1E 82 12 3F E5 83 66 B7
 4C DD DB 3E F8 1B 2F EB 75 D6 D8 9E 30 BE C0 35
 67 11 91 20 95 30 26 78 25 19 96 26 F5 11 B8 2D
 97 6B 94 AD C3 DF 55 C8 99 72 0E EA 78 A1 AD 68
 17 21 79 9D 89 80 7F A3 EF C3 BC C3 FF 9E 93 BB
 2E 83 0B CB 3B E5 85 BF E6 AA 89 3C 8B 7D B9 3D
 2F DB F4 62 7F F3 48 EC F1 8D 49 F7 8C C5 0F F1
 FE 90 CF 85 1E 71 0F 4E 1E D4 F9 60 3F AB 3D 1F
 FF 85 2F 47 74 53 51 AA 48 C0 ED E2 94 FC B8 57
 5E CA 89 7F DC 42 3C 16 62 3C 6D 7A B2 53 A4 13
 BA B8 6A C9 3A D1 D6 50 15 27 1B 1B E3 87 0D 72
 8C 20 41 B3 B9 AD E1 CC 3A 39 D8 A3 29 D7 FE 3C
 B5 75 C6 DE 69 90 AD 5F 4E 61 10 E5 F7 53 99 7E
 88 40 F4 38 1B 2E CF 11 DE DA 94 8A AF AA F0 22
 93 EC 77 9E AD 04 F3 E4 71 E0 57 1F 8B D1 61 22
 97 27 95 CA FF C6 12 34 59 7C FC E5 65 E6 C0 D4
 49 74 9E 97 D8 8D 32 0B 3A 87 43 69 8E 43 9A DA
 5C 89 D2 1A 3C 22 08 B9 68 B5 74 7E F8 F7 D8 4F
 51 B7 3A 0D 00 13 B3 71 F5 5D 1F 1A 83 40 40 CB
 E4 6C 04 F9 98 77 85 D9 C2 3C 17 50 4E 33 DE 54
 B7 C4 09 1A 6D 08 30 51 33 A8 E2 63 7A 2D 65 1E
 C8 B0 55 FB 81 25 3E D6 BA 6E 7B BF BF DA 26 48
 E6 CC 3D AB F4 68 B3 AC F9 6F 90 DF 8D 60 BD 7B
 05 37 82 0F 1B 48 AD E2 78 8B 12 DA F4 63 30 70
 A7 3B 59 39 67 DF 35 5C 73 42 1A 63 18 42 72 78
 D7 E2 00 14 8F B2 39 61 21 E6 1D 59 EC 7A 5B B0
 2E 86 07 D9 4B 51 A8 C6 F6 76 CB 4C C8 A2 25 EB
 0A CE 51 C6 CD C5 27 7F 60 B7 2B B1 F4 DA DC 5A
 AE 5D 7C 32 C5 19 DF A7 7A F0 F4 54 3E 15 FD 48
 A7 BD 0A 11 6D D3 5E D2 8E 81 C7 6F D9 01 26 42
 F7 A6 9C 57 10 DE C7 0E 7D A1 6B 40 B9 C7 BE A0
 2C 41 EE 27 32 D9 8F 91 DB 9C 8F 1F F5 EE 9C 98
 EA A6 04 81 B5 EA 12 C0 75 8D FB AE CE 1F AC 05
 CA 87 18 1D F1 F2 EA F1 99 89 E9 A3 CE 38 ED D0
 D0 56 36 B2 E1 B5 72 41 E8 58 08 AB E8 0E 5F 94
 B0 37 3A B9 30 10 33 BC 24 59 1D 33 63 B8 88 2F
 63 B9 47 B3 C2 72 22 2A 02 10 33 2C 8D E3 5A 73
 A2 6B BC 61 31 71 10 9F 64 C5 92 B8 B9 21 91 E2
 0F 95 18 46 84 EE CE 1B C0 71 94 B6 95 13 3D DD
 72 39 BE 18 6E 56 4E 0D 45 60 22 23 5D E3 C8 ED
 87 3F DD 46 3A 40 2E E1 90 D1 20 35 44 8E 87 9F
 67 95 47 6C 7C D4 B6 7E 24 10 FE CE 2A 62 8A D5
 05 8A C3 77 62 1F 2A 69 76 E3 EB D9 10 FB F9 F4
 B9 9A 95 2D D6 6A 72 E6 8C D2 3A C9 DD 72 D8 D6
 FB 56 DB 85 7A 4A A7 D0 0B 26 52 43 EB 0B E9 F8
 31 AE 14 D5 06 8D 04 A1 E3 00 FB C4 DC 58 5E 41
 68 D2 A3 32 3E D0 88 85 82 8A 5B 20 0D 77 6C 9A
 22 42 52 1F 96 6D DD 8C 7B 4D 5E FC F6 1B BA 38
 47 3F 17 C0 AD 88 C9 1F 9F CB 26 B5 86 08 13 C3
 4D D3 B3 81 EC 37 03 F0 9B 5C 2F 42 4C 04 9F F4
 49 80 EE 3B 3A 14 B6 E8 9F B1 86 50 A6 8C 69 79
 FD EC 6B D0 81 62 06 EF 0B 58 26 55 48 AA A0 D5
 5E CD C8 D2 B2 D0 DC 6E 12 EE BA 74 F4 2D 69 EC
 44 99 1F 31 F1 06 FE A2 F5 2F 0D 98 0C 3B 1E 02
 0E 22 9A C3 D1 79 37 D5 AB 20 9C 6E 95 8F 49 E7
 A7 FA 96 E7 33 2B 74 24 4E E5 D4 0E 3F 30 BE DC
 8B D5 22 E2 EC 1C 5A 3D 70 F4 A1 DD 02 6A B8 74
 0F 15 FC 89 83 57 72 3C 7D 32 ED 85 70 7E C6 D5
 B9 E2 81 31 D9 3B F0 9F 3B F0 97 44 1F 3A FE EF
 75 A6 43 09 11 D9 27 0D 36 AB 92 E0 CA CF F0 66
 B2 74 56 63 9C 23 49 2E 58 83 C3 F8 A6 89 F6 75
 B7 11 EC FE 02 CD 7B 54 21 30 06 51 ED 3E 7E 86
 CD 07 64 A5 AB 63 DB 09 1C CF 67 09 A7 8C 85 B2
 E1 20 AA FD 76 8D 75 20 19 11 6D 26 28 4E A2 3B
 93 DF B9 7E 92 3B 4D 7B 87 E7 B6 2B 58 5D C8 E9
 27 3B E8 6B 02 5F 41 1B D4 BF 21 69 BC 2B 12 D7
 E4 AC DE B2 05 9E 49 C4 F4 D3 F7 73 D1 14 84 88
 86 E6 85 EF D8 A7 69 BA 7E 4F DE 6C E5 1E F2 0E
 FA 56 ED 21 31 98 20 4D DC 9C 06 95 64 C1 E6 23
 8C 22 99 93 BA F7 F8 17 FD FE EB 3B 96 FF 78 D9
 2C 0D 7D 61 AD 97 EA 1B 77 E8 BB 87 03 5B 2D 3D
 28 8A AC 6D 50 D8 F2 98 FD EE CD F7 72 BE A5 B9
 51 92 F9 55 3A 7D 9F C3 1C 33 0A A7 C4 3E F1 10
 F2 F6 82 3B 26 8A 78 2C 87 CA 25 B0 52 77 4F 66
 33 39 9B A8 56 B1 35 15 C3 45 76 6D 2C EB 7A 60
 D3 60 21 24 A8 D7 16 7C A7 02 55 95 69 6A 81 D2
 87 3E 16 E4 5D 4D AE AF 04 BD D0 CC 7D BE 35 6F
 C3 4E 8A 27 9B 2C BE CC 1B 66 33 D6 56 7F 18 1A
 62 77 A8 DA 8D 5E 77 A9 58 1B 07 74 0F D1 60 FF
 03 53 9E 5C EC AA CC 1F 8B 05 72 0F B4 D9 C0 BC
 21 DB B7 E7 8A 98 C0 9A 87 59 72 F4 54 CF 4D 18
 62 16 A1 E0 8B A8 77 C2 E2 E5 62 4B 54 08 E2 8F
 68 55 5B FA E3 26 18 C3 45 3F E9 99 A8 02 38 CC
 94 7F F0 8B C9 41 52 FD 97 85 48 B9 3B 65 5C D0
 2D AC 91 66 E7 3D E8 11 C0 70 CB 4B 2B 5E 2E 47
 DD F0 5C 83 11 82 31 50 8E 51 B3 22 98 ED 72 A4
 B6 A2 7A CF 46 48 F2 55 4F 93 FE 6E 85 BC 86 7B
 92 28 52 4A F3 8B 87 8C 0B 60 7A 26 47 B8 D4 1D
 EE 0A 66 9D 51 06 D5 19 ED 3B 48 A3 10 EE D4 DB
 56 13 7A 01 52 BD 4F 6B C5 5B 69 22 41 FF 88 F7
 42 62 14 7E 59 8F DE 2A 2F 0B 22 DC 43 F8 AF CC
 CF 6C 23 FA 16 5E BC 92 FF 55 EF BD EF 43 83 8E
 B6 D8 C7 60 75 3C 9C 35 4B 71 F3 82 B7 89 E1 6D
 AF 21 43 87 62 16 49 D0 07 81 EB 07 B7 99 F9 23
 B3 1B 14 15 36 F7 74 6B 44 CE CC E3 76 BA F3 9D
 C2 FF 07 6F 2C 08 A5 4F FA 58 4F 81 3C 3C 01 B8
 08 86 71 15 C1 A5 80 D3 56 E1 E5 5C B9 3B 03 C4
 B6 11 1F DF 80 34 41 8A 28 52 AC 7C B0 B8 1B 1D
 9B 71 EA A4 AB 5E EF 2D FE D6 B8 6E AB B9 8D 44
 11 1C A1 33 EC E3 97 AA 77 B7 D0 01 D7 C3 44 B8
 FC 4E FB 9A 6A 2F 66 52 1C 39 CC B2 E0 74 67 1E
 9A BE BD A2 CC 09 BA 1D A6 40 B4 AE A8 71 C1 3E
 EA 58 02 7A F2 E5 79 B7 6D B4 55 DC C1 96 46 99
 9B 67 D9 BF 78 94 80 4A 7A 46 72 61 3D 4C 25 47
 E7 F6 4E 5A 4F 18 B7 98 ED 4E 2D CB 41 1A 4B F2
 BB DE 1A C4 B0 D3 D1 54 D2 3D F9 69 46 5D F6 E9
 B8 1F 25 D0 71 74 5D BD 6A 2C 43 F8 B0 4B B3 B3
 E2 DA CE E4 C4 9C D3 1C 3F 10 EB 84 8E B9 07 30
 98 0E 9C F8 3B 31 19 36 C2 B3 3B 29 2F 96 39 44
 9A 60 63 C1 BF A0 00 C1 00 5B 35 CF 56 77 EA ED
 AE 3C 7B E7 77 99 47 28 2B CA 5F 47 8F 6C 38 2C
 53 D5 80 77 55 3A 32 E0 7B ED 2B 77 5B BE 68 41
 E4 98 17 BE 74 6C 90 50 4E 65 A2 CC 9A 96 45 07
 EA 87 18 61 8A BF BE D1 84 7C 71 81 D8 A8 26 23
 BE DA 4D B3 79 4B 37 C9 33 20 53 DF 2B 6E F2 B6
 B8 4C 63 E6 F1 0F A1 36 56 FC 80 E7 E0 0A 66 3B
 25 D6 AF 2E 0A 3F 45 09 D3 9C 00 D1 10 47 70 81
 41 10 CA 1C FF C9 E9 29 C6 D0 3F 8F A1 23 78 15
 76 FD 9F 77 F0 98 F5 42 89 95 AB EC 2E 04 F6 2E
 45 03 0B 92 5D 32 DD 20 C2 BE C1 76 EC C5 5B 0F
 CC 0C D4 30 EE AC 53 08 57 E8 74 70 AF 31 DF 26
 9F 7F 80 95 DC F2 59 63 A1 E5 07 CD 61 C9 4A F5
 C7 F0 99 C8 D5 65 14 4C B2 F1 B5 53 43 D6 8F 94
 F9 41 48 FA 03 FF BB 1D DA AB 75 2D E6 EA 7F 5B
 07 33 1B B4 C7 89 1A 65 CD D0 40 2A 1B D6 4B D9
 6A 79 7B 7F 55 9E 65 A1 22 BB A6 4A CB 4A 9A 3F
 C4 68 9A C2 86 2D AE 4C F9 16 72 E1 A8 2E 92 98
 18 D7 4B DD 63 E9 A3 57 EB 0B 21 47 E8 05 7B B0
 8B 90 C0 DE 79 9B AE 34 9C FB 79 A0 B0 F2 AB EC
 E7 51 F4 4B A2 D7 8C F7 47 6F 9A DB 18 25 43 C5
 2A 11 B5 01 FC EE 6D F1 2A 3F D8 53 FC 30 9D EF
 4B CC 7E 3F 27 CB 78 D4 C9 08 D5 DB 84 42 DA 59
 E1 FD 93 6F 42 88 72 79 89 72 34 4E 86 4A 35 89
 6F FC 4B 5D 29 8A D6 11 01 C9 F3 27 E3 2D 50 0A
 59 E0 BD 22 DA 1D 67 EA 09 89 06 71 03 04 5A 4C
 70 CC F4 AA D1 09 8B 4E 0E 64 96 83 76 BE CE 32
 7A 5E A2 9F 1B 20 B8 12 6A 98 59 1F C2 BD 23 D5
 B4 BA 01 C8 0D 8B EA 04 62 EC E8 B3 A0 15 F1 A2
 4C D5 2C A5 41 BF FB 72 40 75 8D 25 57 51 E8 BC
 40 0E 3B AC F8 3F 4F BE 05 1D 49 87 CF 5A 35 F5
 A4 31 13 73 DD FD 74 46 A0 EE C1 86 F5 B2 0E 0C
 05 1E 49 06 F0 D5 FB C8 C5 96 32 38 F1 23 4F B8
 FF D3 3B 9F 17 DF 35 0D 55 FC 25 20 86 3F AA B3
 D5 7F B9 43 ED BE 5F 39 34 B6 C3 04 59 6E 91 66
 CC 58 84 87 89 58 48 67 D4 61 2A FB A9 EE 5E D7
 82 E4 ED 95 B3 9F E3 1A 8B 4F ED 0B 06 79 EF BE
 52 EE 24 BF 6A E3 5A 2E 08 D1 86 86 B5 E0 77 39
 C3 EF F1 5B AC 0A 3C 06 B3 70 EA 89 61 A6 4B 7A
 96 C1 CE B9 58 F4 D8 E6 BB C7 9F 62 31 CC F2 60
 6E 53 AF 5A 76 04 C0 44 F1 56 D1 2E C0 57 94 3E
 D4 F4 EA F8 B3 59 30 FF E1 B3 C3 DC D9 68 F6 A5
 7C F8 36 85 51 C5 F5 70 B5 7A 04 5B 8A A9 F6 A1
 5B C6 B6 60 76 E9 57 26 F9 C1 F8 78 4F 83 8D C5
 C2 D0 30 BD 4D 50 9F BD 63 A9 FD BE D1 3F E4 1A
 47 F6 64 A0 53 B1 71 83 85 76 ED D0 C0 EF E3 0D
 F9 F8 50 8C EA 3D C2 1A 8C 19 F3 55 90 F0 10 6B
 4E 1C 30 1C 51 E8 9B C2 75 DF 69 65 5B B8 6E 1D
 39 96 7B E4 95 7F BA 38 16 84 37 FE 33 B3 A1 D1
 FB 17 0A 5C 21 29 6E 24 B1 A5 AF 6F BE 45 0F 34
 40 19 85 C8 20 FF D6 DC BE C1 8F C3 AA 78 96 44
 F2 E5 6C DA 2A 99 35 A2 EE BB FD 93 90 76 FC D7
 09 AC D0 2C 01 06 9F B7 E5 DB 3C 4B F0 0C 0E 3E
 9E B5 13 D6 F4 F3 E7 B8 3C DD 23 2C 5F 15 BA 38
 01 DC 7D 82 49 D3 BB 47 F7 D4 FC 4A 10 A0 CB 4A
 AC 1A 47 C7 A2 6A C5 37 07 61 D9 A1 D3 70 F8 3E
 AA 4D 07 83 3C 31 1A 4B FC 01 70 F0 4E 05 F1 93
 98 50 12 E6 2F 26 B3 CE AC 9C F5 A3 51 28 39 0D
 6A 71 07 D3 08 5D 2F 91 09 0C C2 0D D8 C1 74 56
 67 14 39 D0 6F 26 5D 48 F5 0F F5 1E 4E 36 7E 08
 2E 4D 96 DE 2D 63 53 AB 52 61 D6 D3 59 CD 02 FC
 85 B0 70 86 37 0A 60 9F 50 E8 61 0A E2 3F 82 B3
 78 11 D8 07 38 E1 CC E9 43 7A 87 8D 0D C6 1B AE
 55 56 84 DD 41 B6 C5 59 80 38 BC 3C D6 BD B6 1D
 62 DD 41 3C CD 18 10 B6 60 C7 FD 45 CB 1A 39 EC
 9C 6A 19 F3 76 91 87 33 3E 51 68 F9 42 8A 7C 97
 DA 20 2E E3 49 04 50 56 32 4A 44 C6 42 65 61 FF
 24 C9 5A 4C 9A A2 B7 E9 45 99 9E C2 A4 46 7A 74
 AF 12 08 70 E7 D6 FA 6F 0E FC 6B D4 5C 04 F7 CB
 3A 29 8E 66 A7 EC 5F 55 30 B5 7E A6 55 6F DE 6C
 F2 C6 2D 20 09 BE 19 C0 BD B0 57 7A 21 FF 7A 47
 5C B5 CD DE A5 FF 31 77 33 67 60 DF 2C B1 DC 84
 9E 14 E9 0E 08 43 2A 0D 91 F4 57 12 0F 2C 45 96
 57 8B 28 C3 87 1A 2A 0D BA 61 4D 60 32 35 3C AA
 30 DD AC F3 7B 9D 8E B6 4C 96 91 A2 B7 6E 59 CB
 64 6D AE E9 06 73 18 AA 38 9C 45 DE 32 02 88 A3
 D9 94 5D AD BC 57 85 B9 B9 24 C7 36 58 53 86 CC
 FB C6 93 08 C8 84 E9 6D 34 E4 F9 5A BD FE 44 CE
 3A 7A D0 A4 85 E7 EE D5 55 0E 5D 9C C5 20 A6 B4
 6C 71 1A 55 59 6F EB 03 1A 4E 62 C5 6F 9A 26 CA
 42 0A 85 36 BF 57 41 F7 E8 6B 82 49 01 BC EB D4
 25 C6 C4 DA 8E 85 00 88 8F 02 0D DC FA 6F CF 11
 EF 70 F9 BC D5 0F 00 FA 7D 88 C6 63 AE 72 D8 99
 EF EA 8D CD D5 80 84 1D 26 24 C5 85 53 DF 8D 18
 A1 CF 9D 7D 16 F6 B7 10 1B 80 3F 39 3F 5D F5 D6
 13 67 27 05 05 A1 C2 9C D7 B3 11 DA 43 80 B1 EC
 47 BE 06 BA 33 6B 8B EC C7 1D E6 97 48 59 D2 7B
 F1 1E 4E 2E AA 2A B9 C2 8E C8 AD 77 27 B8 35 E4
 CC AD A2 0D 89 E8 A3 84 91 E8 4E 43 A2 93 B0 CC
 CE 24 C8 B6 C1 71 0F B1 F3 EA EC 03 F3 73 DA 66
 50 DE BC 54 A2 73 07 F3 04 97 7C 45 1A 23 A6 33
 74 BB BE 9D 9C 61 67 42 71 30 47 25 70 1A 6E 1B
 DF 6B C6 07 74 B5 BA 12 E2 9F 89 FA 1E 5A B1 45
 51 C1 93 2B 6E BD 2D 70 39 04 AC FF 6B 00 C9 57
 52 DD 75 A8 C0 F3 EB F1 03 0E 1E 90 C8 2F A1 06
 01 35 BA DE A0 14 4F AC C5 DD CE 85 8A 9C DC C3
 76 FD E0 F0 BB 27 E3 9B B8 6F 00 44 6F 0A 5F 62
 3D D3 0C 92 C6 E8 74 5D 01 AD 2F A9 11 16 37 F0
 60 09 54 5F C8 E8 AB AF 57 D2 9C E6 CF 31 B8 5F
 38 3A E1 A4 09 D2 13 62 72 11 05 D9 CE 2C CF AD
 79 13 50 A4 A1 4E 7C D2 53 61 44 C0 13 36 EB FC
 8D BF BD 81 2A AA BA 86 D5 FF 12 7A 0F AE 87 F0
 49 F6 25 14 95 C5 F2 9B 37 51 FD 1E DE D8 3E 6A
 47 D1 A5 46 70 BF 6A D1 32 8B 90 17 9D 33 FD 34
 D9 99 F7 C2 03 43 D7 D3 2A 72 ED D9 CE C9 D4 57
 56 C8 C2 9B 64 D1 5F 40 6F 78 6C 24 94 2F 83 0F
 17 9D 2D EE 3B C9 BB E6 CD 17 5E A4 47 65 05 75
 E6 FD 8D 6D 3E 96 C9 ED CA 73 19 14 C1 83 EE 37
 E3 13 10 17 59 DF 79 14 F2 D5 07 98 EB 10 33 CA
 26 1D 38 EE 07 B7 43 01 D7 4A DE 69 40 27 B6 FB
 60 1B 18 AB 63 35 BB CC 55 11 F8 4A 9C F9 A5 6C
 60 DF A1 8C C4 FD 89 7B 90 E3 08 14 B5 70 DC 52
 A3 33 B1 F1 76 4A A2 09 7C B5 A1 40 69 68 0E 07
 95 AC 51 11 04 9D 0A 14 AC 70 B5 24 AF C2 1B 5B
 78 9A 92 99 E7 AF CB B4 FA 21 5D 0E 8F FA 25 52
 D9 C6 F3 AC 11 04 62 BB ED 98 00 63 55 70 68 65
 6A 7A 59 DE 09 A8 45 E3 F7 3A F0 BB 0E E3 71 6E
 99 05 CC C0 38 9C 19 A7 81 FA 42 A9 31 B5 16 F0
 89 E6 1D 32 5E 02 B0 C1 80 C1 2E C0 19 CB 90 50
 35 C4 18 EF A1 1E B4 4F D7 5B 3C 39 10 7E E5 2F
 0F 1B B4 E3 4F 17 5D 65 CC 1D 6E 69 14 F6 14 50
 C8 C1 49 CD 63 0D 6C 14 CD 41 E5 3E 1F CB DB A4
 EB 30 38 96 B4 25 86 9B 87 A5 15 33 4D 56 1D B1
 8D D7 1F 4E 97 5D D8 8F 11 1D 3D 1D EF 5F 86 14
 F0 56 99 6E B2 D2 F9 45 E1 35 64 54 6F 4E 8B 27
 7A 0B 91 AB D6 8A 22 61 36 BD 3D 6E 0E 98 A7 21
 5E 3B D1 E1 ED 90 B1 44 74 00 50 4F 7A 00 36 09
 BA 36 27 D4 C4 A4 D1 49 93 C1 DD 3D 62 DB 6F 81
 5C 08 8E E7 35 7A 8E 93 5D 44 7F 56 C6 DA BA A2
 09 0C 5F EF 90 A9 1B 76 C6 B4 F0 AE 4A C6 42 5D
 97 77 72 1D A9 69 12 C9 37 D5 AB 18 9C FE BC 4C
 23 DD FB 8C B6 ED CB C4 C0 48 4D 92 81 D8 3E 29
 38 20 8A E0 D5 FC C7 B7 D3 88 B6 51 32 54 2F 28
 A1 0F 31 22 57 0A 90 7F 31 1B 03 30 B7 5F F8 1C
 07 4F 81 BA 2B 9F 24 40 44 94 AD B1 7E D7 7F 91
 D2 75 F8 9C 53 A2 15 0F 9A E3 12 FE AE C9 FE B6
 E0 AD 51 FE AF C1 24 6A 25 5B 2D 00 85 C3 61 6F
 E9 03 49 B9 28 80 A1 93 34 DC A1 83 00 FA 48 0D
 8D EC 2C 34 69 F4 8E 36 42 62 ED 7A 7D 0C F2 DE
 9D D2 C6 92 31 BA 89 8D C0 E8 AF 43 19 83 2C 3B
 53 83 1B 20 83 AD DB 77 1D 78 11 ED 21 0B 04 54
 FE 2E 6B C8 80 58 C2 C5 0C C1 F6 E8 62 C5 0B CA
 9C A0 9B 6F 4C 08 08 53 1E B3 A5 A4 59 6A E1 6C
 0E AF 2B A5 93 75 2F 39 58 B1 56 0A DB 2A 92 DD
 49 62 7D BF 38 D1 84 CF 9B 76 BA 04 5B 63 C6 1F
 C6 4B D7 2C 0C 62 0F 37 7B 8F B9 C8 33 EB AC 32
 0D 5D 52 F5 0F E4 CD 80 5E 9E 3B A7 6D 0F 67 A6
 16 06 6A 5D C5 3F 1F 8E 79 00 38 E7 9D 42 FA 06
 E0 76 66 B8 C3 37 2E 4C 05 D3 C0 C2 A1 4B 1A 80
 3E 6A CB 07 EF C9 ED A2 CC 23 12 54 C9 52 4A 1E
 15 FA B4 03 2C 7B B9 B9 8B 33 9D 9F 40 B9 33 77
 45 34 E9 74 0D AB 39 E7 1A AD 73 C6 C2 FE 27 A6
 94 22 02 D4 9C 2B FC 83 61 A0 4C 91 56 7E 3F 9C
 1E 71 A5 17 BA 08 87 86 EE AB 24 ED FB 0E CC D2
 14 C1 F4 61 A1 3F C7 D9 9F A2 82 EE 81 C1 56 61
 1A 61 C6 47 01 0B 8C A8 5C 60 F8 D7 F6 3A B3 CB
 C8 31 D8 BC 7F 1F 1B CB CE 10 F4 BC AB 94 59 EF
 CC 2A 21 43 8E A1 5E 71 E1 81 F7 5A D4 77 7E 28
 5E 7F EE E9 6F 48 46 9E 2B 37 18 96 13 6E B2 C2
 61 E5 5D 04 28 AB DF F2 47 70 B2 A2 C9 5F 89 61
 B0 73 3A 45 37 8A 06 F1 F1 9F DC C9 20 62 9E 41
 CB E2 AD 84 C6 4A 36 D9 66 98 91 F2 B4 4E E6 FE
 53 4D ED 46 99 5B 5A 86 CC 77 0B 27 A2 D1 D2 80
 F1 CD 54 44 C0 C1 0E A3 61 16 C7 46 66 C5 76 90
 30 79 E9 14 5D EA 2F 1D E1 22 41 C9 EC A1 D3 72
 FA 33 B4 E6 31 D0 F9 89 E2 A0 02 1C C4 13 ED BA
 20 5A C3 00 E1 07 B2 E0 E0 71 76 72 3E 50 0B 80
 42 6E 8E A9 38 C7 A1 96 B8 F7 A4 E1 2D B1 E6 37
 2A 0A ED 25 7D A8 A4 15 F1 9D FC EF 89 81 7E 9C
 BB 85 82 A8 F2 B5 27 82 F7 7C 85 1C E1 4B 94 57
 4F 73 53 86 D5 98 F6 F6 19 41 74 A6 1F 4A 47 2A
 88 DF 31 1B A3 19 2C 74 FA E7 63 72 56 73 09 A7
 5A A6 04 64 96 B7 B8 58 53 27 71 BC C6 A0 B2 9B
 D1 28 A1 7B 29 35 AA 3C 60 16 15 44 B2 7A C5 B6
 52 4D CE C6 6C F5 7B 75 C2 97 E9 BE 7A 69 2B F1
 3B FF C4 3D 9E 63 F9 84 1F 04 42 7F 8A 97 60 16
 5D 53 CB A9 88 61 C3 37 16 41 49 70 24 C3 EE A0
 1B 4B 00 0D 52 18 8D E2 20 F7 D4 44 0C E4 25 E1
 82 64 6F 01 5B D3 F8 F2 F3 84 57 F9 7C 5B C5 21
 18 1C BC 3B BB DE FD 36 F6 D6 C0 C2 F7 12 95 53
 8B BF 89 B0 B6 84 16 39 D0 B2 0F B2 5D E1 B0 4D
 00 A0 7F 81 F2 5F 66 CC 3D 34 BA FE 72 F3 46 26
 EA F3 2A A6 F4 73 25 C0 D8 C2 88 8E BB 10 6E 44
 99 E7 62 D0 0A BC 66 A7 AD EF 9C 54 23 61 5E 37
 A4 C6 6F A5 B2 88 7B C6 48 3F A0 F9 40 D3 6D CC
 CC F7 1A BB 5F 46 5F 68 B6 19 BB 44 EC 50 44 9B
 C0 26 D2 FB 36 67 C3 9B CC 79 68 2B 0A A7 6F 3E
 36 53 2D 6C CF 49 30 C6 9A 27 91 D7 D4 EC 7C 94
 18 8C 03 3D 5A 84 4F 6C 87 18 9A 95 AF 1C D9 7F
 52 01 11 49 EB 84 48 4B 6E 12 C5 DD C0 18 66 17
 F2 DA BC 6E 5A 2C 3F 6B DB E7 72 83 4D D4 BB B6
 F2 DD 85 9F C9 0A F8 93 8E 3E 65 0F 77 30 A5 4C
 41 5C 3F 77 5E 18 D3 5B 23 22 4E 05 E7 23 A4 AB
 FB E6 80 57 59 AC 25 A6 20 35 EE 13 E0 1E 54 8C
 C6 60 F4 E8 30 6E 3D 93 2C 4B DB B3 D5 58 F8 6B
 9B 1F 82 66 0C A7 07 B6 83 38 B0 7A 08 92 29 26
 CC 17 FA 06 FE 13 23 AE A2 C3 D6 70 58 FA 2D 16
 8B D1 6D 25 5A DD 33 A6 66 49 69 BB D5 B7 AE 98
 47 6E 95 11 BB 00 BB 70 CD A8 EA 01 AA 56 6F 28
 18 22 75 D6 0C E6 27 E7 8A 21 D0 8C 54 48 C7 08
 78 DC 3D 33 45 79 73 2C 5C 61 97 B3 9D 90 FB F9
 C6 30 8A 56 3F 5B 73 7E F2 49 6D E7 28 2D A3 08
 10 F0 A5 FD 62 F5 AA 5B 42 14 50 42 20 EE 01 5C
 53 88 A1 A5 93 F5 D8 DA FC 4F 6B 91 49 2F C3 25
 61 C9 95 76 BC 37 25 7A F2 C5 99 3F 52 C9 A1 3D
 48 19 52 FB 65 7C BB 42 88 33 4A 66 11 39 DA 5B
 CE 24 D1 96 43 C5 C1 AD B9 7D 90 E7 D6 47 F7 56
 56 A8 15 52 05 01 7E 26 34 C7 E7 C4 C4 FD 50 6F
 FD AA FE 20 B7 C2 54 1A C1 B9 95 76 88 1D A3 97
 8B E2 17 93 60 A8 0E C0 C0 68 24 61 16 1B 32 8A
 8C E8 59 34 83 89 CC BD 58 95 B7 CB 50 69 46 BD
 FF 79 C4 D3 59 65 2C F5 F3 E5 8D 92 57 C6 96 25
 32 28 56 81 40 F2 F1 F5 64 41 89 90 13 88 A9 CE
 39 A9 47 B5 18 C8 AA E1 79 81 5F 23 21 3B 1B FF
 5F 52 B6 4B 4F 2B E3 7F D6 69 3A 4C F2 B3 51 6A
 B5 F7 7B 13 F2 F4 FF 98 EE A7 07 EA 8B B7 94 B0
 A0 D1 4F 65 DC 99 87 01 61 84 33 C9 A1 1B 87 4F
 C3 11 D0 F7 61 74 9D B2 FF 69 72 92 37 FD 5B DB
 6F B3 D5 1C 21 5C 83 89 09 DF 98 4E 75 25 A4 EB
 1C 30 43 1E 81 F9 31 09 FC 3F 26 54 D2 52 CF A4
 53 FB 6C 52 E7 70 8F 85 B5 20 4B 95 E5 2A FB 3B
 C4 76 A6 31 BC AC 40 1B 34 89 23 8C 86 04 E8 E1
 1D D5 EE 2D 62 FA 06 16 C6 37 13 01 18 F0 BE 21
 7C 88 A7 FB 5C F6 55 25 92 04 0E FD 4B 3D DB B5
 BB 5F 91 D7 5E 18 D7 7E EE 7A 9D 47 BA 46 48 B8
 5A 98 F2 BF 26 72 C7 1A B1 18 92 D6 3C F0 E1 99
 25 7E A6 AB 2F 40 59 48 B3 EC 53 28 AE C7 36 C7
 0E D8 2C 0C F8 B4 63 CD 72 80 33 00 81 BE 0A DA
 36 7E 37 AB DA 94 38 FC 23 7B EA 46 5E A1 B4 BF
 E9 B8 D0 C7 4B 08 7E 7C 2A FB 88 4A 5A 35 36 A3
 AB 00 D8 AC 9D 47 A9 7F CF 97 76 31 BB 47 FF D1
 C1 62 48 2D 88 2F 28 AC 88 21 0F 4A 23 05 D7 20
 D4 08 84 05 24 17 29 20 DD AC 0D CF 9B F8 20 D6
 9C 2E FF 47 CA CD BD C8 DD CD 65 24 39 6E 87 B2
 AE C1 F9 5B D5 CF 83 93 2D AC 30 24 E2 B9 74 6F
 4A E9 D5 D7 15 60 20 2E A9 14 9E 66 34 C3 FD 46
 F1 C3 24 5E 54 1E 12 43 9E 27 89 93 BE 8F 0C 12
 77 47 71 AC 90 2E D1 40 9C C3 91 E6 13 C0 E6 53
 AF A9 B5 92 61 39 74 83 27 96 D9 AB E1 BD 8F F3
 BC C4 B8 99 44 9D 1F AB 0C 99 75 63 12 A8 31 00
 68 F5 9A 61 AC 04 6D FE A3 CF 90 23 23 AD BF 88
 8F 8E F7 65 42 27 D8 25 4A 30 81 76 BF 16 B5 A9
 60 AE A4 19 93 24 F1 E0 2F FF 6E A7 D6 1D 15 79
 75 43 F6 87 34 B0 5F 43 B4 F7 57 86 45 8F 9A F1
 DE 88 4B 27 BF 00 D4 07 BE F9 8B B9 86 F2 3E A5
 07 DA 9D C6 98 70 E2 A5 9B 2B 3A E0 E8 E8 60 EA
 AC C3 78 5E 80 5D 62 77 E8 D8 D2 C9 77 A1 98 49
 CC A2 BD 30 77 25 B0 4F C6 3B 4E 01 3C 99 89 E4
 83 84 D1 2A 53 60 50 1C 46 2C 67 6F 41 CA BA C7
 E1 56 30 F1 E3 7E 11 77 B5 96 15 69 DD 21 28 68
 B0 6B 53 59 EA 09 6E EB 6D 76 0B 5B B6 17 3D C5
 56 66 9C A9 43 9C 17 91 F2 97 B3 FE 58 4D 46 DB
 23 BE B3 66 A9 6C 3B AA A0 A8 0D 1B D9 37 96 00
 1A 8D 59 A6 1C F2 37 37 11 10 62 7E 24 2B B1 ED
 D2 E8 1C 14 45 52 19 B5 11 32 93 4E 3E 5C 9B 27
 18 70 CA 22 6C 15 20 91 4D 34 FA 04 85 CC 0D 7C
 FE AE 9C A4 0B A6 6C DF 1E EE 49 8A C9 E2 A6 86
 27 6D 09 1C 3D 31 17 64 F5 61 3E 4C C7 75 5B 26
 0A 36 6B DF E9 87 5B F0 C2 D8 C9 79 55 CF 9B F0
 CB 15 C0 E4 1E 04 CA 64 2F 4E D3 CD 7B 43 36 79
 AE 34 3E 42 C2 4F 84 3F 8C E5 CB 53 8D 48 FC 1C
 88 D6 C2 20 52 50 BD E5 AF 82 80 1F 97 4F 3A A0
 FA 3F 5C 38 8B 1D 3B 14 57 37 A3 F9 2A D5 EB 50
 81 91 1B 4A DA 77 2F F8 80 0C 27 A2 03 0B 6C CA
 4F 2E E2 4F D9 CD 34 90 79 25 FE 4B 3B 37 FB 78
 5B FA FE DB 43 60 02 9A 03 F3 65 A8 90 02 68 4C
 48 48 BE E3 13 F4 42 C2 D6 A8 F2 97 A4 EA 74 DC
 42 D4 51 88 E1 97 77 B6 F6 5F 1E 8B F0 03 00 85
 A8 47 00 E7 90 8E DC 1D 0A B0 85 9D 9E F9 62 2B
 9D B8 19 2E D2 22 0D 4A 5D 23 8D F1 3A 83 0D 0A
 1A A5 C0 E2 B7 1C E7 14 6F 4A 0F 69 57 94 57 91
 A4 AF DC 3E 89 EB 94 E7 2D 62 23 8A 67 EA 3C C5
 86 2D EA 09 0B FE FD 9D 54 B5 E8 B3 26 EA 46 34
 39 38 26 B9 FE F5 6D 07 9F 7E 59 BE FC 1A 5F 12
 62 97 F2 9D C5 22 18 72 DB C5 E6 FB 9C 26 3C F3
 D6 74 77 68 08 34 C9 8D 41 E4 1F 36 D3 3A 5B 73
 FB 53 B6 60 ED 76 F4 EB 48 90 7F 2E DE 8A 2D 50
 80 6A 49 6B A7 B2 58 00 51 09 F1 2A 18 32 47 53
 A5 50 9D 0C 83 E3 B3 AA FD A3 DD 25 1F CF 1B 05
 04 7E 60 79 48 99 43 C9 CC 6F 49 67 69 E3 D7 F8
 11 8F EA 50 A3 D2 4A 3F 01 7D 4C 1C 2C EA CE 16
 CB F9 E3 F3 59 79 E8 24 56 77 D3 C0 C5 10 65 45
 B9 96 5E 34 55 A9 5C A8 8E 03 FE 47 27 5F E3 3B
 12 C1 EC 38 FF 55 39 29 D1 D6 DB 76 78 39 FB 1D
 63 45 2B 09 18 38 71 A5 BB 86 94 54 6D 5F AF 8B
 BC 8C 93 05 F6 52 82 E9 C4 68 0C 91 38 C9 F9 A3
 B9 14 4F D9 88 B9 25 7A AC 8E 08 33 F9 9D E9 47
 D9 61 F6 C2 58 4F 97 88 C3 B7 1F C4 7B AE 92 62
 16 E6 82 F3 4B 99 4B 02 52 45 97 21 F0 0C D0 66
 0D BC B7 0A 88 36 10 F9 EE 48 E2 E5 C5 DD B9 0F
 6A EA 0C 48 B1 68 C6 89 A7 E3 E0 09 F7 B4 2E EC
 7A F4 A6 A1 F3 F2 AB AF 65 59 47 29 8B B0 0F 19
 70 15 0F E7 18 C0 A7 DC 5A A2 C3 72 83 A3 8B C7
 40 67 98 42 FD D4 DB B2 07 A6 CC C9 23 67 1C A9
 A0 49 5E 20 C9 EE B1 24 8C 71 28 13 9D 88 25 F5
 73 EB 49 FF 67 CE FE 01 E0 D3 28 00 FE 16 C4 C8
 C8 EA 5C 99 B9 BD D1 B0 0B AE C4 B2 67 2C 51 95
 69 86 C6 19 52 48 93 81 AD E6 1E F5 48 AE 76 58
 69 DB 3B 24 84 19 8D E9 A1 5C 3D 18 2C F4 0D 1C
 D8 4C 5E 34 F1 7B 58 0E 4E 8F F6 65 E1 07 B7 E2
 50 FE 65 09 38 73 51 10 48 62 A9 C6 5E 3C 4E CB
 55 D1 7A 35 BD 4B 25 58 7B 08 3E 41 D1 EB 8A 69
 45 5D E6 29 A9 07 45 31 FA 2A 42 DD E1 9F D9 F9
 2C 25 17 9D 06 3C 39 8C C6 71 2A 5A 24 11 D8 3C
 0A 76 3B 90 14 44 4C 19 7A 28 A3 B9 E7 51 B4 A5
 15 43 EC 73 68 46 39 45 E7 CF B6 2D CD D0 7A 5F
 4A 91 AB 21 2D A3 D0 34 83 71 42 6C 0A CE E4 4E
 FF 5A F9 92 F7 46 2F C9 D0 91 59 11 BF BF B9 43
 E7 FA 56 1A 05 51 B9 DC 2F 8E DE FA D7 B0 A9 8F
 19 EA 34 C0 A3 86 32 C6 CC 9C 22 9B 41 73 41 82
 F9 BA 5E F9 3D 4C 1D 2E 86 85 58 5E 5F 15 4C E7
 5B B6 A5 81 0C 49 FF 05 86 2B D0 41 83 5E 03 F8
 C2 32 56 FB 97 9D 13 4D A1 15 F7 D7 7E 90 89 D5
 18 18 00 33 8B B0 25 1E E0 59 18 E9 C7 B2 F7 06
 5B D0 7D 36 4D DC 13 1A 90 63 83 7E A4 6F 0A 51
 86 0A 83 C4 9C D4 8A 9D 85 E4 7B 8B 8F 13 95 B6
 6D C8 16 96 59 A4 91 97 70 DE 35 FC F6 04 D4 05
 FD B9 BC BD C5 2E 0C 29 73 B0 0D 6A 83 91 C5 DF
 ED 7A C2 56 F3 DB F2 49 C4 FD 6F 85 02 E7 FF A5
 EE 1C 78 59 52 53 E8 48 09 73 A3 CC AC 58 02 03
 AA 15 DC A9 84 BE C8 7E 68 39 99 6A 12 FD B6 60
 CC 23 43 FD AC 23 92 59 4D C4 4F 11 9F D3 F8 7C
 EA 1A FA BB 65 50 4C E9 F1 AA 51 57 D1 3B CD 9C
 5C 8B 69 96 1E A6 BD CE 47 E8 AC 82 3A D9 81 B9
 E3 CF 51 A3 98 56 89 93 8E B3 13 60 A7 EC C9 C0
 70 4F 7D F6 C4 D5 4F 44 80 75 0D 31 78 91 DB 90
 22 A8 42 CB C9 E7 8C A6 6C C3 C2 6C 58 D9 37 7F
 26 C9 41 54 DF 7F 9A 2A EF B9 DE 43 B8 38 31 BB
 E9 61 ED DD 13 77 C2 57 1C 60 4E BC CC 2F B0 17
 63 6B 11 45 43 FA 32 07 14 C3 C0 66 DB 62 8F 2B
 63 9A 7B E7 B5 0E 35 CA 86 55 6C FB 0D 83 C3 2B
 B8 F0 38 89 1B 9A 96 5A E4 AB E8 3A 32 4E F9 7E
 3F 54 0B 6E BA EF 0B 72 A3 41 EF E8 06 03 AF CB
 B7 90 03 06 7C D0 78 C7 1C 43 07 26 68 4F 70 DA
 87 3D 3A F1 21 AD 3C F1 53 69 79 07 3E F8 2C 00
 F1 C7 86 40 B7 00 99 4A B3 10 BD A5 0E F4 21 B3
 F7 01 8C 2B 4E 41 66 82 11 5F 98 9A D9 D1 CB 8E
 90 1C 90 34 89 24 A3 05 2C 47 E4 57 3C FF 14 9D
 35 7C E9 20 98 62 27 A1 F5 B6 3B 30 6B 26 6B 91
 4E 32 C5 8F 2A AA 80 81 B8 47 04 81 E9 1C CB A9
 FC DA 16 40 C6 E1 CA B0 11 81 B4 D5 5A 02 E5 32
 56 E8 AC AD 6E 76 17 C5 61 33 EB 7F 7A C7 50 C8
 43 A3 88 FB 37 80 2C 7B E6 4B 08 91 29 D0 65 96
 89 1D 60 AC B3 42 C9 56 A6 B1 F7 53 AB FD 3D FE
 6F 87 D5 6A 39 8A 97 24 6A BC 18 1F A4 B7 97 97
 0B 4D F1 43 63 9B 78 1B 14 D5 F0 07 7D BF 3F 02
 29 8C 27 AC 6E 2E 7A 53 7B 02 4E 70 FC 86 AF 0E
 A1 1B 07 B3 D7 B2 3C 60 0A F8 79 FE 4E E4 0E BD
 B7 2C 2C AD DD 38 96 2B 57 92 AF 09 79 12 AE 91
 E3 B4 72 34 74 4A CD A7 C5 A0 EA D1 99 42 28 87
 5B 81 D7 F2 54 71 EC E0 77 42 35 DE A7 FC E7 E4
 94 CA 76 79 A1 7E 45 CF 85 C4 2A A2 C3 D7 4A C8
 E3 C7 18 E0 56 48 EA DD 73 7B 9D 6A 05 00 5B FF
 3E 71 65 DA E5 36 D6 41 36 3E CD 08 16 50 C2 13
 AF 93 AB 7D 29 71 61 67 F9 4C A1 48 4D C8 E9 CD
 F3 B5 69 14 FD DA 12 2F 76 8B 6E 39 74 44 C1 76
 46 55 11 7D 3A 08 D7 53 82 92 88 03 DC 8B 2A 87
 AE 42 8B 8C 63 F9 DD 31 17 51 73 1A 6D FD F5 00
 77 02 7F 89 2C E3 FD E7 AD 83 E6 54 0B 3A 87 25
 27 6B 84 42 FC E6 8B 79 95 45 BC 20 F4 F7 9F FD
 DF 34 B4 18 23 81 99 6F F9 AA 23 5D 46 12 39 85
 96 2C 25 C7 EB A5 91 5A FB EA 86 37 63 EB CE A3
 4A F5 4A DA B9 49 96 4E 23 88 BF 23 E2 49 7C CC
 CA D0 19 EA 97 9A B8 9E FE 50 E1 BF DB 46 86 BB
 DC C3 BD 2A 60 1A 5B B7 83 78 45 B8 8B 61 9E 92
 3A 8E D1 B9 70 E5 2E B7 78 82 DC AF DF 3E A3 0C
 78 CC 7D 19 56 79 52 56 13 E4 06 21 93 29 B3 AF
 21 3F CE D3 46 9D 09 75 D4 5A 92 EC B9 1D 6B 6A
 F6 82 D6 55 17 56 CD 6E EB AE 2E B6 9C C4 18 2F
 01 BA 01 72 2F 10 96 DC 09 7B 96 30 FB BD E6 0B
 16 D9 3F 62 28 BA 31 FD 2C C5 8C 40 B2 5F 2D 95
 7F 49 AA 5B EF C4 EC FE 4C 6D 36 A0 11 4C C6 14
 6A E7 0C D8 EA 1E 41 88 58 FB 20 AE 02 DA AE B7
 79 E4 1C 79 65 47 24 FE 8A 05 A1 05 17 1F 3B 7E
 D8 EA 5C 4A 8D E0 F6 13 F4 5A 9D 79 3A EA F2 F2
 BB B0 76 29 B4 3B EA 07 A1 02 CA 97 8F E2 CF DB
 F6 71 00 58 8C 8F EB B1 54 14 CF 13 1B D4 80 74
 0B 1A AD C9 60 D5 56 0A 0A 2B A7 94 BB 5F 11 1D
 51 5A D0 1B BB D0 15 17 0B B4 A2 DC 69 C8 FC 89
 9D 1B 1B 0C BC 51 5B C6 65 8A A1 D3 79 EE E0 94
 AE 37 43 F7 93 44 6C 68 97 A6 31 57 2D 80 8A F0
 CF 99 14 CB 9E FD 49 5E 24 73 E1 37 42 FC AC 76
 80 76 08 8F AE E8 04 9F D7 83 35 19 07 A9 1D B3
 B9 FE 88 0D AC 6B F1 63 CA 8B 5D BD FA 4F 98 E7
 6B 17 3E 11 CB 81 C3 3D E6 43 F0 B8 8E 2B 94 2C
 4D 6F 63 6A 87 E6 71 E4 71 C6 42 90 4D B9 45 79
 A1 37 86 EB 6A A0 3F AC C8 05 A6 B5 CF AC C9 09
 70 94 22 C5 10 A7 9D C3 26 E2 AF 39 F0 4B 79 D8
 CE 76 84 CB 21 7E 81 1E 04 A9 3A FE 8D 36 1D E1
 57 49 1B 1E 56 EA 1E 88 8D CC 32 75 04 F5 5D 13
 D1 36 69 5B E6 CE 3A DF E0 FF ED A2 B6 E5 43 ED
 E1 09 58 F5 88 EB FE 7C 3E 0C BD A5 A7 72 CB 13
 E1 18 71 C8 DE 35 2D FA 13 0E B5 7E 02 CB 68 47
 98 04 36 F2 79 7F 9A 28 84 BE CF 7C 0B 51 12 45
 14 D3 27 5F 00 02 20 E9 9F FD 17 B0 82 12 B5 7C
 96 3D 38 CE AB 5E E2 25 FB B2 40 A7 4F 45 9A FC
 71 AC 5C 8A 51 43 0B C6 E9 32 30 A9 15 20 60 74
 A7 8E 64 6A C0 8B F2 8A 1E 70 D9 D3 83 70 26 84
 8B 73 68 C8 A7 D4 44 B9 AF 1D 7E C7 9E ED D0 9B
 52 66 AE 2A E2 91 32 C1 A0 16 BE 3D A7 F4 60 F3
 67 10 5C 44 55 DF E2 79 E2 DB 71 F4 87 21 3A C8
 95 19 E4 B6 09 4D 6E 85 1D E6 5B AA EB C4 F5 48
 0D F0 9D B5 9E 5E 1B 41 F1 C1 C0 54 C4 17 0B 52
 29 E2 DB 44 EF 6B 0C 9F 69 32 97 24 40 2A 0C 51
 00 21 87 51 63 48 5E E1 6A 49 27 97 46 DA 3B 96
 96 9A 93 8A D6 D5 81 8D EF 73 D4 58 8D B6 65 FC
 67 1B D1 20 23 06 6B BB 06 5C 92 2F 9E 52 6A F7
 3B F4 0F 36 66 1A 9D 3B 72 BB E2 EF AA DE 5D 18
 85 4A 76 B0 6F 79 53 54 6A EE 0B 59 F1 98 AC 17
 0E FC CB AF 18 A7 65 8A 98 A3 F8 D6 95 6B 08 F6
 FD F6 C9 8D 98 E1 A0 46 26 5B A6 5E 3A 0D EB 35
 2C 1A 43 E2 C8 59 D1 0A 2D 62 C2 39 9C AB DC C4
 16 79 D4 8B 2A 7D 9E 6F D7 E8 A0 2F D9 A2 CB 9E
 53 EC 8C F3 F5 27 D8 F1 07 01 80 70 35 0F 75 C3
 CB CA 2D 64 12 51 4D E9 0B C0 88 D8 96 0B E7 5B
 10 A3 7B D9 AB F8 C1 54 56 88 64 DD 6F 28 58 5B
 73 58 BC B0 1D 1B 41 65 E7 B0 3B 22 FB 51 AF 38
 91 F5 09 DA FC 3A 81 1F 01 E5 B7 D9 DB 3F 18 95
 FA AB 9E 7F 8D 97 D7 DD 1E C4 17 2B 37 4F 9F EC
 6F AD C6 B4 AB 14 72 82 BC CA 28 52 11 61 4F C1
 03 3D 0D 18 9B 01 90 22 68 25 9B BB 1C 72 6F 6E
 FE C3 7E AB 2F 91 CD A0 89 C9 55 2B 47 A7 B4 18
 67 67 34 20 16 6D 8F 4C BD 63 00 7D F6 79 70 84
 80 D9 29 E8 70 5E FF 0D 7A AD 1D 43 DC D7 30 C2
 E5 0F 6C AD EB 6E 6C A1 58 B4 7B E8 27 08 1E 5C
 A6 8B 52 EB 74 C8 BB BA BF 66 1D F5 01 A4 7D 49
 77 F9 E3 CC 49 FC 61 25 25 0E BE E6 F8 68 4B C9
 F4 D8 DC AA 89 CE 09 D2 70 D8 F4 19 42 39 22 42
 B7 29 CA 3A 7A 80 87 2F 67 74 90 52 B3 9B 50 B8
 29 49 9F 12 48 BC EF F8 AB FC 0A 3F AA EB C1 22
 1E A8 6F F3 E8 61 3F 94 A5 1B F5 2A CC 5E E9 59
 F2 B0 3F F2 2D AF 52 64 15 1F DD 83 92 F3 F4 08
 E8 12 12 69 A1 06 CD 15 48 90 3C CF A3 40 7F 5B
 77 52 0F 48 85 C1 FE B7 58 AD 72 F4 A4 D8 BB 98
 7F DB 33 14 86 87 33 4F BC CC B2 61 26 EB 55 A1
 E8 D0 89 68 0F F9 65 21 59 99 83 AA E6 E3 A8 64
 9B 6A CC 4D 96 5C C7 66 B2 8B DF 20 9A CE 74 AF
 5B 46 86 67 B9 30 F1 EA 30 5E 65 FB 7C F2 36 36
 5A 56 2B 6D A9 F9 CE 6F E8 37 98 66 CC DC DA 36
 19 81 55 8F C4 AE FA 76 34 E9 13 98 98 74 C8 FE
 87 BA 20 F2 C4 EC 42 F9 DC 6D FE 40 A1 A7 C0 46
 15 3A DA E3 A9 08 5B DA 5B 92 02 B5 7B D6 B4 C4
 4B 06 57 57 D8 85 D7 0B 0C 79 76 9D 41 D4 58 D0
 EA 7B 98 CA 35 E9 51 BB 72 B2 3B 0F 14 2D 3B 80
 F5 8F 43 44 B0 4D 8E 0A 30 C3 14 D1 B6 7B C5 04
 8D 31 21 65 F0 F2 DC 60 53 DE E6 81 11 87 B3 70
 17 F5 E5 FA 1B 9E 59 D4 7B 1C 03 35 66 A6 47 9F
 56 98 BB 7D 71 8B 1A 39 F9 B3 72 0D 24 13 5B 94
 85 84 1E ED D8 66 D1 D7 E4 7A B2 7B 0F AB 4D 20
 25 D8 A6 73 07 B0 CE 07 19 DF 38 C4 E3 04 4C 8C
 F6 A5 DD 65 94 24 C0 D3 98 DF 4B 09 AD A5 EC 68
 8D 6E 8B 35 7A 3E 49 55 2B 1B 3C 39 93 14 A0 39
 7E 45 4C 5A 8E BC 68 DA 82 FB 85 97 4B 85 D8 72
 BE A8 21 E2 E3 0F 26 10 94 41 F1 13 B7 A2 A5 9D
 99 88 25 48 7D CB F8 7D BC A8 C1 25 BB C2 80 BA
 E7 12 DA DA F9 F4 7D 50 0A 12 4C 27 B9 17 A9 88
 DA 27 BA 42 AC 86 C9 5C 08 0F 7A 63 2F 0E C1 5B
 95 4F D6 E5 C2 B8 38 C9 90 2D A7 5C B9 E6 FC 5B
 47 FD 51 8C 68 EA 32 43 6C 19 B2 57 FC 2B DC 40
 86 FE EA 6A 3F 9A CA 94 97 0C 34 04 6F E4 11 0C
 52 17 7B DF 2F A5 50 F6 6E 4D 36 21 B8 06 5D 11
 E3 35 D0 DC B6 8D EC CA 2A AD F8 A7 72 B3 74 74
 34 5A 5E F3 59 F6 16 EC CF 8C 42 BA EF 68 F2 2C
 F1 A4 A8 B1 1A 2B BF AA B2 6D BA 09 47 ED F6 52
 6D BD 2A 34 FC 31 27 E7 9D 98 98 49 04 15 79 D0
 39 B5 55 E2 5C EE 13 61 04 10 02 27 5B 58 00 CB
 E5 78 03 EB C1 14 B6 C0 3D FA 2F DF 2B E9 42 18
 A3 13 22 F5 55 B2 D4 7B DC B5 4D 8B F5 2E 43 7D
 F4 6D BE 6B E5 92 AF C0 16 9B 6E BA 99 35 47 0E
 AB F0 D0 DF D8 ED 5D 0C F9 7D 8B 56 05 30 99 64
 F8 2B 6B 48 DB FF 72 99 67 E2 79 25 70 41 E6 D1
 4D 9F 20 C2 4B 56 A8 BB B1 23 F5 97 07 C9 10 81
 BB 37 A8 5D 9C 50 5C 70 CD 36 53 EA 5E 9B 3E 6C
 30 DF 6E A9 CB F0 EF 63 BE BC DA 1F 00 92 57 96
 20 C0 17 91 7E 9F 05 C3 2F 9C C0 99 FF B6 24 B1
 E8 20 AE 07 57 F9 CF 73 F8 9D F2 08 1A A2 06 5D
 C6 4A E9 A8 54 0F 39 E1 8A 8E 97 1F 39 31 BA 3D
 4A 9B 9D AA 45 B7 13 57 53 D1 42 2D 11 2E 49 8D
 4B 50 AB BA 41 62 34 50 C7 BC 44 E5 11 3B 90 FD
 3B 72 D1 42 84 15 1A B8 22 2C E9 A9 C2 51 C8 EF
 6F 0D 2C 97 AE 46 23 69 D4 AC 60 FB DE B7 8F 89
 92 4A 98 CD 61 F8 11 A9 5F 6E 84 0E 43 5A F2 12
 23 2D E1 90 B3 5F AE D5 2C C4 7D 31 1B 59 23 32
 73 D7 7D 3F 94 61 2D 13 96 61 16 AD 6B D2 FB 0C
 59 A5 FE 63 8C 4B 4F 79 6A 34 93 4D EE E1 CA AC
 2A 8C FE AD 2A 1D 26 9C 5A 7B 3F F8 4F ED 30 1C
 76 7A 3A D1 1F 45 A7 4E 4B 49 13 A7 61 0F 6F F5
 BE E6 F2 17 6F 54 97 81 3C ED 1F AE 4F 29 80 33
 EF BE 19 76 7D DD F9 52 05 4E 7D 4B 0D F3 E1 61
 92 B7 56 2E F4 C8 5A F3 D4 4D 83 98 8E A3 08 3E
 08 0F 7E 17 0B 8D 47 45 82 67 5D 27 7E 94 F1 E5
 A2 7E 35 EB 2D 05 64 AA 26 52 8F E5 C6 0D 52 7C
 63 FC 5D A5 BA E1 DA C3 68 4C 7D 13 ED 52 61 A3
 C2 76 BE EA F7 C8 5C DC 70 5B FA 90 E7 BE 20 CF
 23 5B 00 4C C1 3E 96 19 A4 5C 11 07 36 64 BF D1
 69 57 83 6B 74 BB 62 0E DC 9B 9B 88 F8 70 34 31
 46 11 2D 51 9D D8 56 B0 EF B6 29 42 FD CC E1 6C
 88 69 40 4D 73 36 8F 27 84 22 13 8E B5 0A 7F 99
 F2 A6 A4 17 D2 FB 78 BA 60 8F F5 BC BA 95 DA 81
 CA 18 C7 C7 B8 76 AA 70 3C EA 24 A0 D2 97 DC 86
 1F 8A 3E D6 32 80 62 CE 6F FA CE F2 05 01 D8 AE
 E3 1D 3A 1D 25 7F 69 03 6B 0B 59 BD 8C F8 02 A3
 5C 3E EF 06 29 1D AC E5 33 F2 15 47 F2 C9 8B 6B
 6A 2E 77 F0 48 A8 F1 BA 40 B3 8D 6E 54 E1 98 05
 49 9F 60 29 6E B1 02 1C AA AB 01 8E CA A8 8B A2
 98 2A 76 CD 3C 08 BD CC 45 01 5F 12 FE 8C B6 5F
 4A F5 15 FA 4D 9C 22 FE 82 78 12 2C 25 FC 95 36
 70 15 BD 5D EF 7B 4C 7F 69 50 2A 27 BA 0D 37 C6
 1F 15 7D 87 15 39 13 CE 46 46 2D 30 3C 5C 5E 20
 1D E1 27 F7 94 28 2C 4A DE 21 F3 4E AC CE 5E FC
 12 04 54 53 BC 76 CE 1A 0C 6B CE 93 F6 D7 09 29
 3B 1D 35 34 35 8D 31 E9 82 5B F9 68 1F 06 18 98
 D8 0C B5 C6 CA FD EB 14 61 0D DA D4 B3 3A 9B B4
 2D 49 46 E5 37 8D 08 2A 88 21 C8 2E 81 F3 20 04
 70 E4 67 F3 31 A0 71 97 F8 EF C7 E8 52 51 17 EC
 E8 02 D7 EB 45 2F 5F 47 9B 76 BB C6 14 DE 05 D1
 5E 42 76 5D 0B 3D 8E FD 5B 8C 89 73 D9 BD 43 59
 B6 80 A3 70 F3 EB 42 B8 B8 BD EC BA 0E 1A B1 D5
 31 46 93 1C E6 71 C0 70 8F CC A4 F0 8F 92 12 C8
 0E 55 35 41 B3 CA 02 3A A5 18 6F 05 87 F8 82 9A
 B0 07 91 8A 0C 85 F7 29 A1 EA E3 AF 14 F1 2B 91
 AC F6 60 B9 1E 99 43 8D 6E FE 5C 8C 27 E3 14 EF
 30 79 BE E0 48 BA 7B CB 74 60 22 40 0B D9 32 C4
 65 AE 11 9D C4 2B 16 F0 F2 63 5C 7B 05 84 0A 04
 E2 A0 10 A8 7C 5F 21 06 86 63 2A 22 A3 D4 B2 1A
 A9 0E 22 AC 34 AD F6 F0 9E 8A F0 0B F6 79 50 09
 FC AF 3C BE BF CF 18 FD B6 B7 07 B1 0F 0A 50 B6
 6E D2 BE B9 7E 61 0B 86 21 11 BC B1 8D E7 A7 9D
 03 70 62 40 5F 35 22 DB 62 12 D7 EC DA A2 4A 30
 1E BA 15 D2 6B A5 A8 65 A4 D6 52 DF 04 73 B5 A9
 84 42 4E 41 3B 2C F0 F5 EB 3B C5 9E 9B FA BE BF
 DC DA D1 76 FC C2 56 8C 0B 06 EE 75 4D 53 A6 AB
 E0 1A 71 18 F1 3D 02 41 83 CA 29 57 C0 23 01 DF
 1C B4 C3 72 C3 E7 5C B2 8B F3 15 E4 37 06 43 A7
 13 8E 94 D1 E4 7C 24 4D 64 85 01 4D B0 FB B2 EB
 7F 12 28 E4 33 5A 6B FC 96 D3 77 67 8A A9 E5 D5
 0C 7C 5E BB AC EE 6E CB 2F 18 43 6A B2 7D FB 1C
 8E C6 75 F5 BA 2E 13 16 8C 06 D4 65 16 0E 1F 3F
 EF 54 60 38 C1 AB 5D 34 60 4F DD CB 42 6C AC E7
 33 51 8F FC 1E CC 94 E3 55 0D 54 7A C4 37 B7 7A
 0F B3 9C 9A 70 CC F8 A2 D4 4D D2 AA 97 B4 7E 76
 85 F5 D8 38 A8 50 BF B5 EE 90 EE 13 DA CD E0 F3
 B4 32 C7 68 28 4B A4 7F D8 94 E9 23 D2 52 D0 79
 21 2E 1E D9 4C 02 27 8B BD 01 8B 8D 69 FB 36 26
 41 4C F0 E6 B1 F0 BE 6D FE DC 1A 31 9D 9D 84 38
 D5 E0 38 3F E7 BD 5A E5 F5 86 B4 8E 90 09 D8 89
 29 EE F8 4A 1A 51 E4 57 69 4D DA D0 A6 35 50 82
 30 AB D8 70 8C B3 68 7B A4 06 2A 51 33 E7 E9 27
 96 82 6E 28 99 5E 94 A1 27 D4 0C EF EB DA AD 37
 C1 6E 00 1E C7 D7 1B F9 C7 FF CA 6C 0C 21 B7 92
 57 41 95 6D 95 55 46 00 AC 6F 48 1D 62 96 25 5C
 D8 3B 54 41 46 8B 1B 6B 1C 07 C5 93 3F AF B0 77
 85 A1 F9 33 9E 52 78 FC DD 5F EF 52 40 A4 6B A4
 B2 6E 97 37 46 88 FD AD 19 FA 30 A3 C8 C1 1A 2B
 69 2F E2 8E 61 7A CC 72 50 AC 83 77 8D EC F5 7E
 0D 6A 3C B6 CB 05 9B 08 F9 18 1A 69 D5 33 58 F6
 C4 4C 0E FC 10 6E C6 7C 61 36 7B 7F 11 21 E4 71
 8E BD 21 35 78 BE D6 A4 4B CE 8B 8A 69 B6 5E 23
 46 81 7D CA 5B D9 32 C6 48 49 51 42 CF 1E B9 8B
 49 8D 9D 4A 96 FF C0 02 EA 60 E8 C2 BF FA 72 CB
 8A B1 4B 9E A0 75 35 46 DE 5F 68 8E 8E B6 CC 0D
 DC ED 0F 54 99 11 D7 55 9A 1D 54 D3 B2 10 04 3A
 68 F0 DB E4 63 F1 19 81 E5 76 B1 59 22 3C 73 7F
 6A 77 37 CE 67 17 B8 36 FF BE 3A 1B 02 DA 8B 1D
 3F 86 A9 6E 56 43 9B F4 F6 41 FB 78 78 58 C6 56
 44 D8 09 F6 7A E8 68 D3 62 D4 A8 28 9D F2 78 CB
 0F D5 C0 30 B7 F8 A5 F7 61 2B B2 FD 51 5C C1 63
 F6 3F C2 84 90 23 34 31 18 05 AF BA D5 9B 19 32
 81 C8 39 79 86 62 AB 6E A5 AB 05 A6 8C 13 FC FC
 91 A4 25 DF CB AE C5 E4 D2 C8 99 B2 99 7B EF 61
 F7 22 1C B2 C8 AE 84 B1 D7 96 AE 4F 89 BE FA 08
 0F E8 F4 F3 FA 46 62 27 30 D0 5B 69 05 BC 60 65
 25 9B EC 94 5F 35 AE 68 72 46 39 F7 4A C8 98 AA
 53 07 72 19 4D 9B 77 FB 8A 31 A3 E7 D4 BF 7D 80
 A5 80 D9 0C 6A 67 F5 C9 F7 09 2C 76 92 6D CC F0
 05 2C C0 3A 55 80 BC A1 28 8D E5 E4 06 2E 70 AC
 74 8E 81 3C BA F6 98 5F 8E 05 7A BF 86 B9 69 83
 05 BC F3 D9 BD 5B 8A 6A 6F 34 FE 23 A6 E5 A1 6E
 CB 10 54 85 FE B4 9B 53 3A 39 58 D3 0E 4A 83 25
 1B 03 1C 15 AB FC BC 04 06 EA A4 45 65 BF 0A 2B
 15 1B EB FD 94 B2 8F 9A 96 7F C1 BE 8B C9 65 88
 3A 09 6C 4C 48 F0 6F 36 F0 FA 41 2F 33 D3 6F 33
 B7 C4 BE 7E 02 54 56 48 89 C9 8F 81 D7 B5 31 A8
 2A 0C D9 AE DB 92 5D 5E 12 BA 85 CC 8A 59 80 66
 E4 06 98 25 E5 B3 08 5E 17 07 CF AB 78 72 EE 83
 BF 64 13 90 16 C5 AF C9 01 9B 6C 13 53 69 EB 76
 0A 54 3B 54 BD B0 94 95 8A D1 FC A7 3E 36 0F 86
 13 D1 A0 A5 0A A4 83 7E E3 E9 EC B5 CA 11 CA 25
 FE 13 1E 1C BB 00 FC D1 D2 F2 3B 06 70 6A 31 FC
 1E 1F 91 51 95 C3 E4 F5 86 9F C4 5A 44 A8 2B 13
 A9 A8 8E D9 7C 25 BA 40 D6 C3 F9 D0 BA 2B C2 1B
 F6 86 97 06 5D B3 DA F5 8F E0 7B AB A0 03 E9 FF
 60 5A 8D 06 3E 91 BB 10 89 9D F7 6F E2 15 EC 9F
 85 02 4C 81 A6 B2 2F 38 9D A8 97 BA 5E D7 14 35
 08 F7 FD C9 DD 1D 02 9A 3F 1E 79 CC EC 14 33 FC
 3D 71 D3 F8 A3 6F 07 C8 E0 36 F3 E1 12 1B 91 BA
 F7 98 76 92 B7 39 6B 8B 03 42 84 99 30 F5 A7 27
 E6 CE 88 F6 8E E3 BA C4 E2 A6 5D 45 80 18 DD D8
 9B 65 54 07 28 62 A6 5D 20 98 D1 8F 21 FF B1 5D
 7A 4D 7A 9B D8 89 74 E8 0D A1 11 B7 35 F2 13 CE
 6E 39 4B 67 8C 6F EF 1A 5E 6D F2 AD 2F 84 B3 79
 72 7A 24 32 8C E9 8C E8 4C E7 72 3F 9C E5 E5 0B
 34 7B 50 53 5D 32 E8 C4 50 BC 77 9F A1 22 5C ED
 BE 10 DB 12 43 50 33 CB 10 3A A3 AF 82 6D 96 E6
 33 E4 1C A4 5C 5D BE 9B C5 0C 44 E3 55 A1 BC 78
 F6 EC 0F C5 63 59 04 C5 3E 68 3B 2F 36 7E 1A E3
 B3 F5 88 8F 5C 0B 04 13 E0 85 9F 61 3A 23 D3 65
 F2 58 66 69 D3 62 56 18 0B 22 2E 47 FA 19 33 FC
 30 C0 1D 5E 05 81 52 EE 07 51 57 B5 C4 A4 AD 01
 57 36 E7 43 8E F0 50 BE 2D 51 EB 78 96 D6 83 33
 A0 89 59 4F 5D 6E 1B 65 45 B2 3B 5D 97 76 CE B4
 EC 46 E2 5E 3F F3 E5 88 CA D0 E4 44 4A 76 A0 39
 D7 33 DE 2F 70 6D DE D8 2D 59 BC 06 22 86 96 E6
 DB 91 92 2D 8B 66 5F 05 2E 0E A7 96 66 DE 30 D5
 C5 68 07 6B 68 02 01 3F D2 7F 0F 5A 1A 64 8A 25
 2C 32 DD 7D 99 C3 59 67 9C 65 01 BB BE 2A D2 19
 11 92 2C 27 7E 47 6D D9 8A C9 D8 0F DA 0A 1C 58
 07 6B 37 68 B4 BD 29 27 31 D3 F6 D3 CA 84 57 2A
 74 63 6D 84 E5 9D 85 F2 90 19 04 12 5B 04 A4 3B
 C5 DE 03 20 5B 63 18 5D 43 AC 69 43 4F 97 C0 77
 3E 10 92 F8 D9 2B 00 DB 11 54 1A E4 C0 4E 8B 38
 1A 43 40 0B 0F EE 44 1D CB 97 3F 10 39 D0 2B 0C
 C1 8D 89 78 66 36 B6 E3 FD 3D BB DD F6 EE D2 EE
 79 41 E8 D8 67 75 C7 C9 5B AB D6 B0 14 1D 16 47
 DC 5B 4B 50 39 DA 3A EC EC 8D 6A BA 42 7C 6F 88
 B8 DA 26 A8 88 F8 CC CF 4D A1 B7 FB 33 D2 5A 2F
 05 8D 20 05 23 13 10 D6 30 40 F5 1B 65 90 19 91
 F6 8E A1 51 49 85 78 85 5A 70 11 E8 B3 90 53 60
 4A 89 A4 03 B9 4E 87 B2 16 7D 09 5A 3D 06 84 19
 48 B4 C5 68 C7 94 61 C6 C3 02 53 A1 31 0C D2 93
 D9 FE AB 35 64 9F A9 42 C3 FF A6 75 66 A2 36 81
 BA A7 29 F4 6A 63 2F FF D0 F2 14 E8 8F A2 83 90
 67 E1 57 AB C0 97 B6 93 D5 B6 AC E8 F9 88 0D 0D
 37 86 A4 9C F2 68 34 0F 98 A1 7B A4 AC 69 AC 91
 3C 64 29 87 69 21 87 C1 F8 8A 3F D5 0A FD 10 73
 00 42 AF 0D 4D F1 1B 17 28 11 75 A9 C3 A2 C6 A4
 AE 82 BE 7D 83 69 CF 8C 30 7F 73 DB 40 69 E9 0C
 6E 77 32 13 C7 DE 49 86 DB BC D6 D7 0B DC 83 D4
 32 0D 08 0A 80 36 92 C7 B0 BE D2 E3 59 0A A7 02
 42 7A 84 2B 17 65 D5 E5 4C 3D D1 B5 3D 12 C1 A5
 1C 48 6A 40 29 BC 1E 2E ED 36 45 6D E1 65 FE 40
 10 A8 22 85 B3 BF 9A 1C B6 8E 00 93 42 87 1A 19
 CA 24 62 2C 50 F4 86 BE 66 4B 06 E1 B6 06 C1 3F
 FF 7C F9 CA D2 B0 5E 82 C1 4E 34 C6 B3 0B DC DF
 5C 04 07 65 4C DF 11 C0 47 EA A3 F2 37 4F DA AE
 62 37 2F 3C C3 F4 DE 92 72 0D D8 7F 43 0D 5D 48
 B6 77 66 00 4A E2 77 A9 25 1C 5B BB FF E6 31 74
 B1 B8 50 67 5F B7 45 50 07 0A 60 46 4C 7C 8D 34
 E5 BB 82 FE 80 D5 74 D8 60 9E FA 9F 5B 3F 25 48
 EB F8 A0 B4 08 35 77 E0 B1 A2 A6 36 96 59 6C 8E
 18 D6 A6 7B E9 F1 72 1C 68 FB D6 87 B9 A0 7C 03
 D0 68 B0 31 F2 3D E2 7E BA EE 92 61 1C DD 1F 29
 7A 95 80 89 82 9C 0B DA 2E E8 8B 1A 51 94 8A 95
 44 B6 C0 22 4D 56 FC F3 0C 76 4D D2 D5 09 A7 FB
 61 64 C9 F0 DE 64 7D BA 9E 64 D8 95 2B 03 F7 58
 46 AF 7B F2 A4 51 6D EC 0D 9B 92 5D D9 CB 32 8A
 23 B7 5B C7 92 53 5C 88 97 96 DB 23 DF 21 26 21
 13 E0 91 9C 7D 1B 59 01 C5 38 86 13 53 59 28 2F
 89 01 11 56 1C 26 D1 16 7E EA 0C 90 3F 47 D7 22
 C0 E8 1C FD A4 9B CE A6 F0 8E 0E B7 24 9B CF 7B
 26 8E E9 B0 BD 59 69 C3 6B 9D EC 0A 15 44 4B FE
 C5 EA 3E F1 D2 42 53 AD C3 06 AD D9 8D E7 B2 A1
 A3 A0 C8 C0 8C 04 B6 2E 6A C9 BE 44 12 2F F7 AD
 32 D3 4D 77 8F 7E 26 E2 E9 3A 6B 6D 6F 6D 71 F0
 41 71 CE 49 F9 EF 4E E4 C6 4A 73 BA 30 C3 2A A3
 D3 6E C6 64 62 50 64 37 6D 08 23 2F 2B CE 5B A9
 9A CF AE 63 7E 6B 16 94 E7 DF 1D C5 C1 95 01 23
 CF 9E DA 68 B0 76 1D BF AD 98 35 BE 71 7E 69 CF
 D9 2D CB 7F D6 3E 6B 4D F2 A8 AC A0 1D FD 48 79
 B0 DD 60 9C 35 C9 A6 86 9D 49 67 40 C3 A7 D7 F8
 52 FA 49 55 A4 9D 8F E9 85 1F C6 62 0E 98 62 80
 DC 90 0E D0 57 6E E5 A7 89 10 7B FF 2D C1 E8 CD
 AB 76 D1 28 E5 90 59 75 84 67 95 C5 8C CE B9 87
 6D 5D 88 4C 70 DA DC 7E 20 2C 01 D0 7A 3F A8 82
 9E 0E BA 1D C1 F5 6C 0A 74 60 29 2A DB 9C 59 0E
 DA 46 C1 A6 F4 14 EE 03 D1 F4 C7 58 0E 7F A4 07
 70 C3 6E 79 79 AA AB 37 51 74 4E 65 41 9F CB 67
 3C A0 B6 E6 AD B5 3B A2 C8 B8 D4 E8 EC 28 05 07
 69 6E DB EE C5 AC 45 80 C8 61 6D B8 F4 0B D1 C1
 B5 AF AC 54 5A EE 7D 20 B2 FE FF D4 2A 4D AF AB
 AA E4 A7 52 87 EB 13 93 B0 B5 DC B8 CC 7F 3D 1C
 9D F9 3E 5E 1C D8 E8 22 59 23 68 ED 1F 2D CF E6
 3C CA 98 A1 51 52 71 4C E6 57 6B 45 50 D1 5E 15
 65 25 EF 98 0C 54 DF 5E 47 86 5B 7E 9F 51 A5 8B
 B5 A1 E0 FB 13 6D 4C D8 D9 05 3B 6E A8 6E 3C 67
 0D 2F B8 93 2D E2 99 CF C0 A7 72 DA 93 9B B1 3F
 2C DD 3E 06 66 06 E6 A9 8E 49 A8 7F 44 A4 D5 61
 D8 EE E9 1B D3 AE 75 53 55 66 FA 8B CF 0A DD 28
 3D D5 58 84 7B B5 A3 A3 47 38 F1 AF F8 9A 71 16
 C5 5E 53 A3 54 2B 02 BF 69 90 7F F7 55 DA 5E B4
 AD 85 24 F6 27 72 52 9F E8 DF ED D9 83 74 9A 7D
 32 07 D2 2D DC 9B 04 D7 0B EF FB 97 9E 65 0D A4
 93 B4 34 13 71 96 FB E1 1D 52 43 1B 35 99 C9 1E
 76 FA 48 3B 79 44 23 9D E2 2D F5 F3 ED CA 45 8C
 BF 14 9C 86 81 0F A2 9D C0 20 86 5F 55 1F 37 A0
 D2 75 11 91 0A 85 72 AB 1C 04 F4 A0 E7 24 1C F2
 22 EF A7 7E 76 D1 68 62 67 41 08 9F F7 87 4A 0C
 AC 2D B1 9A B2 9E 6F 64 9C ED E5 4F 2A 06 AA 9B
 61 A4 39 C0 21 A4 2F DC 25 6E B1 BD ED C2 1A 65
 39 76 40 80 86 B9 F2 78 46 29 F1 9E C7 29 64 DD
 E2 A6 34 9C 06 A5 49 6D E0 C1 F3 F0 8B 33 11 E0
 7D 3F 29 9B 16 5A ED 30 F7 6A 32 C6 B1 A5 84 3C
 59 F9 6B 4E 68 33 6E 2E B6 87 AE F4 5F D0 6D ED
 3F 1B 5A B6 49 B7 3A C2 14 36 E2 38 A8 AC 45 D1
 06 11 17 F6 65 2C 43 2B 01 D1 8D 2D 72 6D AD 29
 65 1C 90 96 AB 12 3B CE 1C 25 F4 F5 02 6B 80 90
 50 D1 E9 FA E3 4F 1B 02 C8 41 C1 73 E8 DD 5D 7B
 10 99 9C ED FF 07 89 CB 52 C4 3C 94 57 46 99 EA
 6D 59 F0 66 27 46 16 6C F0 15 1B 8E 84 DD 00 F6
 DF 47 F1 BB 36 E8 22 5D 2F A5 22 00 01 C1 1D F3
 A7 84 E3 74 6A BA F4 E7 DF 9B 41 84 E0 30 4A 47
 83 18 17 46 D4 ED 57 3E FE FA 94 7A 02 CF 4A 5C
 A7 B4 17 17 4E 7A 38 23 65 53 FA 87 F6 6C F3 56
 AE 4B C2 87 1C D6 37 CC 0F 66 EF DB C2 89 34 82
 B8 0B ED CA F3 81 F9 9F E2 3E FD D2 96 80 DB 16
 EA 87 51 98 E1 07 03 75 59 48 A2 67 B5 ED 13 72
 00 D7 B3 B8 E2 B7 66 B6 45 2C BC 57 2C A8 36 C5
 37 EC 2C 92 AF EC 4E 8F C2 BB D0 26 AC 81 0E 52
 13 85 5F E0 DD 58 A0 81 28 68 FA 5F CF A1 8C 7D
 47 0F 20 45 9F 1E 31 6A D4 FB 79 1D 98 68 2A 85
 37 D4 DE D0 A0 44 2E C3 CF 89 D7 C6 62 5E A8 BE
 09 CF EF 80 C6 6D C2 A9 5A BA FC 58 DD F4 69 5E
 05 4A 0D C7 7E 67 62 CA F1 A5 A8 6C CB 7E E3 3C
 12 E5 05 34 52 57 13 CD 5E 3E DF 63 AD 56 A3 48
 B2 C5 79 1D 54 50 51 DB 69 DC 58 CB 7F 1D 2F 0B
 C2 7A 82 F3 C6 AF 6D 37 87 76 D6 19 DA 97 63 6F
 3F 5B 28 A5 1B C0 98 A0 E4 50 26 E8 DB C0 D6 42
 3D 21 36 54 98 20 4B 41 36 A3 F2 58 4D 0E BD 03
 6E B8 D0 47 5F 54 28 6F 70 BF 39 52 7C C3 6B DE
 2C 6A C3 68 7D 38 7A 6C 43 BA BB FB 20 D9 72 7C
 A3 8F FA 0E 58 15 CB 83 A6 B9 50 AA 2A C7 69 3A
 E3 B7 10 D5 E3 D1 6D FF 23 4B 12 EF 0A 00 18 60
 BC D9 81 C7 C4 E0 F6 17 51 0A 53 11 B2 FE 7B A7
 59 6D 63 14 53 41 77 C7 2A 1F 84 E9 6E 15 B5 55
 EF E5 A0 CA 29 2B 27 A9 C7 EB CA 19 E7 9D 6B E2
 85 9A C1 7B 9F D7 61 2A 38 6B A4 00 78 7A 5A B9
 AB 98 BD BA 57 18 23 FE EC CA C5 61 65 65 9F 8C
 A0 15 DF D1 61 CE E7 6D 2E 4B 68 25 BF 75 C2 A2
 50 A0 F8 96 13 7E F1 15 09 F5 E7 9D 40 9E 3E D8
 34 9D 3D D3 C1 02 54 E4 E8 D8 62 5A EF FF 8B C0
 31 99 15 EE 43 1D 97 34 37 0E CD 68 81 42 AE 53
 09 54 CE 6A 36 CC 44 6C D6 28 E1 5A 26 14 71 55
 C5 74 B8 E4 3C 29 83 C8 76 A9 48 84 E6 5A F4 A8
 3C 08 19 90 23 DE 41 40 77 E6 D5 8C E9 61 AE 1D
 42 24 07 51 39 6D F8 0F FD 98 EA 49 CF 5B D2 C8
 22 E0 D5 F6 CD 72 E4 AC E3 46 FD 6A BC CE 8D 34
 D0 B8 62 67 8E CF 5E 3A 80 8A 1D 14 73 0F 30 44
 F5 01 76 C0 7A 99 AF 9F 95 A0 65 20 E1 BC F9 45
 CF 34 C0 FD 5F C1 53 C0 03 57 6A 7B 21 FF 44 9F
 37 9C 1A B5 5C B7 3C 2F A9 2A 82 AD B3 B5 4E E0
 66 75 A3 BC 28 6D 8C 7D E8 2C 5C 6C 60 D5 2F 2B
 14 4E CD 51 14 D4 AF 25 29 00 03 59 5D 45 FA E3
 0B 18 A6 48 C2 01 75 90 37 BD 46 17 91 45 9C DA
 B1 4A 9D EA 2F F7 48 CD CA 94 62 2E 7D 4B AE C3
 A6 A6 90 B5 F8 04 05 98 18 C1 79 D8 35 EA E6 A6
 FE 2A C8 D8 1A CC D5 36 7C 68 90 AF D6 B0 59 34
 19 A9 DA 09 F1 B1 83 33 BE 18 2C D9 DB 7E 75 07
 73 B6 39 05 2E 58 97 37 5D F0 57 2F 46 F3 99 F7
 DF 7A 14 53 9A 55 95 0E CE BE 4F 2E 38 A6 47 FA
 10 BE 8E D1 03 74 F8 84 F9 7E 94 41 AD EA 0A 63
 E3 77 B0 3C 3D 23 B1 C2 FB FB 18 86 91 09 F6 96
 28 82 64 02 63 D6 42 B0 D3 65 A4 97 68 08 2B 14
 DB C3 F2 3D 8A 9E CF AF 06 8A 04 AF 76 E9 EC 21
 07 05 51 41 45 B1 E8 00 69 3C F2 16 F4 A9 8D B9
 7E 6A 28 7F 5C E0 C4 25 06 13 AB 4E 65 3C 36 98
 6D 85 04 76 34 F1 08 A4 8C 1D D9 CF F9 0D E2 83
 E8 CD AB E9 5C AA 36 B2 F9 DB F5 B0 0C 6E D4 75
 65 E6 F7 F8 78 91 F7 25 FF CE B3 4B 5F EE AC DB
 65 76 4C C9 53 03 9C EF 9E 3B B5 C8 ED 15 54 23
 0F 7B 74 28 15 06 F4 42 6E 49 CC D1 07 2F E2 D1
 76 F9 D0 44 26 32 37 8F FE 80 4D B9 DC D2 80 32
 64 56 69 82 B6 6A 56 E2 96 1E 93 3A 72 72 02 F0
 6E 19 C6 D1 67 B7 60 ED BC 1D CF 55 18 FF B9 77
 81 44 98 F1 DD E8 A0 C3 07 84 4C 32 33 B9 77 D5
 8C 89 90 77 C4 4E D8 25 1F EE C8 CC 1D 62 69 01
 15 6B 81 FF BC 79 A6 07 D8 CA 11 9C D1 A1 C6 3A
 28 C5 B2 F3 AB BB F4 B9 77 81 FC 1F 8D 2F 85 36
 D3 C6 2D 9E F8 3A BA BF B7 04 20 48 D5 62 E8 32
 30 D3 EF 80 78 8C C0 C2 97 55 E2 C1 45 EB 50 FE
 56 34 1F 58 19 D7 5C 82 D6 15 52 AF 9D 61 B8 24
 BF C0 52 31 F8 BB 81 63 6B EF 4D E8 1F 71 AB AB
 DC 70 DB 0F B5 7D 8E A6 07 A8 A0 23 7F 33 82 C9
 96 23 B1 46 7A 75 24 27 7F 26 2D 6A 2D A8 81 45
 E6 D8 19 92 AC 2F 0F EA 02 57 3C 23 6E 08 B0 F4
 D2 AA E7 FA 65 E6 C6 4C 37 3D 49 81 93 C4 83 7B
 88 25 1F C8 95 CB 7E 06 F7 3F E8 C7 15 A9 11 9F
 9C 23 92 18 29 CA F2 8D 0B 5C 57 DC 11 E0 46 1D
 03 10 A3 D1 9F 12 08 08 90 19 CA E7 D7 8F B2 97
 A8 82 3D 1A A1 38 9B 65 F3 7F E6 B2 08 6E 4A 5E
 1F E4 00 C5 23 A4 CB 90 09 48 CF 11 FB 91 3C AD
 1A AF 2B 7A 7D 62 4B 9A C2 57 EB 4B 1C 14 40 E1
 B5 0A 0B 28 8E 04 C1 82 29 5F C9 1D 2B B2 76 B8
 CD D6 D6 45 E1 DD 1A 0F 2F 6A 76 FC DC 88 41 BE
 BE 8C A9 A2 D0 2E DB A1 B8 5B 00 6F 46 73 3B 41
 31 F5 E8 87 CA EF 82 3B 6D 4D 50 DE 4D 07 D9 1B
 08 46 6B 6A D2 56 E9 7A 9A 03 58 D0 AE 19 12 64
 4B E1 60 03 AC E5 3F 3B F3 C6 97 F6 F2 C1 03 54
 72 B4 C2 31 12 1A BC D5 D5 DE 60 4D 4A AF E3 24
 FE 4C 00 1E 26 68 C9 A9 2B D8 FA 3D 02 AB 99 C8
 A9 EB AC 62 9F 0F 1A E0 D4 0C 2A AF 0C C0 10 AB
 33 14 79 5C 4A 85 8E B1 DA 55 6C 5F 10 11 62 4F
 5A 1D E0 60 9A 56 23 D0 B1 30 B6 41 C3 7F 75 23
 32 0A 47 97 03 D1 C9 6D FA 3F 58 AF CD B9 FC E9
 62 2C 6E 52 C2 BB 8A A3 E4 AB 21 4D E2 BE EE 51
 35 C5 22 84 3F AD 05 69 C0 08 11 00 91 91 CD 02
 88 53 47 3C 9B 92 5E 9D F8 EF 44 F7 63 00 4D CD
 90 AC 34 09 13 C5 D8 94 98 EC 8F 6A 07 96 AF F2
 EE 06 6C 3B E7 AC EB C9 71 BF 9D 6B 4C 49 A6 9B
 A5 F1 99 01 C1 72 14 DA 5E 95 CB 37 ED 9E 75 32
 9D 16 A1 E5 88 01 50 BF 22 84 80 C0 E6 88 B3 89
 EC 89 5F 9F A1 2A 31 CE 92 39 38 80 18 4A 90 58
 F7 31 6C 67 33 0E 32 A8 9D 67 C1 41 1D 99 2C 65
 3A 27 30 BF 95 20 7C 69 B4 AC 88 03 03 42 F9 D9
 E9 31 1F 3F 61 9E CE 0B 9C 7C 64 BF 4E 25 D2 BF
 80 F4 A7 64 FF 72 A4 B8 8C 0B A9 32 DB A5 03 2E
 EB ED 7F 3B DC B0 EE 9B F6 24 59 B9 F6 42 03 1E
 3B 49 FA E0 27 49 D5 4D 59 1C 0C 4A B5 8B 85 F4
 29 2A A0 01 D7 DB BC 36 E1 65 B5 A4 C9 C5 BD 4B
 4A 48 AB AC A7 66 4E D3 24 AF B0 E7 96 2D 7E DE
 9A 65 EF 83 1F 0C AE AD 10 33 40 4E 2E 9F A6 F8
 1E E7 E4 4E 20 9A 85 E4 6E E5 DA 45 58 DC 02 03
 12 D1 07 55 45 DE 23 5C 02 5D 28 0B FD FB 27 2F
 C6 C0 AD 0A 0A 84 89 69 68 94 39 FA DA 7F 6E 53
 0D BF 12 BA C2 C4 9A 61 1A B4 7E 51 50 15 A1 F4
 54 17 F8 89 11 C0 37 65 0C 51 7A 2D 98 AF 7F 22
 09 C6 5A 25 7D CD 96 9E 4E C4 73 7D 4E EF 79 5E
 A7 C9 05 E3 F9 93 2D 45 C3 56 E8 BE 18 E9 F8 2D
 9D DB F2 20 64 92 46 92 48 D7 A6 55 0D 2A D5 4F
 EF D9 8C 64 89 49 B9 F3 C6 B7 30 EA 32 FC EB 5C
 57 C9 E9 47 AE 2F BD 49 61 61 EC 0F CC AE FA 12
 F8 DB 7A 7F 2A 23 01 40 A9 82 9E 88 6D 6A A6 23
 0C 5A A8 0B 4D 9F 16 BE 81 58 03 82 72 E3 61 C0
 7F E1 DF 84 06 F4 46 EA 36 DB 80 B0 AF AB F3 6F
 24 6E 77 BC FC 39 7C C4 88 3F F5 CD 1A 3B 94 9A
 7C B9 4B DD 0F 1D B1 D3 41 64 7C 19 FB 7C 99 CC
 AC 64 58 A2 CB A7 E3 81 09 8E 34 7C 7B 39 9E 66
 20 79 AF DE 7E 35 14 31 C0 2A 5F FD 06 BE 1B 44
 9A D0 C2 65 A3 F2 7E 13 B8 A7 6B CE 12 C6 B5 91
 60 A6 2A BF 7C EF 7E 9C 4E E8 7E 6C 07 B0 69 77
 22 76 35 1D 72 0D 99 CA 61 E6 8E CC BC 99 E8 47
 05 8A 93 72 46 87 07 EB D3 E7 FF D1 86 A0 C9 54
 1C BD C4 E9 4F 76 32 07 89 8C 74 B4 6B 1D 1A 86
 89 B0 1D 89 A8 FD 5F E8 6A 9D 5C 59 8E EA 1B 45
 5A AD 5C AB 6E 2F 90 4E 8F 5B D7 18 A5 32 EC 80
 8D B6 AE 49 AD 57 7D 43 2B 77 77 EB 90 87 7F 4B
 DF F0 A7 66 F6 02 53 D9 91 BD 37 81 7F 37 DA 6E
 FB E4 94 9F 45 70 DC D4 1A F1 F4 A0 BB A4 31 E8
 89 C9 D2 29 AB 32 17 42 1C B0 5C C0 27 52 55 24
 22 9A 87 9F 19 5F 18 99 4E EE 98 04 FB D0 95 8B
 51 A1 3E B2 E7 B6 1D 2E A3 91 7C 5D D3 31 A3 C9
 CD 4A CA 5C ED 55 28 74 BB B5 43 7F B9 0F CD F2
 4F ED FC 10 87 1D 6F BE 16 54 0C F5 E8 14 BD 89
 0F DA 03 5B BC 2C 5B A8 BE CD EA F0 14 C8 15 D0
 55 35 5F D8 52 72 A9 78 28 07 A1 47 18 70 9B 77
 3D 72 65 D5 07 67 CB BB D1 F0 98 61 69 95 B0 FB
 B6 AA D3 5D 7B 24 B3 C7 28 6D EB EC DB 97 DC 0E
 3B C3 FA D8 E3 DE 92 4F 1D 43 5D 94 B2 3D F7 BD
 9F 10 A1 9F C2 20 26 25 B4 26 7D 69 EE EB 68 FA
 90 47 9A 11 06 6E 55 58 E8 A8 86 7B B2 04 2E 73
 13 4C 3E 5F 9F 25 6F 9F 20 94 F5 70 2B FF 22 32
 7B CA 02 9D 7A AB 59 6F 16 94 8A BC 7D A5 2E 14
 D7 6B 8B 8C 05 61 C8 11 01 32 19 F1 6A 9E D1 87
 C3 EA 69 A0 58 70 93 7C C7 68 77 E1 3F 60 B2 3C
 7D 15 DA 2B EF 82 B4 1F 1B D2 81 DF ED 82 A8 60
 13 2E 83 55 3E 4E A9 46 9D 21 C8 E2 40 4F CF D6
 9A A9 DD 4E B0 5D AB 2B C3 D7 C3 14 6B 9E 12 D8
 A2 E3 06 32 0B C7 59 92 27 DC A6 8F AB 4F A0 54
 84 1A FD 54 02 34 3A 27 BB 12 95 36 43 46 58 23
 56 2E F0 4A 17 F2 29 30 CB B1 3D 40 6C 63 CA 17
 4F 7B 47 F5 F4 42 BB 54 1B 8E 2D 68 D5 53 DE CF
 0B 14 4E DF 5D FD E8 C6 DA 21 7B DC 6D 74 38 46
 78 71 B5 A0 12 F3 37 92 DE C0 42 DE E1 6C B0 25
 A3 37 88 E3 B8 F5 4D BA 4C E2 47 D5 01 C6 A7 89
 06 D2 99 59 03 24 82 6D 80 C4 8C AA 9C 2B D6 F8
 E3 D8 15 1E B5 E4 18 3D 44 84 26 D6 73 B1 36 EF
 98 B5 64 B6 F0 29 82 01 C3 39 54 5A 6C EF 21 DA
 C6 18 7E 27 76 86 C3 3D C7 8B 3B E5 03 34 E2 09
 4F 09 7A CC 3E D7 3E 1E B2 96 5B DA B8 73 96 67
 04 5B 96 C5 4A 18 5A BA B7 A6 95 3A 38 DC 99 4A
 BC 04 71 A5 D3 FB 23 90 C4 24 DD F0 61 05 D5 9C
 59 71 DD 42 62 6F 1C 6F D9 D6 E6 FF C7 14 87 6F
 6F 3D 40 8A 9D 75 DD 58 E8 C5 FC 92 F1 20 D3 BA
 08 87 30 CF 1F 6C 8A 86 AA 61 24 FD 3D 99 13 C7
 F4 3B 5E 46 EC A8 17 81 E4 B7 40 87 F2 F3 CA C4
 75 83 DC 57 F4 AC 64 E5 CF 27 46 71 49 0E 0B 0C
 F0 22 FF 77 54 BC 02 69 AE 29 08 A5 F2 A0 2E 4E
 B2 A7 CD BA 31 ED 03 BA F6 34 8F B7 65 35 D5 95
 22 82 AF 88 E7 FE D3 FB 1D 8F C3 01 CF 83 58 32
 72 E4 0E 4F 20 EA 2E F9 5F A5 1C 49 97 D7 55 11
 6F 11 F1 75 8C F2 F6 B5 FC F8 4F D2 42 EE 99 E9
 DD 6C 75 4A D7 1C 76 C6 6E 03 FC BE C2 72 9D 10
 2A 68 7B 4C B7 26 60 97 31 3F B9 67 D6 E9 DA EF
 BE 25 C8 0C E4 4B EF 02 23 23 AF DD B8 83 02 A5
 B9 79 7E B7 BE C7 47 06 C8 4C 1F 15 41 85 2B 7A
 28 EB EB C7 E4 E2 28 A0 23 D7 6B C8 21 67 2B B2
 81 24 0E 6A 77 90 D1 1C DE 27 B7 CC A1 F9 7E F9
 12 4C 2B A9 7D 27 48 8D 1F 9F 3B E6 C9 49 3D B5
 A0 8D C5 CC 51 B8 71 E4 54 29 06 21 E7 DE 26 70
 E6 2F E9 90 0F F8 9E E7 C4 FF 1B 52 D1 87 4C F0
 D1 42 D6 27 57 9F 01 85 9F 1B C0 2F 58 C9 4D 21
 89 3B 5D 86 AE 23 EB B9 FB 76 17 1D 42 AC 4F 87
 17 31 4A 3C 55 C7 BF 8C D5 2B 1B EC A6 1D 66 60
 C0 3B DC 28 58 12 56 90 1D B5 E0 ED 62 C2 E3 22
 2D 6A 99 C4 AF 7B 03 49 DA 7F EA D1 27 D3 C1 A0
 22 D1 B4 5F 4D 9A 33 69 C5 C6 A9 BE 32 BF BB 2D
 31 A2 31 95 21 18 C8 94 B1 B6 72 A6 6B 05 97 14
 5E 58 F2 36 7A 39 08 1A E8 2F 4A 7A 5D A6 E7 E6
 11 C7 EE 16 52 CD 61 D5 1F 13 5F 44 75 A2 26 DF
 B9 A1 67 E3 F8 61 2C 9A 3C AE 6B 43 57 59 C5 B5
 AD F6 38 31 EC FC 06 69 A8 53 FB 2F 04 62 96 1D
 6A 0B A2 59 69 8F 43 C3 13 A3 0B F7 33 4C 2D 46
 65 38 A0 F0 52 EA D4 CC D7 72 09 0A 20 9F DA 9D
 F0 65 23 6A 9F EA 65 86 44 72 12 72 00 EF EC E8
 F9 95 52 8E 1A 8F 15 74 2E 1A 9B 6D AF 2F 9A 28
 BA 78 2D 81 20 BD 1A DC 42 63 87 7A 5A EB 4E 17
 1C CF BD 68 AC AD 8E 36 51 9A 90 66 3C 18 93 44
 E1 08 7C 91 0B 98 66 C3 98 00 BD AB 51 02 73 2B
 BD 7B 6D 05 73 FB 2F 3C 9D BF C0 1F D3 67 66 38
 35 6B 7B 04 7D 72 A7 0D 29 2F D9 B0 87 74 06 0D
 57 80 9D 1F 52 08 A0 08 C7 20 E4 51 3F 9F 05 98
 C6 6E D2 57 74 9F 0A 66 81 F7 42 06 5C 19 E2 E3
 72 F0 78 F9 E3 A8 2E 9E E6 48 4F D9 6D 6E 60 52
 D1 34 03 34 67 2F FA A0 CB 82 16 E3 AA 4D 03 5D
 87 61 70 CB 9E FD F1 85 7F 1B 2F 05 2E 5E 17 AD
 DA 39 DA EA 61 04 DD F0 F9 AF A5 25 B8 64 98 1D
 92 7F 2C 5C 04 E0 1C 03 0B CE 96 44 2D 50 5A A9
 E0 AB C4 2A 7B 8F FE 63 12 72 F4 2E AE 82 4E D4
 D5 68 B4 6E D0 3A A0 92 D4 0F 7F 93 51 38 70 91
 D7 D3 59 53 5B 26 0D 44 40 A9 EE E4 13 0B 3F B1
 F1 6B 34 BB DE FB B9 F9 D0 38 D9 F9 3C C9 74 19
 08 31 1C 12 02 61 E5 12 2B 48 91 53 E0 EF D7 B3
 20 F8 F2 1A 9E 9C 3C 55 54 A0 5D 85 BE EC 2A DD
 D3 39 9F E0 1D 5A EB 85 26 94 D9 84 F6 90 CF A9
 99 EE 4C AE 34 9B 7C 6F 52 AE CD F2 8A E1 23 5B
 0B 16 35 0A 79 DD 3C 7E 2D F0 71 FE 21 B7 65 3C
 C4 E4 6E B1 E9 67 10 1F 49 F5 19 6F 70 87 31 AE
 37 14 A9 9F F4 E9 FF F9 9B CF A5 4C 5A 29 78 22
 D3 AB A9 EE 59 99 4A 16 61 98 D8 2C 62 C5 B0 A4
 95 E1 09 BD F7 40 A5 55 DD 15 22 14 80 88 7F 18
 50 1A D2 7C 7F E8 A7 46 CD BB 6B 7F C9 67 DC 34
 EF 24 BC 85 2F 33 9D 61 4B 7B 3B 53 90 4C 10 73
 10 1E FA AF FD 1C 09 6A AE FE 9E 52 F7 CF 21 E7
 60 CE 67 23 D3 66 30 35 71 E7 8F A9 FD 3C F5 BC
 DD 08 CE ED E3 2E A3 AA 86 6C 23 BB E9 43 AE 29
 62 BC E9 97 43 5C E1 AE C1 A5 BF DB E5 2B 2F 1A
 1D 73 79 AE 22 A3 1E 69 63 CA 9E 13 D6 5C E3 E8
 64 E4 A4 CA D4 E6 0C FA 60 F8 55 EB 13 FF B8 A8
 5D 64 63 61 62 9F 13 13 68 B7 3B C4 93 E3 4F 15
 E0 6C 2D 9F F8 F5 FD BE 29 E7 82 88 D0 8C 98 5D
 D2 24 86 05 87 BD A6 1F 18 A0 CD E9 82 BF E7 96
 46 9A A2 1F 16 50 01 6E E4 32 38 01 DB 1A 85 E8
 3C A8 8C 1D E9 E6 29 26 D6 F6 DC 1C AC F5 3D EF
 FA D7 37 21 59 FF 1D 2A BC 97 91 22 72 6A 03 6B
 74 A5 0D 53 98 43 3D 52 71 11 81 EE B1 DB E1 B7
 54 83 B9 0D D6 7E 12 64 1D 94 1B A6 DA 8B F5 FA
 C1 78 5A C1 16 1F 8C 44 81 6A 87 DD 02 6A F1 CF
 41 04 B0 7B 72 B8 FF 14 85 39 F0 3B 72 33 32 37
 31 BA E9 07 CB 05 59 30 01 7C 0D 9F C5 D1 68 49
 A4 C8 6F 3E 31 60 A1 6E A3 0A F4 A1 90 FD 6E 9E
 C8 E1 E3 52 F9 72 B7 FB 4E 00 0C 18 5F 51 4A 1B
 61 34 2D CB 19 91 C5 C4 4A BF 0F 27 59 A8 81 94
 D3 A2 53 2F 48 F5 12 71 BE 42 04 EC A5 A1 FB 8A
 E6 6E 2C E9 61 54 D5 EB 7B 82 6F D0 6C EC 37 90
 62 FE FE B5 D2 85 F6 47 69 3C CB B0 1E F8 04 E9
 5F 01 A0 3B 5F 89 FA 04 1D 51 75 4D FF F0 A7 59
 FB A5 7C B9 AD 38 8D 4B 8D 66 69 54 27 98 6A F1
 25 78 29 EE 61 77 0B 1D 2C C5 09 0A 12 25 60 ED
 BB C7 96 B2 7E FA 3F D3 B6 F4 1B 1B 25 D0 33 4E
 A5 B5 2B A7 18 D4 C7 95 4F 9F 94 84 5D 25 D5 E8
 65 11 32 98 E5 67 84 1B 69 33 14 6E 98 6D 81 58
 6E 3D 40 45 90 C3 08 E7 FF 2E 2A 0F B6 B1 0D AD
 E0 58 02 68 44 ED 2E D1 2B 59 59 EA B9 AF 7D 26
 0D 11 DA F4 57 41 FB 4A 0A 2D B0 D0 C9 F9 8E 48
 F8 E4 56 90 C1 47 D3 63 BB 0D 1E 0C A9 C5 54 81
 98 5C E0 10 E7 35 BB 4E 68 13 E0 D1 55 2D ED 18
 6C 94 8E 01 9B FA 20 52 8B 4C F0 ED 05 4A 18 6B
 0C DB 65 0A 98 D0 47 83 FD EB C6 98 8E 09 8B 44
 3D 65 3F 55 3D 92 FC 58 7F 65 00 0D A8 1B 1A 59
 E0 E5 55 E3 BC 3E 7C AD 08 FF 76 69 DF 1A 87 63
 EC EF 60 16 D4 B2 8A 91 3F 99 84 56 58 10 86 D3
 CD CF 45 94 B6 53 0D CB BA 86 45 F7 3D 30 52 6B
 6E 91 CE 6C A3 06 37 3D 75 62 22 86 22 0C 21 F4
 76 2C 78 B6 B3 A1 46 A1 CF 4F 5F 60 A2 33 23 D5
 DF 99 10 D9 F8 FF AE D3 C9 E5 97 C9 86 66 46 F8
 A0 B2 B0 6B 8A 04 DB EC 79 EF C1 09 B1 D3 F9 D2
 A3 51 76 8E 64 51 80 AE 1C C4 DA 4D 95 BE 53 34
 AF 9C FE 1D 89 11 58 DF 53 24 3E D2 17 DC 7F 71
 2B 09 7F B1 C4 9E 69 14 16 A7 C9 78 90 5A FA 78
 7E 0D 08 8B D4 35 9F 45 7F 0F 04 9F EF D2 C7 6C
 22 26 F2 73 C4 8F 33 E4 65 0F 5C A0 A3 73 B1 DC
 7E 5A 94 08 72 79 5A 98 DC 94 D6 1F 61 59 97 66
 A7 D0 C2 6A A0 44 D0 F7 00 B5 85 A7 8F 90 C5 B0
 A0 7D 1D 51 84 0D 96 46 22 52 BA A4 CF 69 72 6B
 97 AA AD 0C 53 E2 34 A2 E7 F1 05 CE 8B FB D8 B9
 1B 04 DD 52 A1 D9 E9 5E 47 BF C3 F7 A7 E5 FA 5E
 14 55 0E 0B CB 1D 0F 05 EE AD AA D4 21 77 12 48
 9E 61 86 8D D0 60 91 00 86 A5 04 FF 04 AF 6C 0F
 45 34 29 82 C5 D6 E0 88 C2 3A 60 B3 D5 F2 C5 58
 62 F8 E9 F7 96 69 58 00 E5 D8 BF 90 62 22 57 81
 47 9D 9E EE 33 89 05 2E 7C 85 7E 87 6A 04 E2 70
 5C 02 F4 DC 18 58 BE DD 38 CB 7D 17 C6 AA 96 16
 59 DF 02 2E 9A 4A 7C 42 28 3F 3A B1 BC 60 2C 73
 42 D2 CA AE 00 B1 8C 56 16 52 8D C4 B1 06 FD 4C
 46 DB C7 EC 19 9D B5 61 57 1F 49 9A A1 5C F3 FC
 82 BE A4 66 06 1C A8 6F C4 A2 91 E2 19 38 4A 8C
 2C 24 2C 26 1B 77 54 05 58 93 54 B5 50 DB 4D B9
 86 4F 7F 99 71 D9 57 72 1C 37 5F 78 26 F1 05 F3
 63 92 93 3E B0 75 39 35 09 5D 04 8C 86 19 12 4B
 8B 94 F5 AF A2 04 05 3B 07 0C EB 0C 71 6E F8 03
 96 94 9B 47 6E 93 2B 88 A6 5F 2E 08 61 25 34 FD
 57 51 56 11 6D 58 01 90 D9 4A A9 41 1E 67 E4 10
 64 7F 33 12 D5 D0 85 2C 88 F2 7D 80 2E 1D C2 8D
 D6 39 7C 34 DC 9B 92 55 31 6A 24 CB CA 04 42 EF
 86 87 96 DA E3 08 AE 83 1E 5C D4 73 64 1E DC 85
 6F 96 7E 59 C3 A5 09 D9 EC ED 1D 7E EF 7F BE 8B
 BA 5A 6F BD 05 AE A4 D0 34 9B 67 FE 89 D4 84 06
 4C 7D EB 6D C7 55 28 4F ED 9A 1D 5A 34 D5 E8 9E
 F2 20 75 67 65 57 6C F7 01 2E C5 98 55 51 64 A6
 7D 54 26 A9 72 1C EF DD A1 89 18 EA D1 9A A0 98
 54 FB B9 A9 5D A8 62 CC 82 3D 3A F4 79 B2 FA 44
 D7 83 A6 93 03 EE CC 4B F1 64 93 9B BF 34 59 A1
 DD 1C 70 57 94 7F FD 97 BC 03 D8 89 5D BA 71 68
 BB 50 87 11 22 F0 9D A8 62 C1 DB 8E FC 88 2D 3D
 8C BD 74 6D 30 7D F9 3E 5E C6 30 00 18 D2 17 F3
 FC 43 F4 8A 63 8A C3 38 AD 79 E1 44 34 2F 60 97
 8E 2C 47 24 A9 F2 B9 C0 F5 FC A1 FB 91 1E 2C 58
 58 35 B8 B6 66 92 1B 79 F5 3C CD 3A 94 C1 14 50
 CD 09 C8 45 FD 33 D6 C6 37 BF 65 7E 8D F2 4E E7
 ED 50 CE 1B D5 7E 03 2E CD 73 0A 13 B1 E8 22 AC
 69 F2 C1 C4 F5 D8 BC 8A 8C 08 D1 85 EC AE E4 61
 C9 74 41 54 D2 29 00 3A 5A D3 2B 41 ED 50 53 16
 CA 59 26 52 EC 99 30 F8 5D 41 B3 AB 78 2A DC 30
 F7 05 32 08 73 5D 7E FD 24 92 7A 79 B8 03 AC 09
 73 2D 78 E0 AE 2C B3 2E F2 2D 57 73 15 E4 C9 A6
 A4 FD 6F 56 8A 89 5F CD 1E 45 3F 10 5C E9 A7 D4
 FF C3 9E 47 94 3C 6F 42 0E 77 A9 29 60 98 2F BF
 43 27 94 2D 43 2C F6 6C 09 B1 A8 40 69 24 83 7B
 A7 97 27 39 60 84 2C BE E8 A8 5C 22 0E 7F 05 5B
 E4 28 AA 5A 29 56 E5 80 C6 05 5C 7B AB 40 F8 E8
 63 81 51 B6 A7 0D EE 9B B8 E9 6A 92 8A 96 BB 5C
 41 05 55 2C 4D 0D 96 89 DC B4 E5 17 DF 8D 95 40
 41 C0 FC 07 C1 70 82 17 91 B6 F7 22 09 35 17 2A
 C2 71 CE EE 66 21 59 B6 AA D5 A8 AE AC 4D 35 DF
 7A FC B3 AA 92 39 5E 70 BD E7 82 5F E7 19 15 06
 84 28 FB EC 43 42 76 12 23 48 C1 5B 39 D2 DF AF
 2D 60 C3 33 B0 11 5A 65 94 EB DE 47 6F AE 75 06
 64 D2 20 08 FE 78 E9 8F 21 AE 91 34 F9 90 3F 9F
 33 30 D7 3A C5 DD 41 EE 08 6A 92 A7 1F F1 ED AE
 57 44 9A E5 D3 43 CA 2C 63 21 61 46 E6 CD 97 D5
 C3 AB 74 B3 34 32 0B 17 8C 6F 30 CB 02 D0 50 99
 BB C3 38 8D 3E BE CD 8A F9 26 BD C4 7D A4 C7 2C
 C6 20 3A 3C 2E 4D 2E 06 2A FC 27 87 92 6B 07 FF
 58 42 2A FB 57 1F 9D 51 7F 3D 7E A6 D6 42 F8 C1
 F2 BC 96 1F 28 68 51 58 26 8F 1C FA 3A B6 98 A9
 64 5F 4A 61 48 6D 2B 20 2A 53 57 E5 28 07 B8 3D
 E6 F1 1F 90 64 6C CB 9C D0 69 8D AD B3 89 54 B8
 1F 14 1F 18 B1 6E 84 BA AE 80 F0 7B 65 A2 4A 75
 D6 F7 7D 55 0A 33 A9 CF EA C6 C4 72 9D 93 AA 7A
 B1 75 11 BD 83 5D AF 3B 3C 3B 5C D8 7E 89 C1 F4
 C8 04 60 EA 05 10 7C 8A 39 C3 46 08 58 47 79 7B
 06 4A 96 6F 68 07 FE 84 1B A6 0E 5C 51 7E 9B C7
 69 2B 96 36 15 08 BE 0A 8E 60 4F 00 BD 21 C5 EF
 20 02 0B FE 12 09 97 2E 15 8E B9 2D 74 D0 67 EB
 2C 4B 7A 3E 1C C5 6F 61 58 A9 45 F1 9E 48 86 44
 22 7E 3C 18 2F 8E 8A 72 31 6F B4 0E 01 4E 69 DB
 6B 8E 91 C2 E0 4F 79 AC 4D 35 94 52 7E 90 92 AF
 66 34 A1 00 67 2B 00 A5 04 61 0D BD B6 DE 4F 9E
 52 B2 0E F9 01 8E 77 7F F4 8C 2B 13 54 6D 6E 56
 38 6C 9A 86 B2 AD 7D B3 5D 3F C9 4D 66 1B 68 24
 6E 98 0D E4 7E 5D 48 5C 28 5E 66 06 30 42 85 24
 C7 DB A0 97 34 8A 7A 7C 0C 1F 6C DC FC 08 09 6E
 E0 EA 0B 59 B2 E4 82 26 40 D7 39 0E 46 FC 30 27
 BB 26 49 E2 67 C4 24 A8 AC 42 E8 23 96 A6 13 63
 75 4B 7E BC 98 7E 2D 40 61 0B 5E 3C 0C BC 46 FF
 0F F6 40 4E 0F 53 D7 CC 05 74 FD 85 E0 6F 59 D8
 BA CC 5D 80 FC 38 06 40 5C 29 00 55 1A 07 24 54
 23 11 62 0E 35 D1 BE D5 11 BE 91 30 20 09 77 78
 91 4F 9D 3A C4 40 C8 38 20 F9 59 7B D5 91 07 26
 A5 E5 12 78 C4 0B 1F F5 F7 AE 6C 56 52 16 0E B8
 D8 F2 29 09 09 08 1F C5 A0 D4 1F 3D 5B 84 F8 72
 5A 58 3F 47 13 7B FD 2B BE BD 5B 87 80 1D 66 97
 93 25 08 CB 70 19 0D 70 89 43 BE 69 45 41 63 09
 AE 8F 5A 11 0A 75 C1 01 FC CD 28 7E 81 BE 00 73
 09 BF 15 D0 70 FB 47 83 BE 5A E0 9A 3C BE 84 2C
 5A 79 44 94 E7 53 60 D5 41 20 63 E1 21 03 AC D0
 39 8C 79 E2 42 98 C4 9D AD 8B B4 6B 74 27 66 C9
 7C CF D1 C1 E0 E5 47 85 9A 05 99 D2 FD 3E 48 35
 74 CB C8 19 F7 0D 63 0B E9 41 77 48 F3 AE E8 A6
 8F 68 24 6D 54 AA B1 44 74 AC 9B BA 32 37 6A 0A
 D2 8B 66 CD 93 4D 2D E4 65 63 64 0E 8F 16 D8 68
 D9 9F F4 81 F0 E1 59 8A 03 5A 35 49 C5 F9 47 48
 51 3F AB 61 DD 0A 55 1E 78 58 41 B0 1A 1E DC C8
 44 4F DF AC 04 0B 0A 1C 0F 86 76 0B 28 D2 B8 D9
 6D 8C 17 3E B3 E9 50 B5 AB 18 B9 F3 2C 29 AC CC
 65 BC 98 2A B5 90 BA D2 63 34 8D F7 3B 7E F4 6A
 D6 49 78 D7 B2 50 D8 F4 3E 83 AD 1E 32 FD DD A8
 B1 ED 7E 9A 07 32 15 6D 86 66 FE F0 C0 D1 77 FD
 7B A9 F9 50 BA 7A 50 E4 3B F6 1E 29 11 DC F5 0B
 01 73 B2 32 00 E7 11 B6 54 DF A9 82 31 F7 4D 98
 AA 29 A5 9C FE 52 71 9A 4D 10 DB 19 3A 89 5C 11
 DA 97 2E C8 63 84 AF 7B 7A 86 EF 97 15 71 8E 28
 6E 10 EB 07 D2 C2 96 EC 5C 18 BC AD 17 C7 E9 2D
 FA 04 E0 A1 66 C2 4A 1D 18 8B A3 39 49 08 E6 9E
 4B 04 A0 DF 50 F2 42 FE 9F 7A C1 F2 2B CC B5 12
 9A 85 70 F6 B8 F6 D2 18 C2 AE BF 06 36 A3 9A C9
 45 4A BA FC 69 C5 0E D3 F0 AA 94 FB 3F A1 87 FC
 F5 C0 C8 C3 3B 03 37 B4 21 42 C4 1E EC 70 22 F4
 3E 85 8B 4E DC A3 07 AD E0 29 28 25 EC 31 CA 3A
 17 0E 03 4A 2B 09 38 11 26 E0 B5 1D 27 39 BA C3
 30 21 6F B6 37 DD 2B 97 5B 24 42 0C 2A 29 E2 83
 A3 8E 45 C9 9D 2F E0 78 E4 14 20 BF 88 A3 FF 70
 26 96 46 32 50 76 3D DF 71 64 EA 4B 55 E8 26 E8
 E1 4F 20 25 73 14 3D 33 12 0B 98 93 35 F6 14 90
 B1 95 40 A7 ED B9 CC C4 D3 97 26 56 FB 79 31 76
 D3 35 97 A0 E6 29 F9 68 A7 B5 36 FE 65 AC 60 EE
 65 BA 72 51 DA 29 10 1E 4E 55 82 2F CF 3F 6E 3F
 F5 1C 9E 5C 3F 7F A1 E6 E5 C5 CA 08 E4 82 D1 8F
 E0 77 F0 C6 C5 45 69 9A 17 92 74 80 3C F1 18 1B
 3B 72 5B 61 6C 1D 3C 58 37 BA 9E 5C B9 63 C8 BB
 C2 49 EA F0 37 64 27 E9 A9 11 6A 7B 5F 4D C0 08
 AE DC 58 DA 63 79 26 8D 64 FD 41 0D 2C 5C B6 7C
 67 BB 40 54 62 7B CF D3 8E CB B1 8B 2B DF FF 81
 22 A6 0F 3E 11 F4 26 85 85 3F 4E D0 E4 81 53 63
 DD 3F F0 DB 56 A6 AE 30 AC 8C A7 8B 89 2C AB D6
 60 AA C7 85 E7 1A 2A E4 04 93 9F 99 4B 3F 6B 9C
 01 CD 0A 60 60 37 AD 45 83 A7 8F 78 6A F2 25 95
 8A FF FD 25 37 1C 74 61 26 3A 45 70 C1 4E DC 2E
 C5 C8 CD 71 50 99 2E 8B 23 4B B8 54 F8 58 8C 5C
 4C 18 E7 E9 6A 65 80 B4 5B D1 56 20 14 F5 81 E1
 20 C7 28 91 FB 25 D2 01 2F 6A 0A 4F 0A 4B 26 EF
 F9 5A 77 04 5B 71 7D 2B 91 CF 29 CD 3A 77 CC 98
 76 D1 95 BD 1B CE 40 36 85 2E A1 7B A2 59 41 3C
 58 5E 9B 9C F8 71 E5 D7 09 96 E1 AB 28 1E 94 3A
 E0 D4 DE 4D 08 06 EC 29 E0 E1 C7 5D AC 73 CF 78
 44 AA FF 68 0B D1 F6 18 3C 42 70 51 5C 27 B8 BF
 55 13 07 B4 8A 5C B1 B5 1B 8B 63 6D F9 F9 37 B5
 80 67 DC 60 AF 8B 93 8C FA 30 CE 31 B4 7F 1C E5
 FD 54 8D 70 AF 0D E2 E5 A6 E5 71 14 D0 E3 38 8A
 A1 F8 EE FD 2B 46 72 25 EE 3D F3 80 A2 1E 2B 53
 A3 5E 95 4C 9E F6 3B 72 85 D4 AA 04 FA 3E 4E C2
 A7 B8 3D CC 75 8F CA FD 31 DA EF 38 4B AA 68 BE
 71 50 0B F7 4C 72 6F 6A 1D 8C 9F F9 A9 D5 D4 E4
 43 03 5C DC 54 9A C3 4D 49 24 70 48 15 53 18 2C
 08 A1 76 6E B5 C1 99 F8 16 77 0E 84 CC F7 02 4D
 54 6B BC 43 E9 1F ED 9C 0B D2 B5 C8 3C 02 27 B5
 5F 4E 81 87 82 A7 E5 6F 11 49 1B 62 59 3D 5C 19
 E1 69 E0 7D 65 18 A6 0B 6F 67 CE 8E 9B 0E DE 7B
 0E B7 51 89 64 A4 76 71 65 F5 83 7F 4E 91 40 E5
 9D 51 B0 F4 0B A8 07 AB 69 7D 3E 32 CF C5 0E 06
 B8 13 1B 89 42 F3 6A DE AC BE 77 67 94 FD 73 5B
 71 0A 52 8C 6A F2 6C 5A 35 99 90 40 5A A2 6F A1
 12 22 09 C5 1B E9 E5 7A 0E 39 4E E3 25 CD F7 FB
 BB A8 84 83 A3 EC 01 8D 8B 1D 01 E4 95 81 B9 28
 45 9C C4 43 89 07 CE 49 57 6C F3 F6 8F 61 C8 3C
 99 40 BF E6 07 72 B7 0F 68 82 FB 6E 1B AE 60 47
 29 1D 84 40 35 3E 80 ED B0 8A F9 13 C3 D2 78 25
 1A 67 66 1F 33 02 04 FB 9E 29 FE 9F C3 FA 1E 78
 71 3E 5E 91 39 DD 56 78 A4 6E 50 7B 09 FB 6B E9
 F7 28 D3 AD D7 50 FF 7C F0 A1 6C FB AC B8 C5 7D
 00 C9 A7 51 4D 36 56 F9 64 0E E1 7A AA 6B 7B 16
 C5 A3 25 F5 18 BA 3A 88 68 6B 23 9C 35 DD B2 65
 CF 9E A2 B9 6B 4E 84 46 67 D3 FC 90 1A 58 23 1F
 CE A7 93 7F A2 6D 08 CA 29 A3 5E 54 9F A8 D2 61
 E5 C5 FA 5E 8C 20 2C 63 51 C8 72 13 4A 7C 88 C2
 82 63 AE 84 DF 8A BA E9 9F B3 C9 EB CB A8 59 6B
 2E 32 13 D4 E0 76 3C 3E EB 19 53 31 D3 C8 50 52
 9E 70 D9 CD 69 FD F4 1B 42 E0 81 92 75 ED B1 21
 DA 4F C2 CE 04 11 A7 AB 4B 4E 58 F4 5F 01 17 9B
 6B A8 03 12 2A 10 67 89 0F 1F CE C1 2C 21 F0 21
 05 19 ED 1E 2C 00 4B 3C 3B 63 A8 BB E3 D9 2D 4C
 31 C1 74 E0 F9 D8 45 63 EB 0D FF 05 1F B9 F0 21
 2B 5C FC D6 50 51 C3 37 36 4F 60 A4 54 BA E8 CE
 3E C8 3B 55 3D AB 1E 43 E2 CD F2 4E C3 25 A5 C7
 72 29 13 96 79 71 19 1C 07 2B FD F3 CC E2 D0 86
 3F C7 E3 7C BA 58 25 EA F0 F7 3A 45 FB 2E 45 13
 BD B8 EA 7A CB BC 86 86 4A CC 43 CA 12 75 9F 34
 BC E7 6B A3 3E 44 93 C4 AB EE DB 48 4F D5 7D 9E
 48 0B 46 C4 0F 96 42 D0 10 39 C1 A3 FC C4 37 61
 C5 67 0E D4 3C 6F 47 A3 C5 0B B8 6D C7 B5 C3 8F
 C0 09 5F B8 EF 9B 92 7F 1A 7A 9F 8A C0 F0 99 46
 A0 B4 CD AA 59 56 70 D9 7F 28 A1 49 04 EF C5 E3
 91 76 68 18 F6 C6 B9 10 12 36 BB 45 E8 CC 94 D5
 F4 1D DF 42 61 71 4A 9C 0C 25 91 17 6E 84 91 7B
 71 C9 73 0A 18 F5 1C 80 C0 57 09 EB 77 FB 75 EF
 27 BB BB C2 0A C9 42 3B F8 F6 0C 87 7E DE DA FB
 F9 D7 3C 96 C1 18 E9 91 A4 4C 9D EF DA A8 20 5B
 DD 06 A1 8D 80 D8 C8 F9 C0 21 87 AB 9A 88 8D 6D
 7D 92 1E 21 E6 78 46 C0 FD B1 89 5D 04 FF 0E 6D
 4B B2 F1 A6 5C FD 88 3D 72 67 B2 D3 77 7B 59 FE
 82 5F 5A AD 28 26 16 29 5F 73 5A C5 FD 82 FC B6
 49 4B F2 7C 0C 52 B2 5C 66 3B D0 41 4D 21 14 EB
 A4 A4 00 02 10 D5 CD EB FF D3 87 B4 81 FC 31 DD
 B2 9F 9C AC 7F 09 77 E6 8B 23 BD 5A 40 A0 2C DC
 BB 38 52 C9 35 41 E8 12 0E 3E 45 90 00 C7 5C CE
 11 25 26 1F E4 A2 19 4B 36 E4 D0 EC 76 35 F2 94
 FA CD 70 F6 EE CF 01 46 CC 09 2A 89 99 D0 56 CB
 A9 A5 FD 02 99 48 C8 C9 A1 C3 19 07 FB 10 AB CD
 FA 99 17 A2 E5 07 F0 6A 93 AE 7D 73 C7 40 06 A8
 00 F3 67 99 D6 EE F7 BF 43 9A C7 72 50 71 D4 32
 8D 77 D6 CF 35 AB 8E 90 67 EE A9 4D F2 D2 9C A3
 3B D0 EA 95 15 CD 7F 6D 3F 4B 55 98 8B 9C 91 E0
 8D 7B 0C 98 32 DA 41 59 07 28 69 05 A7 BA 5A 9F
 A6 9F 43 FC 9F DB 54 07 D5 D1 6A E9 A7 17 14 E2
 14 33 69 53 CF C9 F3 3B 4F 82 DB 36 F3 34 DD A4
 B2 82 CE 61 18 2C 8A E5 ED 8E 00 B5 A6 49 7F 7A
 28 1E E0 3E 13 2F 71 77 A1 2B 46 69 73 2B BF 44
 41 A7 D0 2D D2 DF 03 61 1D 9D D6 AD F6 1B 6D 91
 3A 52 67 55 73 D4 72 3F B9 17 40 B4 3F C0 32 13
 62 A6 B4 40 95 29 A3 56 A8 26 E3 74 8A DC D6 18
 D7 76 13 98 89 38 85 82 D3 18 57 8E 6D 72 59 74
 A3 ED 55 FE A4 82 C8 3E D6 90 DF 0B 0B 43 38 BD
 80 B2 1E EC 04 02 B3 1D 91 04 F0 93 E8 3D FD A5
 AB EB 0C 50 F2 82 79 EA 0F 52 5B 8B 49 A8 56 F7
 E5 75 43 BA 2B A3 D4 80 B8 78 7A 66 D7 F5 AC F0
 8D 90 1C 19 DC C0 9D 15 18 0E 46 2E C2 9F B7 0E
 9D 40 37 A6 2C 32 BF CE 2B CE 2A 66 EF 6C 8C 6B
 65 01 2B 3B 4B BD 2B 58 5D F0 FB FC 44 F8 73 F8
 8D 53 89 4A 75 7A E1 FA 4F 38 79 C0 65 E1 C5 52
 CE 9E 3D CA 7A 65 C0 B8 94 28 EC 8B 4C B9 A2 4C
 7A C1 4F AA 20 93 39 11 95 60 08 AA 25 19 4B E5
 32 30 E8 E5 84 BC 62 FB DD D7 1D 57 D8 03 67 92
 8E 2B 2A 43 1E 2F 7A F6 AE B7 C8 70 2C 15 4E A7
 22 BB 8C 2C 13 F0 88 F6 58 E0 FB CB 75 F1 6A 37
 32 05 28 ED D4 05 3E DA 48 4E CB CB C8 32 FC 20
 AF 3B DC 75 96 97 F8 6B 4E D8 61 BE 6B D4 D5 17
 3D F5 55 37 F1 DD 95 11 97 AA 09 59 20 8F 6C A4
 48 13 01 3B AE 60 A5 02 41 05 47 B0 F7 D7 19 7A
 6E 0F 8F 6E 18 29 4E F2 52 24 AB D9 C6 9A 4D 1F
 48 03 8B BB 79 A0 DA 99 9D EB F0 6F B9 55 DA 91
 CB 80 2C 8F 87 4C B6 C5 C0 7A D0 45 39 FD 71 32
 33 A0 56 F3 38 D5 37 4E 9E B4 6D BC 7E 88 5F 85
 33 61 3A E5 D1 09 ED 1E 41 B6 83 6E C8 94 2D 80
 C9 64 54 5A B3 4E EB D6 04 54 38 7F 38 72 8B 99
 84 05 ED 75 13 D6 AF D6 89 CA 2C 21 D5 54 81 BC
 F3 AF B3 B0 06 11 8A 69 24 4B 04 0F A1 83 77 F3
 C4 00 CD 48 B7 BC D0 02 A9 67 C4 45 D6 6F 23 36
 80 66 1A C1 76 26 9B C4 CF 8B F8 28 FA 5A 2C 9F
 DB 4B D7 2F FC 86 C6 08 66 65 0A F1 F0 1F 0B 89
 22 C5 47 60 13 14 CA 16 19 78 CF 7D D6 26 33 95
 3D B7 98 8B 61 F2 83 3B AF C7 F4 D4 C3 80 26 1A
 CD 26 5C A2 21 15 BB AD 5C 8C 8F 2C 81 54 F2 E2
 FC 06 36 3C D3 06 D7 E7 A1 4B 1D C1 98 B3 74 F5
 A8 81 D2 64 DB D4 99 54 CB 5E 8E C6 44 69 94 D8
 A3 D2 EF 5B AD F7 CF E8 16 23 88 3E 3C 79 0A 55
 3F 2E 7D 82 06 98 FE 00 30 F0 6E A4 55 1C 7A 64
 7E EB 37 D2 B2 51 C7 F9 39 84 4E 4B 80 97 E0 6B
 63 54 F3 08 F9 D5 77 D0 B6 38 8E 88 FD FD 50 96
 5D 9A E7 C8 3C 6B 21 57 2A 7E E8 5A 4E 9F 3A A8
 D7 46 87 C4 D9 A0 97 26 5F 66 FA 4F C4 77 7A 62
 9D C8 55 92 CD 52 79 E0 56 75 12 0B 4F 8B 56 86
 BB D3 16 24 8B C4 33 30 F0 3A FF 99 10 9E F6 0D
 47 97 8C 93 D8 B4 07 0D F0 E7 99 DF F7 48 50 D5
 6B C7 44 7E 00 2B 19 D2 D7 FF F6 D2 66 A6 6D 97
 BA 86 98 4D 44 11 81 44 21 F1 16 04 F4 95 BE D5
 56 81 E1 81 F7 DB B8 5A DA B6 15 62 FA 22 A2 15
 A7 D7 EA 35 8C DE B4 33 D7 F7 D2 FA 3E 3C 98 17
 C8 8A 2B 11 93 A0 7D 92 E1 9D AB 53 87 8E 45 46
 0B 58 D7 BE B5 54 7F 92 2D CE 8F 0D C5 F3 0C 1B
 0A 0B 53 8F F6 C3 70 36 65 B2 FB E2 E7 DE F8 64
 5A A7 A9 C6 40 40 F3 6A 2D 8A EC 1D 48 79 0B 4A
 D8 33 74 07 BC 10 D2 D5 8D 71 77 55 2A B8 1B 6E
 EF 8D 61 FF 0F CE 8D 36 C4 F6 62 2C DA 17 F4 0E
 7E 05 28 82 86 36 A6 3B 0E E6 B4 25 DC 05 BF 9B
 8D DE 46 A0 AA CF 5B 90 E4 76 42 B9 0E FE 81 2D
 6F E5 D6 7D 3F 90 FC 1D 89 9F 7D E1 4B 96 F1 44
 66 0A 48 6D D2 54 67 E5 DF A3 4E 42 DD 2B 1B 1E
 7C 71 88 98 D2 35 12 6F 0A DE 78 90 40 EB 7C 06
 32 AE 8A B2 A3 53 7B 39 A5 DC 53 37 E3 7A EE 8C
 4B 6A 85 0E E7 47 9C 4A A8 23 4A DF 2E 20 52 2A
 F6 84 B1 E2 F0 7C FB 39 23 C5 71 69 CF D9 E7 6D
 11 59 7E 63 F6 F0 51 D6 C3 BE C3 6D 6A 2E ED 3C
 85 43 7B 9D 5E CE 08 42 2A 74 3B CF 0A CB 3E A2
 AD 24 95 3E 3E 01 98 89 49 5A 47 7E 02 C2 AF 64
 71 99 C6 23 B5 D8 31 3A 81 86 53 CB FD E3 A3 FE
 4F 25 F6 A7 64 9D 76 A5 F8 A5 23 FD 9E A0 D0 D0
 C9 E3 7F A3 84 42 F4 41 A1 7D 94 06 AE ED CD 91
 85 A9 2E CB 07 C5 0F 65 D4 FE FB 60 F8 3F 63 95
 B2 44 3E 4E 8F C7 7E BB 50 6A FB 31 75 B9 F4 01
 CB 43 91 34 92 53 24 9A B5 66 93 46 49 33 E4 5C
 C0 9E 4A 04 29 71 1A 57 0F 82 AA AF E2 4C 95 DE
 6F D2 BA FB EE AD CA 50 1A 5B DC 8B B6 FC 2B 93
 77 11 C9 CE 15 DE C0 93 FC 63 05 53 F5 FF AE 68
 F9 45 78 2B 56 8F 39 74 ED 8E 36 BC C4 23 A0 90
 25 0A 11 8F 33 E9 D3 67 56 77 57 6A E6 48 C0 A2
 4F 98 58 CE 32 0E D8 53 AA 7E B4 53 A9 60 AA 68
 A4 E8 70 45 C3 FF 60 28 6D C9 F3 CD E2 36 55 D3
 43 F6 BE 34 AF DB 39 1D F4 F0 14 61 44 54 D5 CA
 12 97 E0 03 9F DF 4D 89 A2 26 47 BF AA B2 FB FD
 18 A6 2E 3B 13 61 E6 2F 88 D1 EA 73 6A 4A A3 AB
 39 71 49 1F 51 CA F9 36 DC D6 C4 39 2D A8 40 ED
 DB F0 6C 1A B2 DE 46 71 98 F6 1B 37 77 B1 FB 4C
 DD 08 47 A6 33 00 AE B5 89 30 24 14 8D 12 AD A8
 80 5D 86 EE 79 FC 99 9B 28 C9 21 F9 24 43 DF 95
 51 53 8C 88 83 0C 45 AE E2 68 63 67 FF 41 8B 4C
 0D 1B AD 9C 49 7C B1 2A 0B 82 89 ED 42 38 F8 0E
 4E A0 6A 96 9F 7F 2F F0 6A 27 3E 28 3D DC 68 37
 1B EC 1D 36 5F AD A2 E5 6B C1 0D 82 64 67 40 49
 52 A7 5F 94 81 10 F4 46 12 55 1D B7 18 16 69 89
 BC BE B5 69 71 B5 47 CD C9 1A 82 0D 7F 24 13 6E
 0C 31 23 63 78 99 D2 94 25 C6 F2 AD 52 AE 39 40
 75 4D 37 71 3B FE 9B C8 C8 EC 00 13 D0 EB 64 6A
 B7 58 FC 35 57 80 4B 6C 58 A6 B4 FB 75 38 AC FD
 CE 50 E5 5E 9E 16 BB B7 F5 64 B0 B6 D0 63 FE 0E
 DF 23 3E C1 07 BB 99 EC A4 6E 50 B2 1B CF 2C 94
 79 5D 74 80 A5 6E 2C B1 1F 7F 77 11 68 15 51 C8
 F1 C9 13 11 41 73 74 0A E7 22 EF C8 DC AE 63 37
 7A 56 87 A4 0F 04 7A 1D 88 D2 10 4E A9 13 28 8C
 AC FB FE 64 B4 52 C0 BC 64 68 BB 05 B7 89 07 76
 36 6C 82 CF 31 E0 57 75 98 B1 54 6A B8 1E 7B CE
 57 55 0B 7E F7 4A 52 3D 21 2B 28 6F AC 7D 88 98
 4D 48 47 51 1D 51 B0 93 7D A1 79 5B 09 76 64 5D
 BC DC 0E E8 0B 2E ED 1B FC 35 36 4E A3 04 83 AB
 ED 95 95 8B 7D 0A 2D 3C 2B F1 BE 93 F4 3A 25 81
 7C A8 62 51 FC 00 55 E3 5C 63 4D 89 1C 6C F5 EB
 14 16 EF E7 A3 C2 07 FF 56 ED A6 F8 70 6E 91 AF
 FB EA 98 9C A4 5B 5A E9 84 FA 2B A6 28 48 29 73
 C1 65 09 E5 88 9C 0D 25 5E 33 FD 6D 1F 59 4F 59
 99 11 F1 88 2C 3E 0E C7 17 D1 29 03 C8 97 D8 81
 9C 50 35 1C 70 75 36 FF BA 77 D4 02 29 8F E5 B1
 64 6E 1B D9 38 CE BB 06 37 03 16 C2 D5 D9 EE 92
 5F EB 98 C6 94 BE 21 30 46 95 B4 B8 E1 E7 02 CC
 59 8D DB 61 D1 9A CB 93 2B 31 A8 A4 FC 32 68 2F
 B7 B8 F1 92 CC 42 76 21 9E 28 E6 48 F3 A1 EA FA
 1D F9 F4 D8 0B 5E 33 25 49 75 E0 48 ED DC 3B 4C
 6B 0B AD 7A 33 16 A0 EC A4 0E 4E 2E 2D 60 F1 CF
 33 5E 03 F4 B1 78 F0 B8 42 75 33 87 77 4F 50 F6
 C4 24 F1 60 5E 9B 65 76 37 13 E9 3E C7 48 0A 9B
 46 2A 0F C0 66 BC 74 67 2A 9F 78 D6 A5 18 C1 AA
 46 07 D0 D7 73 95 81 84 6F 4A 72 62 8F 4E 49 3E
 D1 62 7D E9 43 DC 86 48 D8 E5 C6 24 D3 95 40 98
 07 2F D6 BC E4 26 C4 58 5A E1 30 B2 A0 1C 89 DA
 5C 15 A4 B4 18 38 EB 68 FA 6D DE CE 3E 6D F3 AB
 5D AB AC 50 A2 35 04 6F D2 1B F0 0B 7C 07 0C EF
 02 F4 CA 87 0C AF DC 72 21 D2 98 5F 2A 52 BF 6E
 50 E3 BC 81 64 50 A1 71 80 4A 38 BF 7B E4 C0 8D
 9F 93 56 48 47 7F 54 83 22 C5 8A 01 80 B1 10 C5
 1E 4B 98 8C 07 63 4C 9F 6E 4F 5A 66 65 44 B4 92
 EC 32 34 75 3B A6 5B B9 E8 42 8B A0 97 BF 68 9D
 F3 39 95 ED 91 60 83 74 96 0B 40 C5 BC 99 97 45
 29 18 C5 67 04 73 35 2F 1E BE 16 DA AC E9 7E 68
 00 EA 95 8C 83 C8 D0 1B 52 45 61 52 D6 29 86 25
 D6 E2 1E F7 83 75 29 BD A6 1D 46 6D 28 79 3E 00
 0A E0 DA 74 F1 FA C2 D3 65 49 77 DF E9 38 18 AA
 52 C2 7E A0 F1 7B 75 FE 4F B8 BB 4A 49 8F 18 BB
 06 F7 41 D8 19 B1 58 87 D1 C2 C5 15 68 B4 8A CC
 7C 9E 54 DB 0F 83 B5 DB EF 8F 1A E7 3B 8A 74 7C
 BB 66 FA DF BE 0C BC C1 9E 7F 21 E2 8B 3D 25 19
 3E FD F2 66 4A 4A CF 3C D2 A8 74 14 DA B9 C3 2B
 2D 03 FA 18 07 A0 E8 A8 89 BF 65 22 49 C4 96 9E
 B9 C3 0E C9 5E 09 7B 2E DF A6 7A 8A 57 D7 D9 98
 36 6C 7D 6D 9D 59 9D 16 A8 6F AD 0E 57 A5 27 CB
 24 FF C2 E4 58 30 E3 FD 0F 01 71 6C A4 97 91 63
 23 FC 44 3A 44 BE 60 AD 05 59 6A 38 F4 D6 CB A2
 E2 C3 9E 83 89 27 9C 9F 62 21 58 FA 25 AD 48 21
 87 FB 42 76 95 85 1C 09 E2 52 97 4F E6 23 39 BD
 8A F4 6B 83 F5 70 95 E4 2F 57 0A 9C 9F BA 37 13
 DD CD 56 BC 82 EC 60 9F 0A 65 AD 7E 1C 70 2B 5D
 41 2F 8E 9B 22 87 B7 25 A6 D4 33 CE 07 5C 46 C8
 00 AE F9 D7 C5 37 E6 CA A5 9F 0B DB 12 E9 99 86
 D8 1A 7B B7 1D B5 6B A6 D7 9C CF C2 06 FD 74 9F
 17 0C 28 C1 96 92 94 F5 A6 22 8B 9F F6 32 70 99
 C8 8C D8 F1 BF 94 AB E5 DD B6 34 B6 AF 11 73 E7
 60 F9 E3 C5 6F 6A 83 A9 A7 14 D8 AF 68 8B 7A 37
 97 61 FF 61 72 87 17 C1 67 B5 97 C7 68 7B 52 FB
 FD 8B AC 1C 15 FC F4 1B 1A D3 A2 60 FA 23 F9 BB
 5D 39 E7 AE F3 D3 6C 5B A6 4D 51 75 18 7C E8 18
 24 8B A4 C3 B3 49 EA F1 2E D7 D3 E4 BE 02 49 C8
 EB 7F 1B B1 59 90 28 1B 29 A4 F1 E8 73 F9 E3 B4
 DE A8 4D 33 A7 8F A7 31 5F EF 5E 18 0B B6 7A F6
 90 6C 66 D6 85 9B 39 CC EC 67 D5 90 ED 81 B9 72
 17 AD 9B 5D 12 33 6E EF 06 96 83 22 66 67 CE BE
 0B 8A 47 2D 13 92 62 48 17 35 2E FD 83 E5 91 8C
 ED 4A 4C 04 35 37 9F CD A5 DD C9 74 FD 26 4C 70
 DA BB D9 8B 56 BE DF 2D 48 2B 8D B1 96 D7 87 45
 89 3D FD 51 B4 0A 45 00 63 7F 52 95 D3 8B 22 FF
 62 05 CF 40 0E 62 23 DC D6 09 61 8F 42 73 0D 73
 A2 6C EA F0 A9 69 A0 9C 9E CE C5 83 53 BA 0A 89
 6D 33 82 5E 34 78 C9 E1 48 0B 2B 2A 2D 6A BC E5
 FA 48 28 27 9C 1B E4 0E B0 E4 05 C1 71 AF A1 02
 CC 73 2F 93 9E A0 D4 A4 D7 93 16 A9 C4 FE DB 51
 15 49 8D AD 25 D9 AB FD E2 55 06 7A 7C 26 AA B6
 A0 E8 5E 21 DE 34 94 75 3B 20 28 C6 54 80 13 89
 26 A8 3F 8F 57 F4 F6 EB 2C D5 69 4C A2 B3 C7 41
 95 4A 8C CB 3D 3B 95 FC 63 B4 2A B0 0A B4 0C FD
 37 67 60 44 3B 69 73 66 6F 36 F7 63 58 84 90 AC
 BF E9 42 5B 79 CF 51 04 70 79 33 F7 ED D1 96 20
 07 40 CA 68 A4 C3 8D 28 8E BD 92 AF 1C 1E A1 BD
 85 68 E5 B8 65 FB 96 C7 76 3F 92 26 78 40 0F C7
 A8 9D 85 4B 29 C3 71 9F 23 E8 70 5B CC ED F2 45
 D0 8C 6C 34 92 A9 5B 18 E1 4F 90 DD B5 0D 80 BD
 9A 5A 61 A6 30 66 6E 14 02 DD 88 77 8C 0B 82 98
 A5 5B B5 97 8C 10 BC 14 8C 0B A7 46 0D 93 7A 36
 D0 33 FC BB 49 7C 1D 35 0E C5 11 FB C3 9B E4 CD
 AB 60 AB 69 6E 64 88 63 92 D7 CA CC EA 87 BC E8
 56 16 09 D9 54 A5 B5 1E 59 06 76 EA CB C1 EE B5
 3C EE 38 5D EF 8B AF 75 B5 1C DD F6 90 EF 02 63
 4A 15 12 A3 33 2D BF AB 62 7D 8D 54 3C 5F D8 A2
 17 02 18 27 72 35 79 3F A6 E8 D9 61 B6 71 21 2A
 98 C1 CC 24 DA D4 D3 6D 6B B6 FA 70 A5 56 E0 A5
 C7 D5 EE C2 EC E6 F7 FA 43 38 DB BF 64 4B 29 E3
 A2 FA F9 19 D6 AE 22 06 AB 2E 07 2E 9F 25 F2 E1
 FF 16 9D 17 8F A7 84 D0 15 B7 7B 3B E5 3B 13 2E
 E4 2C 58 58 C2 60 27 6B 95 B2 3D 21 AF B0 66 FC
 96 47 63 FC 85 6C 0B 91 5F 18 16 C6 7B EC 63 5E
 6A 13 AC 60 20 0C 90 08 4D BE FB 9B 7F 30 3F 9C
 5E 50 93 A6 F1 A2 1F D5 D5 B2 22 FE B4 51 EE E9
 A3 D8 D2 EB 35 0B 1D 2B 6D 8B D4 A6 06 E5 2A A2
 54 54 11 4B E2 D1 04 B6 76 2E 38 73 19 7F F2 B4
 7B 3D A6 48 33 A8 BC 04 5B FE DD 1B 1D A1 93 D9
 50 FE 11 93 B3 C5 28 0F 2B FA 5C 7D 6D E9 AB F6
 F4 F4 91 57 EC 50 96 83 72 50 BF A7 47 8F E0 D2
 A6 E4 40 77 21 9D FC D0 F9 71 30 BC 40 86 25 92
 DE 14 BD D1 02 19 01 9D 16 87 00 68 C3 11 BA D4
 9C 33 93 CE A4 CA 49 5D 7E 4B BE F5 C6 EF 29 74
 A3 C5 7B 27 1B 2F 9C 24 81 E7 35 06 FA 30 12 A0
 29 E5 19 E2 5F 34 58 3A 3C E2 AB AB 90 9F 60 09
 CE 14 2E 80 70 76 03 B3 2C 3C FE D8 A8 EC 82 57
 CE BD 7B DA 0E 01 00 59 A9 CF D1 9A 5B 59 56 F4
 D7 D4 AA FC F9 E6 33 9A 18 DB E0 E4 F2 83 14 02
 BD 5D 88 D7 3D 27 8A 1B 6F 04 43 57 30 DA E3 A6
 68 CA 31 45 85 B3 A9 81 30 E1 43 81 69 FD 69 E0
 2A 64 F1 B5 6C 16 20 10 02 DA BC EA A4 5A 97 81
 AC A3 69 59 95 C2 30 FE 4A 98 DD 71 C2 05 66 65
 67 48 3A 42 FB 70 42 37 E9 E8 60 F8 90 D4 28 7E
 E0 FA FF D8 4F EC EB 36 B3 70 EE A1 91 AB 82 7A
 EE 37 4E 1F 71 16 0C 93 2F 47 26 35 55 1D FD B2
 92 62 1D 33 81 F1 80 8D FA 92 FD 36 B8 D3 E2 A8
 FE 8B B9 B7 4A C7 5C CF 75 C2 83 AD A2 C2 CA D0
 E7 E4 16 6B 20 07 01 84 03 BC 60 70 64 0C A4 FB
 A5 06 67 CF DB DD 0F B1 E4 59 D1 C3 8A D6 DD 5A
 59 27 D5 8F D5 FB 61 3C B4 72 03 80 8D 2A 17 31
 2F 69 04 0F A5 37 F7 66 A4 E2 50 12 C9 B8 68 86
 5E BF 09 87 0E FC BB 95 0B 1C 25 9B E4 9F 7F D3
 57 75 2E BA 5F 2F 90 06 01 66 04 8A DE 12 2E E5
 ED F2 CC 1C 07 49 2F 8F 9B DF AE FC 97 09 F6 F9
 6D 8E B6 C4 72 E0 AB 47 5D E1 06 31 6E F9 E5 A4
 A2 0E 63 39 69 DD 1E 23 82 41 DA 40 34 CB 71 42
 20 8E D1 AB 7E 1C 75 53 CB E0 73 98 8F A5 63 73
 F3 95 40 D2 25 85 25 B3 2E 6E 85 8A F9 9F CA 1A
 D4 05 D7 97 ED 2E 74 C1 F4 C1 EA 1B 09 93 D6 E2
 4E 78 D9 74 05 2A B3 D4 95 84 3F C6 46 79 E1 88
 90 91 74 81 2D D0 0A 46 FE 6C 9C 04 0A 06 51 A7
 7D 8B 65 EC 5A A3 28 AB CA F0 5C 5E 30 CE B0 51
 16 BD 34 41 95 F5 84 37 6B E1 CB AF 87 74 13 7F
 F3 0E 43 E6 D4 2C 6C 71 E5 CF A7 31 45 CE A0 0C
 97 25 4E 35 CD 40 3B 25 9B 34 9B FC 98 4F 37 12
 F5 9D 69 C4 07 81 D6 38 92 1E 02 39 C5 DF 47 CE
 A2 5A 9F D1 BD 08 06 D3 91 A4 04 04 A2 D4 07 A6
 1B 05 50 A6 A0 A0 04 BE 7D AB BC 25 BE 43 FE 79
 0C 2A C7 AD 5B B1 1F FD DE EF 87 5C 62 1A 5F 53
 66 56 E4 E3 B5 E4 B9 38 94 B2 49 41 12 46 EF 9D
 D8 7E 6B 59 2C 44 2E 93 6E EA 9D 4E 6D 0A B6 8E
 F0 BF A1 E3 3F BB 4F C8 DA 4B B9 F3 A1 8A 5D 09
 4E 3C 2A F2 F3 D2 79 85 05 22 EA 32 FB B5 36 AB
 82 79 41 90 FC C1 80 3A 41 02 20 50 6D B2 E5 2C
 48 95 39 E0 6F 80 A6 64 3A 4A B2 E3 B1 91 42 1E
 6F BA 64 2F 9F 80 68 0F 5E 69 3E A0 3D AF 13 7C
 4D 16 99 07 07 28 EA 53 C1 B4 73 77 32 8F 83 72
 E5 FF 5A E8 B9 19 8E 79 6B BA F0 07 08 B0 E1 2C
 97 77 49 40 CE F6 57 5F A5 4A 04 DA 4A 03 2C 53
 3C EB D8 1C FE 5C 29 98 5B F6 9D E3 5F 1D 80 A5
 F9 19 3B F3 FB B7 6D CD 7F A7 F2 B1 EB ED 98 06
 BB F1 37 3A 7B E0 90 45 87 29 8C 0A 25 F2 16 BE
 83 A4 08 D2 8D 75 2C 70 3F 4B 68 62 0F BE 36 61
 09 E5 15 AB 49 FF 00 6C CF 9B 07 AF 54 E2 9A 72
 0D E6 B5 3A FB 19 AE F2 1B DC 9C F9 81 5D 4F FB
 7D F8 AB F1 D4 01 EE D4 E6 AE 08 D8 3E ED 69 DE
 60 63 12 95 46 D7 16 2F 49 04 4C 55 40 41 07 00
 60 63 76 0A D6 A7 86 02 95 F5 D2 41 49 DB E4 4B
 AD 26 9A A4 35 A3 B1 C7 35 72 43 05 28 D9 E4 91
 C1 A4 14 76 0B A6 86 A8 10 DF 8C 65 08 37 07 82
 3B 8D 19 8B 06 DE 36 70 B3 47 4A 2E BF 61 9B 3F
 15 58 D8 7F 68 E6 3B 53 E0 BE 66 31 70 70 3B A2
 73 48 4D FA 14 43 13 E3 EA 2B 79 24 39 E2 B0 45
 B1 A5 E3 CD 11 07 03 37 93 EB 56 DE 9A 68 7A A2
 90 F0 5B 23 2C 5E DE 94 AE B9 A2 F8 E5 D4 1C D2
 63 B1 3E FB A1 A5 00 AB 77 53 6C 24 51 3B 94 0D
 31 53 FB 37 29 62 0D 20 F9 EF 53 F5 28 E0 D2 89
 84 AA AB 48 D8 A4 71 CA 76 6F 0B 75 8A B7 4C 68
 68 34 82 DB 0B B1 4A 3B 16 01 A0 58 0B A0 82 F9
 03 A6 6D 74 CF A9 60 DF A1 2B CD 4E 04 ED 1F 69
 FE B2 31 E7 BE 15 44 7A 77 A0 5B 07 0F F3 45 B5
 D6 1B 3E ED CA 10 0B 5F CF EF CC 53 04 DA D2 6B
 5F 0F E7 1F 2B 03 90 5D 96 77 95 6A 1C 20 A0 8A
 ED FE 66 71 D1 34 75 26 16 3C 06 40 3F AB F6 9B
 69 A4 EF D6 83 7F 95 37 76 85 9E 37 AF 27 13 A6
 2A 7E FA 7A 15 9E E2 A8 81 3E B8 FA B5 31 56 5E
 32 0B 60 17 E1 B6 E4 8A C1 16 CC B4 DE 3C A3 7B
 CD 9D A6 C1 1A CB B2 FB 79 AF 85 E3 30 1D 0F 72
 D8 33 87 2B 8C AC C9 AC 57 89 4D 13 02 3B CD 43
 8F 36 B6 53 E1 12 04 68 FD FB 1A 7F 1A C6 7A F7
 86 B6 07 B0 79 CB FB 1D DA 76 8B C1 71 D5 53 68
 FB 23 50 C2 8B 70 86 DB 95 55 69 D3 83 35 C7 D2
 78 D8 7E 96 B8 BD 1D A8 59 92 FE 11 40 05 8F 47
 40 D7 C8 11 24 C0 19 55 9E AD 4F CF 8C BB A2 7B
 46 CA C5 63 5A 88 4B 88 FC D5 1A 5F 7D 97 96 45
 2F 50 83 57 41 20 10 35 F3 6D E8 88 90 02 BA C4
 30 4E FE 68 31 A1 EE 37 BE CB 97 A9 1D 34 38 57
 5C 8D 6F 72 16 E0 1D DD 89 0E 9E BB DC 7F 5C 01
 1A 01 D8 44 E3 F0 9F 8A C6 DC 67 AD EF CB 3F 61
 01 37 54 BA 16 B4 31 B2 E6 0A 4E 45 E7 1B 90 86
 22 06 8E FF F0 23 DF 68 0A 4C 50 E2 8C A3 F7 2E
 0B 4F 8F B6 ED 06 32 EF AA 8A 12 5A A4 F5 6F A0
 3B BB 21 40 86 A4 4A 81 B7 C0 07 DD C3 A7 24 0C
 D6 F6 AB 8D 68 59 58 8A BD 49 F9 EE 16 A6 D9 D2
 FC 49 D7 0C 79 49 B9 44 D1 45 42 60 A6 96 11 02
 4D 6B F1 D8 17 7E E8 E0 21 58 9E 3B 52 18 34 2B
 A9 D7 3B 12 75 F7 96 77 1D E2 34 46 42 7F 82 95
 45 C3 AB 6A 52 A1 4A 7D 88 52 AA 17 3B 47 04 D6
 77 4D C8 B6 C2 A9 FC B7 FE A6 62 04 2E B3 23 24
 08 12 6B DD E3 07 5D 00 A5 12 33 3D 28 40 DB 12
 E0 C5 E5 8F 72 07 01 57 F6 D5 1E B9 F7 14 AD A3
 42 D1 8A BD CF 3E D1 70 7E 12 4A AB 41 78 9B B0
 05 6E D4 22 AB 63 6E FB C0 4E 68 31 B9 F5 5D AE
 DB E1 4E 03 45 D1 ED 0D 79 24 D8 EE 5A 93 60 6B
 25 D4 55 F8 66 6F 1B 07 3D 3E 46 9A 58 EE BF 22
 55 4B 86 99 7C 6B 91 43 80 D8 40 F6 6B 7D E5 BF
 84 97 9C 2F FA 78 4A C5 7D 2A 65 A1 66 66 C7 00
 E3 C1 E1 19 38 E0 4D 99 05 FF AB 3F EA E5 C9 CF
 75 1B 37 A0 AE EC 19 4D 00 2F 8C F3 57 79 DE 4C
 84 A9 59 5A D3 24 EA 95 91 E6 B2 D7 91 07 C6 C5
 8C 1D 3D 01 09 C0 F6 B6 0B 08 61 2C 73 EF FE 19
 51 31 99 19 7C 46 F8 18 C7 17 0D F0 79 3E D3 03
 8C 03 92 BE 1B 95 56 87 3E FB 09 B7 38 84 85 00
 00 C7 8F 70 78 66 74 F7 A7 AB 71 E5 2D 00 54 54
 EA F7 4F D5 69 89 F6 FC 6D 06 C0 0C 93 E5 90 0D
 2B 87 06 16 8C 74 6A DC F2 DF 4B D2 D6 14 BA 0E
 CE 8A FD 3C EE 29 BF 4F 04 64 8B B6 39 76 E6 3E
 FE 25 2D 5A 61 FE E9 26 C5 64 27 FB 9C AE BB C1
 A4 42 83 EC 2A 92 FB 65 F0 57 F9 59 AD 09 D8 3A
 0A BD 21 31 90 65 3F DE 2E B5 06 CA D7 B4 29 04
 92 94 0A 4F A1 59 03 D2 B3 B0 A5 2B 11 DE 3A FC
 18 36 AE 9D 27 3E 34 AD 81 F6 95 64 49 C2 F5 63
 94 5D 0D 37 65 FF 32 9D 0D 04 68 DA E9 5C F7 DF
 AE 81 95 61 C3 35 8D A4 8B 27 C2 83 16 B0 D5 8F
 D0 B7 CB DC 10 21 AD 6B B4 AE 6E C5 CB 4A 5F 2E
 D4 5F B9 5C 4D 39 B7 47 61 7F 76 EA 3F 2D A4 5C
 5A 07 5B D2 E4 9C C0 06 73 38 58 AD 34 DD 71 AD
 FC F5 3B 52 BF 3C 30 9A 9B B6 58 1D 2D 33 79 89
 D2 11 2E 7E 49 1C 9B 4D B7 93 B2 EB E1 2D D2 42
 FA BE 22 A0 CE 1C A1 60 CF 5F 60 29 58 78 06 49
 31 29 CB 1E 45 16 4C EB 31 A0 51 87 64 A8 E5 A1
 ED 03 55 06 74 A3 76 4F B3 36 E6 2A 72 E4 1C 04
 CC D1 7C 6D B6 1B 42 39 0D 7F AB B4 22 D4 0D 1C
 15 DD 0B B7 81 10 EC 86 AB 4A 0E E7 BD D2 FE A4
 DC D4 62 F5 DF 13 40 65 B6 30 14 C9 20 15 34 B0
 03 A7 7B 60 D7 1D 8C 2A 89 C0 A0 07 DC BA 96 B4
 DD 3B CA 6F 96 F0 1A 8E 7B AA 5F 6C AB 65 5C E4
 10 BB 02 C9 08 2A 85 B2 AE 83 FB 5C AB 47 3E 4B
 2E 28 62 14 2F 3A D7 7B 4B A2 7B 30 8F BC 44 21
 FE 2A 48 89 4A 3B 32 BB A9 3F 20 A6 1B 9B 2D 43
 EF C3 D5 32 B0 CC BF 4B AE F8 73 BF 4D 2B 7A 7E
 69 77 D5 11 D6 FD 5D D3 62 69 E8 C1 2E DD 51 94
 DC DB 17 BF FC C9 1B 12 E1 86 73 BB 4A 8B C3 61
 4B 54 77 26 03 AC EF 9B 3E C5 09 95 A7 85 64 7D
 C6 65 5E FE 67 DF 4C 31 0A 7F 35 C1 FB 4D BF 91
 BE 3C 9F 67 7E FB 42 33 73 37 33 D5 9D 54 17 45
 38 CF 4B 1E 8E C3 A6 C5 32 1E 8E 39 44 D3 C8 64
 6E 92 39 25 DB BF 37 E3 DB 2B 18 47 01 E8 08 F9
 23 FC D1 5E 07 94 04 98 14 43 3B E0 FC C9 A7 6B
 33 EA 0C 9E CD 8C 61 36 C2 18 96 AF AC E7 14 8F
 2F 8C 6A A2 0A EC 70 0B 6E 51 9D 79 DF 67 14 74
 CC 75 F6 C5 D0 25 AD CD F0 AE BE A2 62 DE 4B F1
 1E 8D 8D C2 0A 7D B5 44 15 F4 02 EA 6A 55 F2 2E
 84 D1 1F 4B B5 27 36 DA C1 03 FD 60 01 4B F2 0A
 58 A6 9D 9B 87 45 BD 11 5A 83 E0 B6 3A 74 AF 18
 8E 34 96 88 55 82 22 C9 A6 EB 79 F2 B8 3F D3 4B
 59 A7 CE FC E9 B1 F0 E7 FD C8 B9 0A 16 7C A3 DA
 4C F4 86 13 A8 DA FC 92 E0 F2 7C 71 0F 57 6B 6C
 1D AE 99 AA 09 69 55 13 46 E2 C1 3D E2 89 70 B4
 08 9F 04 1D 7F 03 17 62 3E 95 86 FB 89 3F 50 38
 F8 86 00 F8 95 CA 4C A8 90 F3 B3 34 60 23 38 7B
 BB B2 B9 AE 92 64 FD 3D 17 77 E8 73 6E 82 45 0A
 50 BC 42 B1 59 B2 1D E7 D3 28 97 6A 3D 56 A1 B4
 D9 05 BF 8A 33 1A 39 C3 34 CF 32 FC 2E 8F 15 F4
 1D B5 DD AE 68 60 88 B0 FA 8C 72 85 BE 40 37 0F
 EE B1 F4 58 36 D2 1F 3B CA 19 0D DF 14 43 A5 E6
 44 DC 85 55 CA CF 06 8A CF 9E C1 B2 70 B5 DC 56
 FE B8 E7 EE 51 02 92 47 F2 D0 8F 16 30 76 3C 0C
 66 73 B9 F4 FB CD 62 32 62 34 38 95 36 21 DA 1A
 2F 5B 66 BD 89 B7 6C 86 B6 C9 43 B6 C3 92 59 B2
 60 95 68 1B BE 84 E5 AD B2 7B 7E A3 39 67 38 AE
 01 77 B8 25 AA 3C 33 0F 1A B9 8D 14 E7 6B 21 62
 49 48 31 79 18 9B D2 F5 99 7F FA 7F B8 E3 4B 44
 F4 83 4D AA B6 A7 89 C3 F8 CD 6A EC BB CD A4 6F
 2A 48 73 52 3A E2 68 1B F8 1E DA 52 9D A6 05 7B
 80 17 A4 0D D9 E8 F9 B5 4A B8 D3 EC FC C8 7C B8
 4C 8B E3 B2 40 6B 68 5A 2C 9D 3B E1 C5 A9 1C 1E
 E0 70 EB D3 54 C7 8F 72 26 8C 93 49 DC A9 46 B6
 FE EC 3D F6 3E 72 FD 6F 36 4B 40 19 5E 5A C6 5F
 49 C7 C7 26 F6 43 C2 C1 33 ED 18 22 FE 4A 33 F7
 4E DA DB FF B0 CD 0F 34 99 E3 88 56 88 0D F7 C1
 FC 6F C9 CB C9 18 69 37 FE F3 45 7E 36 7B 21 36
 34 58 1E A4 91 5D 70 5A 1F 3B 68 73 D1 BE AE 22
 95 11 65 B9 92 CB AD 58 D3 F5 F0 9E 98 E4 EA 7E
 3F 42 F0 63 38 EC 77 3D 6E F0 02 46 76 58 9F 2B
 B4 30 8E 4F 85 0D C0 39 2F DA 72 BB 1E DE C6 91
 CF 62 54 25 6A 60 6A 40 0D 55 79 5D B8 BF 79 E7
 9A B8 DA 9F CD C6 5B ED 2C 0F 8C 97 BA A0 E5 06
 42 71 CE FF 5F 51 E8 71 A6 E8 06 17 CA B4 4C 8B
 80 27 39 BB 32 76 A8 E6 67 8C 44 DE 2B 9F 39 B9
 6C 41 1F A5 51 79 5B A2 9A 69 58 28 61 16 11 C2
 A3 B2 5D 1F 00 83 84 E8 96 A1 29 CE 85 3E 94 93
 7D A7 56 B1 D8 64 36 FA 98 30 3A 60 FA 44 CF 09
 00 21 49 98 6C 44 2D 63 30 74 DD 6E F2 1B 5D 74
 FC AB C1 09 2C 65 71 7B C1 9B 48 4C 1B 8E 26 2C
 76 80 71 3B 8D 4A F6 0C AB A0 16 91 5D 77 3E 9F
 1E 28 DC C6 1F 27 43 31 04 D0 54 55 46 8B 39 FC
 4A DE B1 18 31 8C 30 79 5A 04 EA CE 2D 6F 01 3E
 0A 73 2E F1 0C 23 7B 68 4D BB D6 CA C1 CB 14 91
 F7 90 F9 9C 46 A6 04 72 57 71 56 8F DB 43 02 BB
 B1 7F 0A 5A 2F 0E EA 61 F9 AC 21 75 58 03 2D 25
 73 87 31 05 B3 1B 03 BD EB 49 EC 6A E6 67 72 C9
 3F 4F 03 3C FD B9 20 17 4B 95 36 8D A1 36 5C 0E
 E4 01 06 DD C5 AC D5 5D D9 27 B0 B1 E9 69 3E 92
 00 00 95 6B 49 AD 56 D0 77 9C 16 A1 81 E4 27 05
 07 22 E1 2C 74 88 26 ED 39 BE D8 46 AC 24 0C DA
 4C 5C E1 A8 FB F2 EB D4 94 AF 48 42 1B 9A A7 80
 51 F0 F3 2B 37 28 7E 12 5B 97 DF 34 E0 A1 AA 56
 6A 34 74 FB 9F 95 0B 7C 1E 31 78 09 03 EE F1 FB
 DB E3 4A 44 A1 A8 05 BB 1A 95 41 1F 78 5E CB 6B
 C2 E1 F3 C1 18 DA C8 92 01 12 B5 5B 31 CA 07 4D
 58 BD 68 25 6D ED 98 D5 0C 80 34 62 1C 35 69 4E
 EB 52 6E 08 2C 3E B7 67 46 3D 71 0D 22 07 7F 3A
 9D 40 BC 0E 0F FE A9 BA 16 DE AB FC 59 01 2F DF
 92 E9 72 41 98 4D 2A 5C 13 C3 A8 2A 5E 31 32 A7
 64 C7 30 D9 3C DB 1F BA 61 0F 52 F0 EA 20 14 D8
 DC 7E BB 8A FA 8F 52 F1 C3 E4 6A 98 86 47 2F 9C
 9E A4 13 92 18 11 9D E9 87 79 9B 41 A4 00 5F 38
 15 4D 0F 0A 50 74 A0 EC AB A0 68 36 12 9B D0 56
 83 4C C9 EA CC 76 F2 5C C4 3B 9B 0B 36 69 C7 E3
 F9 7E ED 48 7E 87 41 88 11 56 FD 13 92 1F AB DD
 8A E3 14 C6 4E 9C 8D 87 94 1B 34 16 B1 51 65 F3
 E3 83 4B F1 27 A3 FB 79 E8 40 43 D2 2C 65 D4 7D
 DD E4 1E 7D 0C 01 69 22 81 0E 82 36 49 14 A9 62
 49 62 6A 66 EC 03 E7 B9 D7 1D C4 78 38 29 2F 1A
 20 BB 84 BB F3 35 E9 72 A2 E3 E0 1D 76 2E 09 9C
 54 BF ED B6 85 C1 3C 58 88 2C D6 4A 64 3F 1F 4F
 E1 02 87 33 B8 09 F7 FE 8A 6E 0E DE AE 8E 4D 1A
 D1 D0 88 49 BE A8 D9 C9 1F 79 03 27 5E B9 4D EF
 4F C7 F3 B6 A3 5C FA 4D 51 B7 98 3A 23 E2 3A 74
 D5 E5 F1 28 0C 3C AA EF 45 0C 71 85 3A 51 42 88
 3C 7D 76 50 32 69 3A 62 AE A9 FD 83 E3 EE 05 BE
 5A 77 90 20 0A B4 70 3F C7 8E BC F6 69 BC FB 50
 69 86 A9 BB 96 2F 7D 07 DC F6 25 19 3F A3 B3 9F
 12 07 7A 2D F9 C7 71 CE 79 06 AA 27 16 94 73 59
 80 35 9D 2B A0 6C 11 DF 57 06 2D 83 DA 5C A4 36
 47 7E B6 3C 66 F4 F6 E4 12 78 EA 1F F9 20 08 42
 11 8A 52 73 F7 40 D7 B6 E9 5C DA BE 0F DF 6D 27
 D1 C8 A3 A0 05 1F 78 AA 67 7F 54 CD E0 5A 94 F8
 F7 EE 4C A0 B8 7D 4E 98 0B DC 73 0E 02 6E 22 21
 01 9C 5D 6D 31 9B DD 7A 49 28 2F B5 7D 67 F0 18
 45 91 38 19 8F 55 D5 50 79 75 14 58 67 2A B4 56
 C0 6D F2 1A 2D B7 90 AA B1 C2 6D 91 37 4A BE 70
 EB ED 12 80 D0 7A 8E B4 5B 11 68 65 21 2D 16 8D
 EC 73 81 0B 72 D5 D2 EE 59 E6 78 64 CD 78 A1 D1
 3C B1 FF 46 73 64 A8 F8 F8 55 7B 70 D0 A7 21 8A
 0E 64 0E 5A 9B FA BC 57 C5 E6 3E 7B F8 6F 16 64
 27 41 83 19 B9 6C CB FE 2F 38 D9 44 5B 0D 7B E4
 C2 87 9E D4 C7 B1 44 8D BB B9 06 E2 00 D0 8D FE
 9C 6B B1 4A 51 5E CC F5 27 EA 78 AC 33 23 89 B9
 57 DC 15 70 11 61 65 4C EE A2 17 B3 45 C8 47 D1
 3D FA C9 8B 91 8E 48 FC 86 F1 B4 4D 0D 68 25 C5
 F2 21 6C 32 A7 8B B3 68 3A 05 F4 E3 F2 8E 7D 2A
 33 70 22 F5 FD C9 8A 6F 04 7D 55 D3 D7 EC 3B 31
 20 AD 3E DA BF 7D 9A 6F DB 74 5D E4 3B 98 0C 5A
 E5 FB 51 87 56 2C 37 10 B8 97 A2 9B 9B 8E 51 74
 A4 B2 8E 58 CE EE 29 E5 00 F8 BD BF 86 3F FB 7B
 5C F2 4F 35 EB 0E 19 F8 2E 97 A3 93 1B AF 5A 18
 1A BE 74 13 0B 7F 91 F4 1E EA 03 A0 80 B4 38 D6
 6D 68 FE BB 09 12 6D 85 6F 11 78 1E 20 7D CA E0
 26 EE 3B 13 76 C8 52 D7 EC BD CF 99 EB 19 9A 1F
 B3 93 B2 D1 6C 56 B1 88 59 53 DF 1A 22 2C 62 8E
 50 83 C7 40 4B 99 FD 49 99 39 5D AB 3A 21 D9 C1
 38 90 C7 CF 4A D6 17 E8 63 8B 86 2D 99 21 7B 7A
 22 67 3A FA A5 0D 61 AD 18 22 D6 1E 04 EA F6 CB
 F1 2D B9 15 84 67 5F 29 26 7E 47 95 78 53 2D 56
 4D 43 7C 0F 52 AD 48 01 FC B6 A6 D7 09 B5 25 47
 A5 E1 8D AF FE 12 4E 3F A8 9D 7E 5A C6 59 AA B2
 96 77 5B CD AE E6 72 DB 30 9C 80 0E 5A CE 66 CE
 69 17 5F 4A 44 CA 8B DB 9C BB FF 4D 3E 5A 70 92
 E6 BD 05 8A 6E 04 2A 48 73 AC 9B D2 E4 9C 94 D3
 D7 BA E5 63 CE 96 9B 26 19 5C EC 3E 4C A1 1A 3D
 FE 20 53 45 BE 1F 40 6D DB 38 14 C2 E8 24 3C 42
 5B F6 73 A2 89 3C C3 41 5E 8F 42 DE E1 33 B8 59
 2E 75 09 DF 4A 22 FF 84 6C 8E 6A B5 6F BE 3B B2
 01 63 0D D8 2C 00 7E 6F A9 75 95 8E EF C9 7B FD
 69 4A 4D 05 BD EC 8B 22 12 50 DE 57 0C 95 D0 CD
 B9 4E 6A 95 E6 96 6F 09 85 63 E0 6D 99 37 4F FD
 A8 CA 2D B2 24 B3 98 25 53 F2 56 7A 40 5B DE 98
 56 BC 00 7F F8 8C 1E CC 2F C5 C7 88 2A 92 98 9E
 D8 08 C3 8D 4D 52 32 0E 5F 5F 88 83 39 A4 0C CC
 18 A4 0D 0F FF 83 59 03 44 D3 17 BF D4 FA 85 00
 4B 99 30 71 86 7C DC 65 7F 56 5D FD 1A 16 BC 46
 2C 38 F9 5B 87 97 71 3B EC 7C 44 7F F8 F1 D7 DA
 77 80 EB C8 D6 26 78 8C 26 87 25 3E 21 E6 FF 60
 A2 97 86 4A 87 0B 09 16 8E EA F7 2B ED 56 2B B7
 5F EF DB A3 F1 D3 B9 98 49 47 3E F8 E7 40 7D 45
 16 0A FB 0A 4D 53 F4 D7 B4 AB A5 4E 4B 9C 93 36
 54 AC 1A 7D 82 F6 02 5D 24 19 69 03 BB 4E 9A B1
 F4 C1 7C C0 4F 29 F4 E2 0D 06 B9 28 62 11 BC 18
 66 CF E1 2D E7 C0 46 1D CE 06 51 C9 4F D7 AA 9F
 01 4A 68 C3 E2 64 F7 9B 80 06 3B CE 9C A6 E4 45
 89 11 3C 58 85 5C D0 5B ED D9 01 75 A6 85 16 53
 AC 2B 7A E6 B7 56 4B B2 6B 2D 1E 9D 48 FA B6 AA
 D2 9E 23 B2 9E AD 74 4E C1 2C B2 DB 80 D1 5B 86
 9D 9F 31 4A B5 41 94 E9 1B 1F 81 94 CB DB F0 70
 BE E9 95 AE 02 1C 88 01 53 DC 5C B7 27 CB 04 FF
 54 6B 91 DA 2C 80 FF 8A AA 2F 1E 2B 51 93 70 AC
 3A 9D D8 A6 96 A1 FA DD DD 04 B3 3E 52 D0 58 FD
 53 8B 91 8A BD B6 5B D9 86 F4 7A 85 29 74 0B E7
 2E 2B 16 52 A8 DD 89 8D 12 F4 41 35 F0 A7 E1 25
 8C F4 36 71 AD A9 71 91 B0 08 98 0A 7F D9 4E 5D
 65 CB 59 50 22 0F 21 8E 1D 21 F7 60 AC FC 26 8B
 56 CF 77 08 19 A9 CC F3 20 EE B6 60 0D 7E DE 39
 B4 EE 26 93 F3 DC FB C2 5B 97 3A 1E E2 DA 98 7A
 34 C2 71 20 B3 B9 80 51 E7 70 93 F3 90 B1 12 AB
 1A 65 E3 C2 F0 4D 9D 0F A0 F5 00 C8 4C 04 B4 37
 19 CA EE B3 51 E8 AC A0 4F 06 FE 52 EC 8A 8B 87
 E4 27 B3 9E D7 FA A0 79 E6 89 53 31 41 46 DB EE
 73 AF 83 B9 0A 5C C8 AD 1F ED 59 93 8F 85 4A 8F
 39 DE 53 3F 48 75 D5 D2 51 A1 4E 8A 4A 09 01 6E
 1C A3 28 E0 36 9F 2A A5 84 DB 36 A3 0A 3F DB 90
 0F 2C 29 E9 84 23 A7 D4 92 B0 A3 DD 46 3F 42 08
 3E 32 C4 58 28 A7 BB 77 5D 54 C3 9B 71 60 A7 6F
 93 AA B6 62 D5 53 2F 8D EB EE E0 03 07 2B 5D 60
 15 33 01 AC DA 4B 79 DF E5 66 03 F0 DE 0E E9 71
 EC 74 5E C4 23 56 EF D2 70 05 B9 98 F9 78 E5 39
 E1 4F 04 22 E3 1E B7 B5 38 EF A9 2C 53 27 A6 F9
 0E B2 F5 3B 73 3A 31 A6 9E F9 86 F4 C0 A5 35 B9
 B9 5F A1 41 14 16 D5 B3 24 40 8F 45 11 1D 41 F2
 6C 32 C4 38 F2 41 82 9A FB 9A 5A 87 80 F6 C8 7A
 D2 50 BA D9 B3 95 EA 3E B5 98 1F 03 3B D5 AB 31
 6F 3E 69 7F 2D 39 EA 51 B2 F1 9F D0 C1 BF 04 10
 EB B1 BB E8 A1 A6 0E 2B 1D FC 4F 13 40 79 E6 40
 9B CF 36 3E 74 9B 2B 24 B6 40 F6 6F 4F 2D 87 B4
 40 10 60 EA F8 4F 81 16 27 E9 CA 3C B2 9E FC 53
 8C C5 28 AE FE EB 0B F4 19 74 F1 E9 D7 AC 1E 55
 07 14 A4 2D F3 38 4E B2 DB DA AD C7 60 CD 6A 77
 DE C2 56 CE 25 69 E3 2A 08 D8 8C D8 92 FB 5D 45
 BB 54 51 52 52 CE FC 49 D2 B2 A0 5A BB 43 05 70
 58 20 1D 24 34 E0 E6 20 6E EA 77 E9 F0 1F 10 94
 16 3E 4E D1 CA 45 77 FF 95 44 A4 5B 58 E3 20 64
 42 94 9F 00 16 58 D1 8F 65 AA D0 72 A4 D1 60 E9
 FE 27 70 FC F7 36 DF D4 54 11 8D D9 76 EA 9B D6
 5E 76 DF F8 96 85 6D 81 4A 9B 96 7C 1D 12 47 B4
 F1 8F 01 96 E4 30 2A 62 42 19 E8 ED 75 35 17 B0
 EA 4C 91 E6 09 0C A1 85 C9 CA 10 D0 67 3D B6 31
 03 59 AB 0F B8 49 11 2C 07 C7 AB 32 22 BE 98 49
 7D BA C9 BF 2A 0D 09 1E 63 EB 9D FD 9C DC 2C C5
 23 CB 41 FA F2 82 14 A3 36 ED 61 6F BE 8B 37 0F
 BB C9 2F 32 33 C0 B8 88 0E 4E DC B6 14 F3 BC E9
 84 3F 92 DA 7E 90 B2 A7 18 1D 4C A4 6D EE 1A 4F
 1A 8E BA B9 4B C1 1A 8A 90 7B EA 09 BF 02 A1 21
 7F 83 61 DC DF 37 AC E8 29 E6 02 2A 11 CA 5E BD
 51 E8 9D 33 A9 94 70 D0 88 82 2B 1F 24 E2 0E 2C
 70 6F 6B 43 E4 1E F3 BB C8 EC 60 1E 1B 23 BB 4C
 3F 31 3A 7F DB 63 B8 99 58 38 E9 21 D4 A1 68 4D
 6D FF 66 F1 99 A7 6F 54 14 35 9A 6A 00 E6 BB 59
 C8 F1 45 A7 9F BC B4 14 21 46 2A 16 B6 4F 2A B6
 C4 48 1E 56 67 FF AC 85 80 B6 88 9E 40 50 15 11
 93 C3 F7 DC A2 46 A3 06 FA 27 32 47 7E F2 BE 18
 62 85 F2 61 8C A3 6F 4A 72 35 AC 01 99 45 E2 6E
 14 9D 60 CB 88 74 80 99 33 67 12 1D 00 03 E4 50
 D5 CF 4F F6 70 B5 77 40 80 45 C1 22 AD 9D A6 11
 64 F4 F5 FA F7 37 A6 54 DA 67 5B FC 72 C3 7A 0C
 77 97 DE 2E 75 89 96 D3 B2 19 45 B5 C6 CE F5 76
 1F 05 96 61 DF 54 AD 36 7B 8C E8 B1 1F 9A 53 71
 4E 50 84 F2 76 B7 6F 70 5B 4A 5F 37 73 CF 3A D6
 B3 F5 1E 54 C9 AE B6 13 BB 91 C0 3E 05 AF F0 7B
 F0 DD 05 8D E4 64 4E 75 81 14 A2 8F F8 6A 6B 03
 1B A0 2B BB A3 DF E4 06 C9 33 B3 53 D6 A4 72 A3
 A6 BF FE C3 1A 22 7E 5F EB 20 6F E0 98 0A 04 6C
 B3 86 65 7C FE 55 A6 B0 E1 9E EB EE 0A 4E 9A F5
 49 75 DD D8 60 B7 9C 3E 65 93 60 9A 7E CE 45 5F
 62 B2 50 6B 0A 0F 1F ED DE 73 A5 AB 01 0F A8 3E
 A0 61 9D 07 36 66 5E BF B7 71 D9 A2 85 09 6B 42
 0C CE 3A 3D 71 B5 14 FB E9 F0 2F B8 2F 08 8C D0
 35 80 F3 CB D7 D6 8E 2B EF EB 21 D6 95 9F 8B 06
 27 0C 36 05 69 A6 6E FE B1 BA FA 6A F1 6D 3A DB
 D9 72 20 27 22 80 29 36 D6 8C E2 A7 6E 3E BB E7
 8B 2C 24 C4 4C CB C6 57 79 ED 33 6D 24 71 12 B5
 6D E8 D4 23 46 AC 6F 71 92 D4 6E 7E 79 44 EB 32
 4C 89 51 96 6A 3E 21 6C 52 E8 AC 26 5F 12 96 3C
 99 25 3D CB E2 63 BD 3D A4 14 E4 CC C2 18 DB 37
 08 FF DC D0 CB C4 0E C9 2D 9B 28 C1 AC F5 50 2E
 67 D2 E6 FB 60 8B BC 2F 72 4A 99 87 1B 47 DA B9
 AB AC 1C 26 AB 8A 55 7B 41 63 29 DF FB 78 D6 BE
 DA 8A 6B 49 4B 1E C9 20 11 93 BD F9 71 18 63 14
 D0 62 0F B5 47 08 EF 82 27 C4 A0 BE 9D 89 9B FA
 0F 38 29 D0 F4 D1 A4 4C 1F 22 04 25 96 B5 B3 30
 86 F7 90 FF E4 85 49 41 EF 4D 7E B6 19 AA 45 0C
 69 B8 DC 7C F3 25 FD C0 62 76 10 30 DF 85 A4 B0
 22 50 AC F5 F8 40 72 60 CC 20 C1 5B 97 4E 95 51
 05 83 D6 B8 67 C9 6B D6 21 CE 5A 1D 0F F1 D4 81
 2E 0C 3C BA 25 6E 43 86 77 9E D7 3A EE 23 12 0F
 86 C8 92 07 4A CC 6B 60 88 BA 6D 5D AF 9D E3 CF
 E1 D5 AA 5F E8 7E 92 74 F9 DB C8 7B 3A A0 6E 34
 ED E2 7F 7B F0 67 95 2E 77 33 47 06 81 18 B4 60
 E4 99 14 3F D5 5B CE 61 B5 9E 05 42 AA 3F 18 3C
 9D 8B 00 A4 0E BF BA 50 31 E9 7A 9C 18 BE D3 9C
 C6 4E 38 85 35 86 B2 40 0F A1 CD CE C1 52 CC 3F
 48 0B C9 C0 36 44 44 43 C1 94 D6 94 DF BD B1 5B
 0B 6E 44 70 C5 79 D5 27 15 CB 53 D4 62 11 33 1C
 3F A1 56 20 4E 5D C5 09 76 BE 2C 8C A0 13 50 3F
 9D 5E 3B 7D 9C D2 7E 19 83 0A EA 2A 40 10 CC 33
 8C FF 2E 37 0D A4 90 3E 02 C4 DD 95 9B 98 9F 45
 3C D4 60 97 AF F0 8A 19 73 B7 D6 E8 D0 D3 97 2F
 CF C0 4E 90 C1 7F A8 DD A9 1B 53 B4 2C 38 E9 8A
 26 6B ED 33 B4 00 35 DC D2 E6 A3 E5 69 F4 65 A2
 54 08 98 8F A1 BC 85 3C F5 E3 19 A1 37 53 BD 85
 A1 3E 6C 8A BD 9D 81 97 82 94 6E 6A 4D 28 5C 25
 75 A3 3C 43 94 31 C6 AD F2 14 AC 03 70 50 CC F3
 DB EB 23 55 DA 3E 06 0C 5E 92 2C 5C E9 78 F8 8C
 B5 17 3F 2A 45 8F 65 1B 7F D4 2D F2 DC 13 28 18
 28 CE 8B 02 06 72 43 EF D4 8F 32 18 36 71 1E 36
 62 D3 9B D7 4D 5B 31 DB 9B 84 4C 44 87 E6 A0 80
 86 F1 F4 B7 84 80 38 7B 5A 83 81 33 58 41 A1 BF
 42 19 C8 7F 35 94 7C C3 68 2D DA BA B3 76 C0 9C
 59 FF 87 14 16 5F 6E 44 07 98 E3 51 98 65 F1 51
 C1 A0 89 74 37 96 84 C3 A5 5A BA 44 39 5B 70 4E
 2E 6E 6C 04 C3 9D A6 A9 65 E6 50 03 6C DD E8 B6
 FB E6 27 C7 7A 3D 72 4D BB 0D EA A7 E6 DB 70 83
 77 0F 99 48 B7 7B 76 A6 DB B9 3E A8 6E 27 1D 6E
 5A E0 03 24 0C BA 76 BC DE 83 34 8F CB 4D 02 BA
 34 57 08 4D 5C 48 38 07 17 0D 12 E4 4F 95 86 62
 3D B6 11 E3 9E 80 1C B4 EC A3 23 7D 75 DD 04 2A
 AE 75 28 16 7A 5C C0 B4 4C A0 E9 AF F1 72 85 DE
 BC 3F EE FC 38 BA 01 8C 9A 8D 73 57 AC 1F A9 AA
 3B C4 C4 9B CC BF B1 D9 4A E8 37 8D 57 6F DA 6A
 5C 9E 5E E3 FB 8A A8 3E 7B 56 34 FA CC C4 33 AA
 D6 AD 8C 1E E6 D6 14 4A 00 F6 21 F7 1C 82 33 68
 34 85 DA 43 6B B1 47 3F 5C 49 62 20 A2 B5 9B 09
 68 D3 0A C6 42 50 81 4B AC 07 FC 73 90 68 1C 13
 CA B5 94 29 01 CC 4C 9D 00 11 65 4A EE 25 3A 5B
 A1 E9 1A 88 06 25 72 21 A3 6F 57 B8 00 3D 08 B5
 3F 2C 9B B7 74 AD 7D B9 8B D4 80 74 06 3E 3E EA
 F4 16 8F 5F 3D C1 D5 20 1E 7E 65 53 8E F1 08 6A
 7F 5E A8 86 41 17 58 97 CE DD B3 E9 B4 45 AB 0B
 F6 18 95 EC 44 D3 8D 46 FF 43 B3 EC 4F 10 11 FB
 E4 B5 72 EB 82 61 61 0A 1F BF C1 B8 82 08 99 97
 D5 59 DE AB 57 AE A2 D9 81 30 53 92 35 FD FB D9
 2A F7 D9 37 E4 6D BD 20 82 42 F4 0F 56 F9 71 70
 DF 5E 61 FA C6 FD F9 97 E5 7C 1F 9A 1B D3 20 C7
 E7 3C AF E2 74 5C 9A 3B BE 34 F3 73 1D 8E CD 29
 94 4C 9E F0 80 D6 D0 C5 86 AD 48 E2 41 B3 5F 50
 2A 4E 86 1C 13 61 6F 42 ED 3D D5 E4 F9 60 33 74
 FD 69 BE BB BC 8A 1D BE F2 CA 34 09 73 0F E7 79
 BB 34 EF 6E 95 BE B6 AB AC 3B F2 67 F2 A2 66 22
 F6 51 36 91 57 B6 4F 97 C9 8B 5E 17 C2 0A C1 82
 67 BA FD 94 32 F9 A9 63 5C 2E 8B 2A 34 84 86 DE
 01 49 57 C6 2D FC 68 2B C1 43 19 BC DD C4 13 8B
 35 FF 3F 39 9E 06 9A 54 CD 37 20 94 E5 9E D7 4B
 07 55 55 45 07 EE 68 D9 5B D5 63 54 39 7F 6E 11
 61 8F B8 A6 D6 7E EE 46 55 4E F0 AE 6B 65 4B 49
 80 8A 16 34 6B EC DC 92 E0 E1 E2 33 65 D7 98 2A
 57 7D 46 8B 3E AF 6A 4D 31 11 36 5B C3 A8 F1 B8
 81 B7 00 87 E8 02 29 97 0D 05 C1 79 42 B0 AE 9F
 3C C4 06 A4 61 B8 3F 7F 52 DF 42 8B 90 F5 2C 12
 5F F0 FC 54 8C 91 7D F6 62 7E A4 91 4F 9C 47 A1
 86 CA 87 28 32 9D E6 5C 4C B4 85 00 B3 A0 E2 DC
 F1 26 BC C4 3D 30 5C E1 EF 23 A0 0D 0D DE A6 C6
 DE F9 A9 E0 8A CB 71 24 FA 4A B1 4C 93 22 2B EF
 E7 3A D2 B0 54 47 9C C3 36 43 B1 27 C1 32 6F CD
 B0 95 D5 5C 3C 8A 21 4D FD DA 6D 17 C4 0B C5 49
 44 17 B4 17 08 34 4F 9A C1 DB 51 A0 14 CE AF A8
 82 CF EA 31 E4 A0 86 C5 F9 F1 A3 7B E0 DE BE 36
 05 A9 F7 70 21 CB 44 D9 EF 2A FD E7 8C CD FD 4F
 0D 6C DB D4 5E 01 50 4C 11 2E 77 68 8F E9 89 C5
 DD 71 F0 24 AE B8 21 B6 13 7F EA 4D 15 39 B8 FA
 A3 20 B0 4F 64 BC A9 F4 B7 8B 5D 9F A1 E2 9E D1
 FF 0A 93 E1 35 FD 5E 0C 9A 35 3B F0 1D 5C 75 4E
 00 0A 66 C5 FF A3 15 86 F5 C8 98 73 B0 EF 01 6A
 99 2B 0C 0E 66 FB 3F A8 1A 39 07 2A 32 02 D6 94
 87 E8 FC AF BC 9B 6C 4A C9 E6 F2 69 0E 6E EC D0
 36 DF CC 50 BA 8C 8E AD 95 DE BD D3 E1 EB 4C A3
 B4 0B 62 E8 28 A9 E0 9A 4D BE 04 9A C8 67 5A 58
 C5 A3 7E BC 5E 30 37 6C 5F 97 B0 07 8D FF BB 4F
 3E D7 53 A1 C1 37 CB 9C FB 06 5B 4A 3D F1 7F 01
 67 A2 46 1C 83 CD 93 DF 81 B0 BE F6 66 00 B6 68
 DB 45 06 69 B6 CF 50 FF 83 78 D9 D3 D3 65 46 58
 F2 48 20 1B 8B CB 30 5D 53 8B 6A 72 D8 6B C0 78
 91 E1 62 BF 45 84 B7 E6 EE BB EA 0C A0 20 33 81
 39 92 64 60 1C 75 C9 99 7A 76 7F F3 50 F5 F2 A6
 A2 31 F5 39 C0 DC 74 76 7C 6D 2B 88 06 5E 09 98
 FA 99 8F BF 8D F9 11 DE AF 41 6C C4 A3 E5 D4 21
 0A 94 F4 3C AD 8C 34 F7 62 96 50 C3 C1 CE BD 49
 E7 5F 32 4F 85 72 9A 52 EC A3 1C 1A 3B 32 99 95
 56 11 8D 0F 49 2D 67 C5 C2 4B A4 83 5B 8E 6A 35
 1D 73 A3 13 59 A2 C2 48 8C F2 5A E6 22 C9 B3 E0
 F0 10 FF CE 9D 9D F8 8E 0E 1D 23 73 CE B6 9C 5E
 B7 6A E5 CC 81 88 97 D5 86 43 A8 51 0A 53 D6 4B
 62 79 48 59 50 09 9D 95 30 79 E3 84 B1 8A 0B 60
 A3 7B B5 B9 89 E1 7A FA 3B 81 45 78 04 62 84 5B
 CF 2E 32 2E 14 39 00 58 FF 80 D1 30 4E CA 31 AC
 8E 92 3A DC 8C CA 85 FA C3 92 1C 32 15 15 EA 74
 0F 3C 22 35 85 37 2E 77 CC EE 02 2C 40 39 9A B8
 D0 30 A8 01 82 B4 BA 75 E0 54 D9 EB C9 B9 9B 7E
 3E FC C5 4B BB F8 D6 D6 56 52 63 86 96 44 F2 4E
 98 5F 96 85 1F 50 41 A2 C0 E3 95 94 4C 45 E1 66
 34 10 7E A7 9A D5 FA E2 B1 4D 58 B4 3C 58 A0 AC
 C9 87 5B 9E B0 A5 31 73 45 BB D7 54 E3 A1 97 A0
 3B 1D 14 FD 50 DC 9D 2A EB CF 01 F8 28 07 C7 8E
 BB E0 B8 23 B4 5B FC 33 DB 86 FB CE 9B 62 80 CF
 CB B1 24 15 22 F6 6F 09 B9 3F 74 AC C4 44 05 DE
 3E 30 F0 F4 C8 31 8A F3 B7 13 B0 3B E3 2E 3A E1
 27 A0 B4 40 5E DB 79 AC CE DD 8B DC 70 69 DC A9
 C7 28 09 8F F2 4D 47 48 BE 68 D6 07 AD 61 41 D6
 3B 6D 52 CC B7 B1 20 8D 5C 3E 84 E6 EA 8A A9 FC
 1F FB 88 78 E5 D0 2A B2 DF D5 E1 C8 76 E4 DC 59
 E7 D0 CF FD 44 ED A2 2A B3 40 47 40 4C F0 FE A7
 D2 9D CB D5 24 B1 66 24 6A 2E 83 C1 0E F3 4C C0
 6C A3 AC B2 57 56 22 64 4F 07 C7 03 38 A6 14 46
 5A 95 06 4A FA 45 5C 89 72 AA 46 FF D9 16 1F 6A
 7F 4B 1A BF D9 D8 2C 3C 37 9F A1 5F 49 06 31 6D
 0D 15 41 E7 7B 3A 25 09 43 C9 0A 2C 42 D3 21 99
 F3 ED 7C 56 A7 1A 3E AB 7B A2 AD 04 A9 CB 81 D0
 B2 1B 45 0F 7D 01 8D A7 78 08 DB 50 29 34 7F B3
 6F F3 02 7D 37 E1 B2 A3 D2 93 47 A2 FC BD B4 9C
 78 84 74 5C 67 34 01 82 21 5D 4B 3D 81 14 62 7B
 59 2E 08 84 EA 91 97 63 E2 91 77 8E 55 C7 02 A2
 B3 2C C6 68 18 32 C9 1D 6E 38 40 04 EE D4 E2 88
 92 ED 05 0E A2 A9 6E 5D A4 40 B5 33 46 65 FA 44
 8A 03 25 4F B4 4B 8D 0C 06 76 A9 65 87 9F CE C7
 41 1E 75 00 A3 65 A5 12 58 E4 0C 80 E3 4C 6D 5C
 D8 17 E9 47 C6 41 A3 AD 72 12 A7 57 2E 86 11 8D
 F7 ED 45 87 6F C3 B5 13 01 39 60 06 3F D0 6C 41
 B3 95 B4 57 D4 45 2D 0A B1 5B 6C C9 E5 EF 6B 64
 AB 16 4B FD BD 0A 87 35 4C 7C 7C 47 61 5D 44 32
 BB D4 08 9E 4C CA 62 CB E2 D0 52 41 DC E9 A0 F3
 B0 F4 7F CB EC 65 81 AA A7 EA B6 2A FE FE 39 87
 D2 DB ED 29 94 8D CD 23 00 F7 5C 30 DD 95 C1 8E
 54 BA E3 4D AE 50 EC 13 90 92 9F 88 64 72 14 5F
 2A 95 BB 70 4C DD 90 A2 4F DA 1C 0B 55 20 32 E4
 33 34 D8 E0 18 8E E2 4A BE 73 B0 10 83 82 37 A9
 CF 1A 44 2B 76 F7 28 14 23 14 3C 78 31 56 BF 94
 3D 60 B9 0D 25 24 3C 7C 57 84 5F 44 0E 61 4E 9C
 43 0F 0B 72 35 FB 04 0A FF E8 9A 2D A7 D6 06 DB
 ED 3F CD FF 64 0F 9B F1 31 C9 EA 0C D6 F4 65 23
 6B EF 37 1A 3A 32 EB EB E2 91 97 05 DC 3D A5 CC
 79 EE AB 34 69 F8 25 88 93 0E CE 1D 05 56 DB 44
 C2 32 61 64 93 B1 90 DB 54 2E B3 14 32 61 DF 7C
 FA 1E 42 0D 74 CE 85 0A D2 0F BA BD 67 39 9C 56
 14 D9 6B A5 56 80 53 7A F7 7F 01 AB FF 08 FF C8
 C3 66 41 18 BB BF 53 9E E7 1C AC B1 87 C4 35 AD
 83 DE DD C9 BC 0C E1 25 ED 5F 77 4E 6B 50 5D 77
 30 09 74 E7 91 DA 62 95 83 A6 99 30 7A 01 F9 0F
 92 69 77 81 2D 68 7C 6C B8 55 8E 58 66 0A 27 E8
 3D 08 39 38 4C 35 43 B3 20 FC A4 88 A8 13 0A BC
 5C A7 69 9C FB C3 26 A9 8B 58 88 60 7E 4B E8 EF
 C5 42 03 EC 68 25 61 BD EB E5 1E 13 17 53 C5 29
 77 83 D7 BD 97 02 1F 18 78 91 6E 19 76 AB D2 C3
 22 FF 45 53 8A E4 4F 0E 60 B1 17 4D 37 43 FD 57
 CA 9B 26 C9 E3 1A B2 9F 03 53 92 4D 4A DD 1E 24
 94 3C 2E 7A 1C A0 98 2A 70 D0 51 52 73 56 E4 9B
 72 5C 21 8A 15 49 D5 CA 34 16 77 C2 6E B0 8B C6
 1B 4C BE E0 77 63 92 E6 BD BF 38 AC 85 A1 99 72
 29 92 3C 5C F0 AB 2A EF B6 DF 66 0C 3E 5D B9 95
 9A 20 D7 69 35 B3 62 90 86 FE FA 66 02 E2 6F 3A
 C9 1C E5 A7 D4 C7 D0 FB BA FD EE 3E 5A 6D B6 A7
 AC B8 25 1F CC B5 61 12 DC 16 45 CC 1B 96 9F 88
 E8 56 D9 DA 33 93 54 85 F9 27 E2 6F 34 23 46 C8
 94 ED 7D CA 45 BA 4A EB 58 93 E3 63 FA DA C0 79
 9C 89 22 1D A6 C4 76 70 1A 2D 34 84 7C 4E B2 9A
 38 98 0B D5 7B 65 75 B4 4E 46 CA C5 50 2A B7 1C
 9B A5 2F AC 8A 16 EF 3F 5B A0 D4 1B AA 96 9A B4
 13 78 D2 67 4F 9B A0 C7 89 66 9D 4A CC 76 80 43
 5B 86 FA 8F 79 57 77 27 9B AC 35 BF 14 68 70 14
 BC A1 5E 65 AA 44 EE F7 3A 81 04 D2 BE 78 06 FA
 C8 B2 BE C7 E7 DD 61 E3 A6 A3 27 D3 1B 07 61 D0
 68 B5 C8 35 A4 D0 E9 07 1D 49 21 E0 C6 D4 9C 80
 49 6E 0F B2 E4 CB 0B BC A6 74 8A 6F 3D 6F E9 99
 66 53 C0 8B B3 16 57 D1 40 6C 44 AA 64 0F C5 2B
 2F 56 25 7E 76 94 B4 35 F9 49 D4 A9 EB 5C 14 D7
 F8 0F E1 04 2E 22 D4 C4 21 52 A5 54 FA 4D A0 84
 E7 9D A9 35 7B 93 DB DF C6 1D A8 B8 40 9D B3 D1
 A2 E7 53 55 C1 C7 FC 8D 9B E9 6A E7 89 0F A6 17
 0F 3F DD 1C E9 F1 52 73 CD E1 54 83 16 47 9C FE
 8E 6A 00 B2 F6 6D 46 DC B7 FB 6B 73 3D 66 E6 41
 CC 86 CF F6 FD 83 92 82 D9 47 1E A5 5C 53 EB 06
 07 94 8A 0E D1 B1 F7 32 0C 97 2A 50 AE 80 94 6C
 8A 98 9D 70 C3 45 79 77 62 AB 6D CC 75 16 EE 96
 54 72 9E C2 C7 59 2F 4A C9 FB C5 B1 D8 D4 02 05
 F6 7B 58 90 3F 53 9D 83 35 7A 87 5B 69 A3 74 AC
 4A 14 E9 8C 0C BD BA 93 44 C1 6C 91 F4 D1 0E DA
 97 FA 41 C4 99 50 49 C4 84 5D 84 6C A8 5D FD F4
 B7 A7 A5 AA 0D DA 1F C7 53 02 B2 F4 D0 7E 5F 69
 C4 05 F9 38 FA DB 5C A8 D8 7E B4 09 45 9C 20 F9
 73 E1 C4 E9 50 BB 5E 90 B9 A3 16 ED 17 53 0C EC
 42 3B D3 5F 9A AD 1D E4 E5 13 75 8B 87 77 34 57
 BB 5D 80 1F EA 69 9D 1F 1A 46 04 7F 66 7E A8 C4
 5D 38 00 33 E9 18 5E AE 20 FF 73 75 4D 08 5C 2F
 55 F5 56 D9 80 24 00 2D 9B EA EF 4E A7 88 A9 21
 26 9E 0A 13 BB FC AF 06 29 1B 88 AB 5D D9 87 DF
 C4 42 58 FE 13 23 51 C1 43 43 7D 64 9C 6B 59 66
 55 7D 74 1B 96 A6 E0 41 AB 4E 22 03 8B 39 5B C3
 05 EC 27 A0 E3 98 E4 BA 6B 86 11 7E 1A A9 59 4A
 0E E9 82 2A E9 55 D0 0C AC 91 9C 69 CF 2D AC 4F
 74 C4 DC 9F CC AB 4B 1A EB 56 85 1B 4A 8E F5 CE
 A6 54 1F 94 E2 38 48 CE B4 5C 32 F1 E7 F8 85 89
 B5 9D AB 1C 90 E1 B6 72 E3 EF A6 D9 FF FA 91 34
 41 3E F0 DC DA 9D E7 BF 04 C8 F7 CB CC D5 F7 86
 B0 CA EE A4 8E 51 50 FE 42 05 11 D6 40 6F 64 24
 D4 E5 E3 E1 35 2F 0C 80 61 4F 1E C4 2B 44 F0 9B
 69 00 0F 21 9D 90 7D 36 07 CC 65 56 07 90 7E 6D
 2D CB 8F 65 AE 00 C0 F1 E4 5B F0 66 B4 36 39 69
 41 6B 9A 60 6F B6 0E C9 81 6E 8A EA EA D1 11 E0
 52 F4 E3 DD 6B 06 83 7D 97 C2 05 22 CC 47 20 D9
 C6 CF 1D 85 60 B7 B3 FC BF A0 BD 9D 39 03 E4 C6
 12 53 EF F2 79 2F F0 9B BA 3E A7 97 30 05 31 C6
 0F FE 77 DC 0D 1C 1E 0E B5 7E A9 B3 DE 16 5E E7
 75 FA 03 0C B8 1D 97 23 57 07 A1 B1 3D E1 5A 70
 C6 39 86 CC 7B FB AE EB E9 AC 77 DE B5 66 2F 4C
 AC 46 B2 79 2B 63 6F 39 05 E0 A2 57 06 FC 62 E2
 28 BC 69 C6 D8 51 83 B1 EC 9C AB A5 0A 4B 34 18
 A2 37 A9 EB 7D 1C 99 22 41 65 36 E1 12 62 65 1C
 A6 85 CE 11 66 01 C3 17 C6 7F AC 2F 5D C6 C2 D4
 68 AD BB 88 D4 A9 2E 23 F9 48 BA EE A2 A9 FA CF
 44 4A 7F 3D 32 4D 8F 8A D9 69 46 50 FE 3E 5E 16
 51 51 65 5E 6C 3C 99 1E C2 15 47 70 48 49 E2 DB
 C4 EB CA CA C3 DA DC AF 94 A5 F8 FE C9 68 47 23
 33 1E EC 6C DD 39 D0 D5 D8 15 73 E2 22 42 8C 17
 F1 08 BF 94 14 F5 ED 81 DD 4E 7A 8F 89 2D 84 D9
 FD 94 1C C9 A1 55 8E 0A 89 B5 94 18 3C 3C FF 6D
 FA A1 EB D6 19 59 86 2A 62 22 C3 C2 A4 A2 AC 30
 2A 18 6A DA D3 3C 5E FB 4F 77 EA F4 30 54 78 AF
 C7 90 6C 1A FD 9B 01 B9 45 72 66 95 7A 81 C0 A2
 89 E6 C2 62 AB 78 34 E0 50 DA E1 AD 35 3D 90 29
 6E 18 82 27 A7 6C 7D 3D 3F 47 D7 12 E6 C0 62 0C
 BA 6A 94 9B B6 B6 82 DA 82 5F 6C A6 5B C6 8F 4C
 3A BD 4A 91 C0 45 53 97 9F 7C E2 1D BD 25 F4 29
 E4 B9 77 F6 2C 92 04 C5 61 85 A9 03 B6 21 D7 99
 F2 E9 F9 D7 96 E5 6F F1 B2 2C A0 1E 60 DA 60 0A
 A9 2B 90 F8 95 42 84 0E 58 12 F6 A5 25 07 F6 77
 BD 02 DC 8B 3D 2E BB EC BC 92 44 2A AE 45 57 97
 F9 6B DB D2 77 C6 80 E4 A0 AA E8 DC 63 0A 84 C8
 1A FB B5 D7 97 8D 6B CA 47 9A 2A F7 FE 9C C2 1A
 70 5D 33 61 F0 17 E9 13 D8 D2 B3 9E CC 41 3B D2
 C3 5B C6 DD 40 A7 59 55 3F 15 EF 9B DE 99 60 38
 8A 15 F9 6E F0 A6 32 B2 CD 66 2B 8D 4D E8 1C 53
 DF 38 23 0F A1 8C 60 F8 05 28 95 B7 D8 24 D3 11
 68 E8 D7 21 3C 8B 68 DB E3 ED 48 DA 48 72 61 87
 92 7D C9 75 30 63 90 EA 9B 6E E6 32 45 5C C9 A6
 54 EC 61 7D 3A 00 30 FF E8 CD 0B A4 3E 52 16 06
 78 00 8C 75 C0 46 95 61 4A 14 14 27 1A 9A 48 0B
 F9 17 9B 0B 5A 63 FA 62 AE 6E B8 E4 0C AC F9 5D
 07 DF 73 DC 3D 79 89 7D E8 92 49 CB 05 43 DF 3B
 45 F0 A1 43 19 3C D7 36 F2 4F 91 F8 02 11 D8 8E
 AA EF 13 2C BA 7D FB C9 30 3E A6 BE 74 C0 E7 C7
 F1 6C 1E E5 F3 F8 83 F0 FD 6C E2 BE FB E7 A7 D8
 28 F2 00 0D ED 27 97 AC F0 C9 9D 42 EA 50 EC 1A
 89 73 3A B9 3A AE CB 6E 67 19 42 50 72 E4 8E 21
 D8 50 86 F8 31 27 CE 8A 49 FD 52 06 8A 75 5A 54
 C1 19 2D 4B D6 38 2B 12 72 D1 44 81 69 98 7A 55
 45 98 EB 5E 49 69 F9 60 EB 22 BF 75 3D B6 06 C3
 12 0D 74 34 97 9F 60 9A 8C BB 4C 0A 73 C7 81 C1
 C8 5E F0 31 13 F2 05 64 E5 67 14 77 7F CB B0 87
 A3 7E F5 98 63 FF DA 7B D3 A5 6E 00 7C F9 CD E4
 2B 46 E6 21 C8 65 3B 90 71 23 AA CC 8A 4C E4 A1
 31 1B E7 3F 7C 8F C1 CA 28 2F 85 22 35 8F 98 8D
 EC BA 89 D0 5B 45 FD 69 42 3E CF 1F 09 DD 63 55
 80 6E D4 14 8E 4A 53 B6 49 B7 E1 94 6A 96 8C 67
 EF C6 C9 D6 FF 7C 72 47 3A 39 EF DE 22 F6 96 8F
 FA 7C EF 1E 67 74 31 D6 5D 19 AB 22 02 F8 E3 93
 BB 36 31 F2 B5 5D A8 C3 3A 68 D6 E1 5B F9 75 4A
 23 77 73 51 74 D7 65 FA 8A 27 CE 33 2F 64 46 B5
 EE 31 8E EF 8D AD B2 3D 9D 84 E2 88 0E 05 8F 11
 2F 95 DE 5E 3F 0E E2 E8 BA 42 CC 94 D7 55 27 04
 2E EA 0E 2D C6 40 58 F3 A3 6D 4C D2 7A BC D6 31
 F7 B6 65 76 2E BA C1 B5 CF 73 99 2C D5 66 57 3E
 D4 29 81 1E 19 0E E5 4E 70 22 5C FB 22 16 23 29
 61 98 65 92 A1 C0 A2 FF 1F 12 9E 6F DA 69 DD D4
 80 D0 BE 18 A1 D8 D6 FC 2B DE 08 21 2F 87 B0 EB
 FD 65 67 0B 45 D3 B7 C5 95 1E 98 AF 61 90 B3 2A
 F6 D4 03 FB 5B D0 E1 75 CA 1B 39 F0 A2 72 EC 2C
 E4 38 26 EF 78 F9 EC 80 06 7E E1 68 4E F1 8C 6F
 05 0B 46 A7 8C D3 A0 35 16 27 18 08 5E 1B 37 FF
 C8 CC FB C2 BA 19 8C C7 B6 87 42 1F 04 9A 3B AF
 80 52 8D 83 6E 5A 6D AC F7 B1 20 ED B6 2C 83 3B
 DE EB 99 49 B2 DE 78 B8 28 8F 47 77 2E 6C 86 D8
 AD 62 15 06 F9 F3 5B 5E BF B5 B5 BF 67 53 1B 42
 8A A7 E7 B6 8A 2D 57 A9 77 5D 2A 95 72 74 E7 C5
 01 78 56 99 E9 D0 0D F0 A5 50 0F 0A AE 01 1A 60
 B5 77 EE 31 E9 2E 7D 8E 2B F8 6B 6A F2 6E A4 D0
 C7 60 09 17 09 34 68 71 9D 4F AA 89 BF 7E 2E A0
 AC 13 24 D1 10 CB 72 B1 37 9B 28 19 A8 BE 5F CA
 D3 69 39 23 0E 98 9A B6 34 72 73 52 74 FC 85 F2
 35 30 3E 2F 7A A4 A1 F9 0F 30 C1 0A C3 BC 7E D4
 3F AC FA 29 81 CE 90 FB BA 98 32 D8 7E 6B 0B E8
 88 5D 70 AD 05 31 27 52 D3 85 CD B9 B0 12 21 2F
 3A BD C1 1E 1C CF DA 2F 34 26 7C 1D 34 23 C4 D5
 2E 8D 2E 09 0F 09 19 49 CF A9 D5 39 07 8E 14 42
 9E 03 45 CA 4B 4E 7F 19 42 65 2C 18 FE 64 F1 35
 99 07 D2 19 2A 9B CD B2 EF F5 CD 39 C8 93 B4 87
 3F 2B 01 23 B0 2B F1 7E A1 D9 9B 67 15 0A 01 B9
 2E A9 A5 E4 58 E7 F9 9D F2 AB 24 00 E8 E6 3A B0
 BE 91 EB 82 DB 75 A9 95 E9 0A F9 C0 73 5C 3D 0E
 61 2C 76 43 7C 85 A1 C2 53 97 6A E4 47 35 AF B9
 F0 EC 76 23 26 9C C3 F1 F6 5D C3 B4 D7 F3 1A F1
 90 8D A0 58 FD 7A 02 D1 C3 7C 38 C0 8A EA 12 68
 54 27 A5 33 4B 49 FF 3D 89 26 B7 3F 77 5B 07 2E
 65 92 9F AF A7 29 5D 5F ED A2 F2 A1 ED A2 F6 2F
 A3 03 84 41 7F AE 81 CA BE 4A 7F C1 4E 3B 5B E2
 BB 54 61 3B D3 E3 83 A1 62 2F E4 D4 52 2D 45 E8
 91 E1 BA 4B 3F 6C 3E 1F C3 A3 7A AD D4 C3 AD 92
 F2 F6 8C 03 AA 23 3D D1 B0 01 B8 C7 84 E1 F1 6C
 CC 1E FA 41 D4 E1 AE 72 F6 BA F5 28 CE D5 12 46
 7A A3 08 D6 D1 79 47 AA B2 32 AF C5 37 E6 B7 F5
 6F 98 17 DF 81 E2 22 B6 C7 E5 D3 FC 9D 8E 02 E9
 AA AA 9F 3C 41 A2 A8 F0 0B 7B A4 02 85 E8 BC EB
 F8 34 89 F0 EF ED 12 1E 59 81 6E ED 63 28 4E AC
 3E 2B 33 F0 8A B3 74 EA 40 84 EC 74 CF F6 1C A2
 43 0E B7 E2 A3 FB EA 24 EB 80 5D 1E B2 DB BE 8E
 97 B1 A2 C2 C2 4F D0 9A AA E8 BD 8A 9E B1 48 31
 7D 9A 76 2C E4 2A DB DB 63 61 55 1D 61 62 9E 83
 BD E3 14 AF E7 0B C6 AA 20 A7 C0 F5 5E 67 31 4B
 1F FE 94 F4 26 79 F2 7A 36 EC 6C 37 EB 25 8F 79
 6B 1C DC 8D E6 68 51 34 82 FE D7 B0 D9 DB 72 A9
 52 E0 A8 5B AB DF D1 A2 B0 A8 26 8F 53 85 97 79
 94 1E 36 19 AA E5 2C 0E E1 3D 92 56 B7 AF 00 DB
 1A B8 4E 4C 71 33 A3 E5 BC 94 3A 71 67 91 85 8F
 FA 95 40 95 9C 3C 7A A1 19 E8 8C 9A 85 B0 DD B7
 51 A0 BE 4C AA D4 2F 78 4F 47 F6 BF 7F 0E 23 4B
 12 74 38 8D 6A 56 3D 9E 05 D2 59 54 F3 69 B3 C8
 3A 13 8A 33 43 6D 47 94 EE 1C 77 F7 D6 26 96 86
 5B 74 14 00 8B E6 6D 37 55 64 78 5C BF E5 84 D3
 F0 A0 9D 49 56 E1 55 0E 81 F5 CA 7B 59 12 F6 D8
 73 6E AC 28 52 4E E9 C2 6C 1E 13 9D 3F 03 81 E7
 6C 25 E1 C9 5B EF 3C 94 3E 5D 21 58 5A C4 B7 C7
 90 35 DE D9 32 F3 CA 00 DD 8A 06 96 B8 22 2A C1
 FC 22 A0 79 E3 C8 2B BF BA CC DF 71 1A 52 E6 9B
 8E 35 64 E3 34 DD F4 50 D5 46 DE E5 26 B7 94 CF
 B6 60 DE 98 64 A6 35 65 BD E3 F5 64 E3 F8 BC 7C
 22 45 D0 72 F8 72 E1 BF AA 58 96 4A 44 79 E2 DA
 00 B9 A6 1B 91 AA 20 01 A1 E9 9E BF EB E1 8D F3
 7F 0D E2 45 01 87 6D 18 4E 87 B0 07 53 95 A2 49
 2D 0F DF 4C 7C E8 47 22 1A AD C9 EB DC 3A 29 DE
 52 74 4F C2 A6 04 CD 2D 51 1A 3D 54 45 32 69 3D
 4F C4 7F 38 2A B8 52 1A 88 D5 1E 36 48 C3 10 8B
 97 07 C2 BA 36 CE 0D 51 15 E5 B9 F6 9C E0 C8 DE
 22 91 7C 2C 49 45 E7 D9 66 DB 28 83 EF E8 0F F2
 2A 77 9E B8 A3 A7 6F BC 70 CD 3E 18 2A 09 81 61
 38 26 7A C8 F4 05 F2 5F 4D AB D4 FA 96 32 BE 9E
 C3 5E C0 AE CB 33 DE AE A2 E4 E3 07 07 8E 70 88
 10 37 BD 89 8B 74 4B 16 A3 1F 11 B8 29 1F 74 54
 81 75 D4 7D E0 7B 89 BB 97 C7 6A E1 1B 81 93 75
 80 6B 7C BC E3 53 7D B2 7D 5C 2E 8B FF 2D F9 FB
 A3 E2 9B DC EC 90 32 B4 DF 31 05 F9 48 BC 28 A7
 F4 9C DE 2F 1F 14 04 3B 73 08 43 5C 96 4A 00 45
 18 18 78 06 E1 B1 6E 69 83 E7 05 C6 C7 14 02 43
 1C C7 9D 51 CF 08 C4 1E 56 7C 6D 88 96 54 B2 4D
 55 D3 AD 07 75 D9 5B C8 E6 B3 92 BD 53 99 C2 95
 32 02 48 80 FC 03 74 D1 38 41 23 23 56 97 B8 82
 58 7D A6 AA 27 31 BE 47 1A 9B D7 E6 06 F4 4C 17
 32 3C C1 9B 1B 85 73 CD 44 D4 5E 02 67 EF 03 C6
 66 BA 2F 28 94 74 8D 88 6B 19 87 82 D1 BE 39 6D
 7C 0B 2A 46 BD 34 89 2E DA A8 03 19 33 04 1E CB
 4F 09 C9 5C BA 5F A2 92 80 1A 33 1A E7 9A 0E BF
 BE B3 CC A4 73 8B 3E C3 3D DA 4C BF E7 4A FF B2
 6A EA B8 85 CF DB 2B DC 5F 61 85 C9 78 42 3D 4F
 66 4D C8 72 7B D6 FA 4E 9B 14 1C 7A 98 76 7E A8
 A1 77 38 D3 49 05 B2 F1 49 76 DB FA DA 19 29 AF
 B1 A5 D0 3A 3C 25 14 13 73 63 6F 8E 3B 02 14 EF
 AF 65 5F 32 2B F6 13 F5 43 2B 17 E5 CB 27 03 83
 C8 9B 0D 27 ED FE E1 8F 4B D3 B3 80 82 65 7D 48
 7D A6 E7 32 38 B4 04 E9 4F 91 C0 3E DD 12 86 91
 B4 5E 45 6F 73 8C 97 A3 0F 26 D5 61 6E E4 64 31
 03 29 B1 B8 E7 02 72 05 DA 54 77 1C 76 D8 86 26
 E8 F2 25 71 0F 0A BB 06 7D DE 78 7A 35 37 ED BF
 CB D5 5C 78 6A BB 8D EB 9C 5B 3A 0D 6B 2F 91 8E
 6E C5 F3 7A 5C 94 60 CE FF A7 47 D8 22 06 06 6A
 C5 50 5E 30 CB 45 32 EA 01 6F 5B 9E AE 11 77 9F
 87 BA F9 F8 70 A9 BE 54 41 63 81 FE D4 E0 BE B2
 04 5C 75 A8 EF F3 12 0D 65 73 DF C5 EE 75 20 32
 24 BE CC 59 8A CE FA D6 4E C7 BA 30 89 DF 66 03
 4F 59 4F 04 D9 AD 2A 30 B4 1F D3 74 70 9A 90 C7
 4C 71 06 39 BF D4 BD AC BE A9 2E F1 0A E6 6F D1
 0D FC 7C 40 26 3F D7 6F 82 64 3D 79 3A 1B C4 37
 34 85 59 71 5D 8A AC D7 96 37 75 46 9E A8 D3 DC
 7F CA 5E E6 63 06 EC D7 66 C5 B1 63 48 63 2B 45
 47 F0 FA BE 72 FB 8D 14 8B 2C 6E 1C B3 93 EF 05
 23 79 F8 AF 93 5B FE A0 21 65 01 DA 8F 11 C3 83
 BF A6 00 C9 B6 0C 02 03 71 2E A3 6C 55 66 A9 C8
 F4 F0 CC C1 8F 10 F7 D0 86 FD 42 E8 5E F1 93 14
 C4 80 F3 BC 92 9A 9B 1E 4E 35 DF 48 03 ED 6A 9D
 34 8F 99 10 FA 93 DC 66 13 B6 75 C6 37 80 AE 4F
 27 4C 65 7F 1F 7E 80 45 D6 7D 11 76 F4 53 1A 5E
 FC 28 A8 DE D7 D6 4C D5 19 B9 F9 5A 13 8A A5 67
 4C A7 A6 EB CA 13 01 19 03 C2 26 9A 32 27 7A D5
 61 D1 75 D9 E2 47 FB 7D 66 C0 DF AE 34 2D 17 56
 54 9D 90 C2 C9 1E 80 A4 B2 90 DD 02 FE 99 3C BA
 FB 9A 27 0C 4A 8D 7D 9E D8 2F AA 7E 4E F4 29 8B
 0D 17 64 99 73 AD 03 1E 63 79 59 D3 83 AA 63 3D
 5C 1B C9 03 C0 6A 41 65 54 F0 06 3F 21 7C 88 9A
 1F A8 ED CE 15 F7 DE 2D EB 03 9D 2A 4A 06 57 A2
 E5 F2 AB 9A C9 11 D5 36 E1 68 DD 43 A1 7E FA 95
 F3 FB 77 68 40 38 D5 F7 90 8A FE 07 CF E0 53 DC
 CB 53 C0 2C 57 9D 51 BC E3 53 8F FE 1C 91 C8 1F
 0F 61 7B 68 E8 94 0E 53 34 F3 D3 84 52 0F B7 1E
 7F B7 D8 1A AA CA 70 6D AF A8 00 EE 77 A2 DA D5
 75 02 91 1F 6E BA 61 EB 0B 92 AC 5F A1 C1 38 AF
 D9 89 25 28 27 BE D7 D5 3B DB 1E 4B 3F F7 63 F9
 E3 A8 5A 21 BE 0D 46 39 B3 75 D5 86 38 9D 51 2D
 07 F7 E7 19 40 63 1D 77 CE FE BF 9E 45 3D 93 1E
 1C 5B 1F AA A9 3D 70 01 19 DD 84 5D 6F 1D 72 5F
 B0 E2 B1 C8 52 AA 68 5B DC B9 47 2E 13 43 58 37
 A5 9E AA EE B2 3B 2A 58 CF 76 6E CA 08 02 F5 4D
 A1 36 13 E8 FC 1A AA 57 1F 24 39 2C 4B EF 52 CC
 9C 85 9C 66 83 C8 28 F7 4A F9 7D 7E D0 C5 7D 37
 EF A9 6C A2 51 0D 7A 05 34 0F C2 60 8E B8 54 A4
 06 3C F5 29 52 7F A2 1D 46 90 D6 AB 9A B1 15 ED
 89 11 48 9F 90 C5 18 1F 14 4B D9 0D 44 BE D1 96
 04 E1 CC 36 58 1E 56 F1 BA 18 CD 0A F5 8F AB 4B
 EB 38 4C 51 16 28 AF 5B 69 80 3A A6 73 4C 78 A3
 E2 97 FE C9 90 97 EF E9 EC 52 2D E6 D5 03 DB 56
 74 DC 91 CF 57 83 7E B7 3D 69 C5 AC F4 11 9C 09
 70 69 DD 27 4A BB D0 F3 1B F1 D2 05 AC 18 FA 96
 25 E8 76 94 3A 76 7C 02 B4 B9 10 6C A9 71 C9 1A
 D5 86 16 5D 2A 03 E3 E5 D5 B0 2A 8C 4B 59 4E 4F
 10 27 59 89 81 17 CD EF 43 2A CB 73 7B A6 E4 75
 48 92 0A 6F B9 2A 35 14 F8 D6 BF D2 DE 38 CC C9
 F0 D2 82 DE E6 EE 45 A0 7C D4 AB E1 BC D9 A2 F6
 7E 5B 6F F1 0B FF 4A 99 6E 49 FF B9 83 08 5E 3D
 7E CF B0 4F 89 16 79 44 9F 26 50 12 B5 DF 6D 1D
 1E AA 06 30 39 37 B3 7B 1F 83 67 02 2F B3 E1 69
 36 44 15 24 31 E3 01 78 66 38 AA 0D 6F AC B5 A3
 7E DD 28 95 39 9C 22 D0 2B B8 9B 9A 70 C3 52 53
 52 C7 68 A9 16 02 9E EA 3C DB 36 8F 99 EB EE 28
 9B AA B0 C7 45 A2 5D DB 81 6F A9 15 EB 9E 55 0F
 9C A8 CB EC 55 67 F3 3A 01 01 62 73 15 4A 63 47
 E8 38 AC AE 3F 31 79 93 C3 A8 8A A4 8D 1B 5C 04
 FC 05 73 C2 81 82 3D 6B 1E B4 8C 01 1F 62 CE FA
 B7 B3 90 1C 3E BF A2 A9 5F 3E 78 F6 4C 12 A6 83
 1A 3C 4E 00 E0 75 94 63 44 E3 23 B8 0E 78 6D 65
 CA D1 10 3B CE 08 1A A3 1C B2 D7 F5 4F 06 45 90
 2D 44 C3 66 B7 FC DB 6D DF 77 F5 E7 1A 81 5D D1
 20 08 6A 6F A1 28 7B 3B 7E D8 8E AC DC CD E5 7A
 20 37 A8 3C B8 AA 32 1A A8 AD CA A9 CB 20 86 98
 A2 81 F9 50 CF EB 16 F6 04 8E 01 8C BF FF DD 27
 CB 03 BC 38 30 FE 2D 8A 33 D5 5B 69 21 2F A3 0B
 81 EC B5 CE B0 80 0D D5 EC 82 20 8C 3B A4 27 51
 1B 2C 7E 5B 82 3C 77 E5 78 19 6F 4D 3F 03 58 E2
 0F 08 0F 10 B0 78 B5 28 83 05 49 CE 19 89 13 D3
 F4 9A 51 A0 9B 81 76 05 59 2D D1 91 DE 87 C6 82
 25 65 07 D9 A4 D9 21 FD E0 29 00 AA 48 72 7D C8
 C9 BB 02 21 2E D0 94 06 83 6F 97 E8 E3 C2 2F 3E
 B7 A2 A2 82 0E F6 EC 0A 9F 21 0E 79 27 9B 81 A4
 7B EE 07 07 FB AD 2B 47 04 11 E7 83 5D 2E D6 24
 91 21 3D 57 2A 21 C4 29 83 61 C3 44 D5 55 32 EC
 60 63 83 2C 53 7C F4 66 17 17 42 22 07 40 E1 7D
 73 93 FF 6D 5C 8E EC 93 8E A5 50 0F 8E FF E4 EF
 91 72 03 E6 A0 39 D6 3E 2F BF C6 05 6A E4 16 89
 D5 BF 6A 6B 3D 03 E6 88 57 D6 E7 79 08 65 A8 71
 9B 75 BC 64 49 F7 3D D1 19 3A 11 AC 8A 73 20 61
 11 E0 D0 A2 3A 51 6E 7C FA D3 17 35 A1 76 18 A7
 38 50 7B 3E 78 21 31 A7 E4 8D 0F C0 72 3F CB 1B
 83 53 F6 E1 06 5F C5 CE 7D F7 71 B8 3D FD 6E D4
 C4 8B 73 37 0D 93 E3 76 60 24 BB BD BB BE 72 18
 0C D9 1D AB ED A7 9C 6D DF 82 E2 76 E0 41 37 05
 40 A1 21 0C C2 D6 FF B1 56 7C 9B DC 93 B5 15 87
 82 4B 59 EC 47 6C 45 F1 49 A0 D1 4C DF 40 C9 42
 CE 39 63 5D 78 2D AE B7 79 89 7F 47 73 83 94 E4
 13 62 5F 39 F4 63 57 08 9E E4 2F 0B 8D 24 35 B5
 E6 CD 70 3E CD E0 6D 7D 9C 96 EF A3 75 43 B5 60
 29 DA B6 9D 7E 85 73 F6 C8 A0 D0 52 DC DE 78 1C
 C2 26 8B C4 99 05 5D A0 4B AE A1 A1 F7 1C 80 65
 D1 26 5D C3 54 5B E7 A9 35 7D 26 D2 EE BF 43 86
 E5 D1 C1 BA CE CF 80 4F 4E E1 8F 36 8C 60 0A 15
 5A 66 0B F1 FB FF FE FE 27 54 54 34 85 C1 D1 02
 D6 56 62 D3 9E EE CC 92 20 91 0B 5F 60 34 CC 53
 AA 27 33 90 BF 76 7A A8 18 6A AD BB 7D EE 23 C5
 B8 01 E5 1C D0 7D 48 E3 2B B8 F2 B0 C5 B1 E7 B8
 C8 78 F4 66 09 E0 63 15 F6 48 51 B2 5E E0 4C 06
 46 A0 04 10 F7 A0 70 73 7C 6D 1B 35 F9 5F 1B C4
 80 01 5D DB FE 49 8F E7 D9 1B DE C5 94 69 87 29
 D7 E6 35 AA C9 00 63 F9 C1 2D EB 83 6A A9 D8 56
 03 14 CD D3 32 E9 4A 3D 4C B8 58 EE FA 7A BD D4
 79 D9 34 C4 33 A1 72 2A A4 D1 40 49 13 A4 AD 67
 0F 82 C6 5A 3D 7F 55 35 2C 3C 36 59 7B B8 48 3A
 7A AF 1B 8E B2 98 99 85 4A 33 4D 12 9B D4 07 0D
 4E 6F A2 CF F5 72 D5 E4 E6 60 C4 DF 4E 19 2F A6
 FF 78 CB 97 C4 C1 15 9B 56 79 7F 30 47 2E 72 9C
 48 89 BA DE 27 19 76 0E 68 18 DE 33 50 7C 6C 6D
 88 E5 1C 33 4A BC 3C DF 4B DE 49 B3 4F D7 47 62
 28 87 1A 77 1D E4 69 B5 AE 1A 19 40 DC 6A 48 50
 90 A8 D1 BF 13 E7 8E B5 9B F6 92 EB EC 3A 44 21
 C0 14 15 DB DB DB 31 36 28 CB 1A 88 E2 3C 7F 8E
 AC CF 94 60 30 D8 CF 83 C1 DA 35 1B F9 38 15 E0
 97 4C F3 EC D0 FC CA 05 6C F0 9C 15 76 F7 97 0B
 B5 20 FA 5C D8 2B AA 8A A2 92 7A 99 21 B6 35 8D
 98 27 04 1D 94 B9 17 D4 4A E6 CA E0 5A EF 3B B8
 E3 94 2B E2 AE CF EB 6B C1 F3 84 20 FC 54 62 11
 08 B9 C8 58 F9 88 49 1B AA C1 E0 62 C8 EC D8 6E
 2D 3C 80 48 7A 5A DB E0 59 E8 1B A1 7F FD 0A 28
 76 82 A6 6D 30 13 AA 55 91 D5 5A FB 29 66 8C 18
 12 5C CE 7C D2 06 4F 12 16 8D 67 53 76 1F EB 28
 F4 9E 70 5E 32 8A 1B 6D B4 2C 62 94 C1 B6 39 27
 22 2A 4A EC 1E 4A 86 AD EA 9E 80 2A DA 96 9F C0
 F4 AE 3D 95 AE DA F3 35 98 3E 84 18 01 0B 61 B9
 02 36 DD A9 06 78 22 F5 CA 75 B5 85 8C 75 C1 C8
 08 23 25 D1 0F C3 D9 28 9F 4A 30 B2 1C 62 B5 A7
 C6 45 E9 75 74 F6 9F 01 50 7C 73 2A 86 F3 E4 4C
 BE AF 66 E4 05 E1 5B 7A 8F 0D E6 A4 E7 16 C7 FD
 56 F2 57 BB F1 53 9E D4 BF 91 74 AD D5 06 AF 7E
 50 98 D2 E9 CA 28 F8 DF 87 59 5C 5E 92 7C E1 2F
 DA D2 EB B2 8E 1F 8D E2 66 1D F7 B8 07 6B C3 0B
 82 9D D6 CE 9B BE AA 56 83 97 37 B3 54 FB D7 74
 24 42 A2 56 7F 92 9F 9C 5A FD F4 EA D4 87 0E D0
 F3 6B C0 46 81 45 78 03 AA 3D 56 F5 62 86 0F B9
 B9 BF 94 41 E7 0D 77 7C 9C 45 66 AA 04 5A 47 7F
 F0 92 95 C0 E1 31 24 ED 68 C6 AA 58 62 44 7F A5
 68 FD 37 BE E9 98 C0 2E A9 57 84 E6 07 7A DC 5D
 56 86 53 A1 08 DF AD 63 3F 2F 6D 4B 49 94 37 9B
 75 9F 48 53 2E D5 C7 88 09 CE 83 00 9B 04 62 E8
 16 7D DA 1B 4F D4 A0 10 B4 7A FD A4 43 CA 1E BB
 57 B2 3E 09 9C E4 8E C4 44 C2 83 33 0C D0 95 3B
 D6 FB 29 E7 86 A4 CB F0 04 4C 07 B7 9D 23 3B 60
 5A B7 1C E5 B6 22 64 08 98 95 05 5F CD 78 D1 E8
 6F 29 DD 11 E2 F5 9A 22 1F D7 04 2A F2 E7 64 F9
 09 4B F4 DD 89 14 F7 01 F8 E8 0E 4E 6B 36 B3 FF
 D0 72 97 25 BF B5 C2 91 FD FD 8D F9 1F A2 1B 11
 A1 C1 95 DB 40 D0 E6 35 02 C7 39 C8 61 EA 96 DC
 F5 B3 CF 3E E0 2C D0 2C 04 E6 86 BD BF 5E 8E 4F
 90 E0 A5 54 66 56 66 B4 AB 31 EF 36 C3 97 31 56
 B6 50 98 E2 87 F0 3B 0C 94 D5 73 81 E6 58 BD 23
 50 15 98 F3 52 09 76 BD FC 43 CC 17 F8 00 9A 24
 6A 76 66 8E 0E 9C E5 C2 8D AB 01 4B F4 CD 87 DF
 A6 FE 2B 7C 74 9E CC C1 58 0A EA E6 57 C8 AF A9
 0B 97 64 B7 13 81 61 16 95 0D 5B C0 F3 2C 7E 27
 64 54 EB D1 4B 58 17 50 FD 00 C3 2F E5 2C A0 AF
 B6 89 DE 08 3E DC 8A 8B D2 AA 81 E3 C9 08 BD 61
 D4 2E 9E 73 B6 64 96 42 9F 14 A2 14 E4 F6 CE 2D
 88 6E 46 7A 48 BB B8 EE A2 93 53 74 A0 9E BF 98
 25 D9 1C 72 80 32 48 6D 97 1E 2C 1D BC 3F 72 62
 34 85 F5 7A 50 96 70 00 8C BC CB F5 D3 1E 06 AE
 FA 8A E2 C5 3C D7 35 E6 33 95 52 2A A9 ED 16 DF
 F3 DE CE D1 E9 A0 9F DD 5F 16 06 85 45 99 30 03
 F1 70 95 AA 34 5F 83 51 A2 42 6C 90 99 9B CC AE
 80 FE 68 9A B5 95 59 B6 FF 5A 4C 86 75 73 F9 3C
 CE 61 1C 96 5B 27 55 D0 8C 77 64 94 60 EE 84 EF
 98 BC 15 B5 19 B6 C2 7B 40 0D 60 81 2B 32 15 B7
 76 37 69 E1 E2 17 6C F9 6C FE 65 85 84 E2 A9 F9
 2D 6F F1 D2 D7 45 B6 66 D3 09 5D 78 1A 0F DA 9F
 9A 25 DF D0 C6 4F 5B EE DD DB 18 A6 E7 63 08 2C
 85 E6 AC 9B F9 CA A3 D5 D5 96 47 DD 20 DE 9B 68
 2A D1 09 80 68 F8 85 63 89 95 6F 07 3C 21 CB B6
 C7 60 E7 77 29 40 8C AE 0D 58 83 62 4E 4A 99 E9
 A8 21 53 B7 06 97 75 22 56 3D BB F6 E0 12 51 D6
 2C 25 FD 21 7F 61 05 0D 42 D1 1C EA C5 90 EE 68
 1F A2 D5 5B 2A 02 56 3F 73 71 30 DB F2 F3 18 F6
 F9 2E 78 73 FE CB D1 71 4A 56 AE EC 41 D7 01 FB
 A8 51 0B CD 37 BE 92 F6 A7 74 64 B7 72 83 45 74
 05 35 5B 39 BE B0 FD BB 0A 2D 2A 73 83 37 D3 8D
 0B 7B B5 F7 C8 3E A9 C6 CD 33 91 EE 2E C1 92 11
 57 AD 62 05 73 16 96 2E 69 DF 6F 90 C1 99 18 15
 0C D3 F5 6A F3 45 C0 D2 3D A7 7C D4 73 EE 15 F6
 0D FA 68 40 90 47 59 E2 5D 45 FD 37 12 B5 09 79
 D5 E3 4A E0 B8 5E E0 84 E7 0B D3 F9 AD A0 49 ED
 00 16 91 24 4A F8 20 B5 82 32 0D 62 D7 02 1A 2F
 76 89 6A 7C 5F ED 14 C1 9F B5 72 BC D3 44 65 66
 FB 8A F4 8D A5 29 3A E9 CE E5 45 2F 87 6E B6 94
 0A 9C 16 76 F0 70 B4 EA 25 1A 81 75 DA DA 3B 2A
 9B 08 42 06 3F 90 91 3B 57 C9 7C 4A 6F D6 DF 81
 47 C9 54 C3 A5 35 97 DF 98 41 42 4B 97 60 B8 38
 46 6B FD EE 2B DF 1E D1 83 37 5C A6 95 75 7C C2
 8E 91 B9 B9 B9 D8 27 15 8E D0 BC B4 DF 39 EF 45
 95 79 BE FE 04 66 06 4E 66 5C 0D 6F C4 81 79 8D
 C2 52 13 75 7B ED 1D 73 B4 2A C2 14 D3 FA 69 72
 50 E2 F6 10 FC 97 65 9A C4 3F BF AB 37 75 8D 8D
 5E E8 39 44 55 BD 12 78 24 29 CA DD DD 7A A3 F1
 7A 7A 5A BA A0 77 5D 9E 49 0C A3 1A B7 55 16 80
 87 8F 0C 21 04 02 8D F8 D4 14 DB 5E 16 53 F2 42
 1E 53 8A 08 9A C2 1E 93 B2 56 29 F2 85 76 8E D7
 26 64 3F 6B 56 D0 4A 89 C5 E5 46 2A 45 5C D8 35
 80 97 37 43 1C 53 0C 83 BE D7 EF 4F 22 C1 79 99
 BF BF 6A 5A F9 D7 A3 2B 06 CE BB 5C 0E EA 5B DE
 BC B1 FF 10 26 5C 57 5C F9 77 83 7D 0C 9F D5 A7
 A4 57 03 D7 C1 EC FF 33 B4 E3 A5 EA 7B 5F A0 1D
 D1 84 63 02 D2 82 0E B0 4E 50 55 40 E5 CF 07 86
 D2 45 0F 5A 96 FB 82 84 B1 60 C7 AD ED BF CE 11
 AC 05 1B 21 91 8F 15 D7 09 D1 88 0A 82 78 C0 47
 71 93 DA EB AB 62 C7 57 BB CE D4 4A 3F 38 93 B8
 62 14 5D C8 55 A3 17 A4 FC 5D ED B9 05 D1 28 74
 02 84 3E 0D 22 19 D1 C7 0B 3C 24 2A EA AA A3 84
 27 44 34 D2 FA F0 EF 15 BE D5 D7 71 D5 D4 1D A3
 0E F9 08 A1 75 35 C4 37 4D 18 F2 C6 02 E9 F8 F7
 84 E8 CC 46 ED 17 F1 E5 8B 01 10 28 76 4D 48 63
 42 DF 1D 7A 30 A7 FC 0D 1F 7C 35 98 02 B0 34 82
 26 71 AC CA 9B FA 3E 99 37 25 0E C5 7B FB EC 1D
 FE F8 2D D4 09 C8 4B 2A 8A EC 37 28 95 69 53 FF
 F8 C4 E1 B8 5A 48 6D B5 00 88 26 FF 2F 59 5C 3E
 25 B0 4A ED E8 03 F8 CA FD DC 7A B4 76 82 98 65
 2E C9 A7 47 1C EA 20 C4 76 D8 50 CD 15 E5 4E 93
 B2 6F 21 87 89 D5 9F CE C4 1D CA 7E EB E2 DB 1C
 C9 CD 03 02 EF D9 A1 E9 0D 34 9D 01 C0 F0 66 45
 C6 89 3F ED 56 67 88 0D 4F DC 80 0D 91 24 4A 3F
 06 6A B6 13 38 81 70 37 FA FF E3 AD 1A C0 9C FA
 C3 BB 05 A4 A3 F2 2A 22 1B 22 CC FF 64 91 DC 8D
 05 1E 6C BF 39 DB 70 55 39 4C D8 F0 6E 31 ED 1B
 15 6C 42 CD 37 74 84 74 88 6B 9A 00 23 47 A9 8A
 0F AA F1 34 CE F3 C9 6A 55 67 9F FA 42 74 BE BD
 64 C2 09 D9 28 85 56 4D 15 25 C1 00 8B BB C4 E6
 B6 37 A5 0D B5 B4 B8 63 21 05 83 4F A0 A9 77 5B
 51 E7 85 30 23 66 52 BC 89 39 A2 C5 BA 2A 9B 31
 1F C7 FD 7A 80 55 FA 99 D1 72 3E 05 50 6E 9D B4
 1C 29 AC 1B 7C 10 8C D0 46 49 4C DB 09 2B 4F E6
 8B 1A 5F 87 C7 9B 20 96 A8 62 AB 6D 56 3D EA DB
 07 D1 2C 73 DC 3A 6D 73 B2 B3 BA 46 08 92 43 2E
 8E 1F C2 8D F2 F4 1C 05 38 28 D8 E3 26 81 58 BB
 CF 10 70 AB 4E F9 3A D4 D9 C0 E1 CB 28 18 1D 13
 CC B1 7B 5C A0 B7 78 28 00 9A 3F CB E0 BA AC 4F
 D1 0F 23 6B 32 4E D2 7A C2 59 E2 BB F3 21 C0 A1
 0E DA 61 C5 1C AD 9E E9 7F 3A AD FE 93 7F 8A 61
 B0 C8 3C 8D 4D D6 B4 06 85 FC 5C CC 14 C4 51 5A
 69 29 8D F6 2A 8D 33 10 79 58 4F 3F 09 27 B4 B7
 50 D0 43 C2 75 B0 17 93 1E 0A D1 2E 58 DB 4E B0
 C2 C8 2B B2 6C BF 1E 6E 03 BE 8C 43 79 5B 35 D4
 00 D6 53 78 98 8A 19 AB 76 25 2A FC 82 86 CF 68
 90 85 B1 09 B6 4C 33 32 28 BF 9B DF 59 DD 9D 9B
 B2 AB 18 EA FF 2E 68 9F 8A 74 3B 69 08 6F 78 8B
 D2 B5 96 40 A3 39 FA 6A 41 81 7A D3 40 69 33 FF
 4D 10 DB 3C 90 58 1C F1 08 1D 40 92 54 CC 0F 81
 3F 31 B2 60 15 85 8C A9 59 DE 97 F2 AE 2E 84 40
 04 AD 6A 65 95 1F 4F 95 BC CC 9A F5 47 68 71 E8
 A4 2B D6 9E CF AC 6C 42 87 DE 12 AE 6F 60 74 84
 DA 58 4B 77 57 B6 B1 36 F7 DD 5C 89 75 A9 B5 F2
 A6 BC 03 9C 13 C2 62 0A B7 A2 E5 4F 81 E1 4E 6D
 38 2E 29 07 2B 57 B6 19 BE 48 5C 08 21 45 D5 CA
 E3 75 B2 DD A7 73 C3 2B 3A E2 CD D6 36 C4 54 B6
 97 02 B4 BB A9 9C 19 8E EC F6 99 7B 2C 86 A9 C0
 40 2E B8 18 0B 85 EF 7D 6F A7 68 7D AC 7E 34 E8
 BA A3 6F 05 35 9B 26 60 72 2E B3 49 F9 9A DF 45
 23 70 4E 71 B5 64 21 28 E8 E9 8D 44 1C E0 1B 3E
 DD 53 F3 DC FE F7 1D 5A 2B FD 0C 0A C0 52 CB FB
 67 3B E0 E5 A5 32 FA 0F 68 FB D3 8F 14 08 8B CF
 79 F4 AD EC 6E 0D D8 66 E2 65 D9 39 F0 38 AE 7F
 44 48 A3 5B 81 58 64 57 06 1F F4 B5 14 87 CF 02
 2C 8E B5 70 45 54 0D F4 69 36 95 8A 8C 1B 97 9D
 72 F0 58 4C 62 69 65 E2 04 0E 9F BE 96 F9 39 DF
 0D 4E 65 1A 56 CA 0A BF 17 8B 64 12 DA E9 33 4D
 06 A2 CF 76 E9 37 F5 8E 31 BF 60 46 66 74 83 C3
 A8 8D 63 25 95 70 CA C6 31 B1 22 91 8A B3 AE 2B
 1A BE 38 CA 26 92 6D 08 4B FD 61 2B 21 3D 7F 61
 EC 2D 8B 13 2D D6 D4 C2 44 B2 11 C7 F6 A4 F5 62
 51 AA A5 C8 C7 9B 33 CE 28 5C F8 E6 2D 8C 9F 7C
 BC 6D DA 5E 10 13 01 FB 54 C1 70 EC 9A CD 4F 2F
 0C FB 9A 17 1D AA BF E1 8A 1D 0D 55 14 19 9B E9
 F2 53 3D 8A D2 79 46 89 A6 3C 10 5A A8 28 16 15
 C9 92 7E 5C 68 4D 85 46 E3 93 71 81 5E FB 89 B1
 C5 FB EC 72 FB C5 F5 2D 69 71 AC 9A 02 FE 6D 8B
 B8 91 F0 EF AD AE D1 B4 63 31 D3 BC 47 E9 B3 77
 03 7B E7 0C FE 47 76 F6 BC 08 6C 3F B9 1C 70 E3
 2B 59 0F 8B F9 39 BB E8 E4 F0 58 67 F5 93 07 16
 36 53 2D 91 F4 32 78 5B DD 4E 37 12 D6 6F 03 6C
 5E BE A8 DE 5A 4E 03 40 BB 47 C7 65 38 0A 2E CD
 9C 2F 1F 91 CE 0C 61 32 DD 3B 87 55 68 DC 5A 3E
 61 D0 CC ED E3 5C E9 72 41 B8 A6 84 F7 00 AD F5
 F9 5E 0F D6 F9 61 2C AF D8 32 51 2E 55 51 6C F3
 03 13 5B 14 5C 7E 2C 13 7D 37 CA 7C 97 C1 F6 1E
 2A B4 9B 41 6C E6 8D 31 09 01 D7 A3 B3 2A 88 37
 35 3D B3 B7 16 A5 89 FA 2D D4 1A F2 C3 01 67 D6
 E9 53 27 61 45 76 BA 15 08 61 93 5D 7F 1A 96 89
 32 C5 C3 C7 D3 26 EF F1 93 E2 FB D3 67 2C C4 E9
 7D EA EB 7A 40 62 B8 28 AA AF 03 5A BD 96 26 89
 01 16 03 26 02 AA C2 D3 31 2E FB 13 CF 3D F9 63
 7A 69 8A 45 DD 51 1D F3 90 1E AE AF 40 E7 23 72
 1F 70 8B BC 29 3A E3 81 CB 35 90 74 79 14 20 D6
 01 76 05 B7 14 D8 56 DD C3 13 FD 65 EC 16 99 29
 9C 7D 53 CA 73 2E 83 20 5F 76 EC 31 9B 06 80 E8
 C8 0F 70 F4 FB A8 2D D8 3D E5 C1 39 C8 8A A6 7C
 DE 6B 95 78 E0 83 14 9D 59 31 9F 58 8B 89 31 28
 F2 EA 3E 49 E5 E7 77 55 43 BF BB 36 15 DA 39 08
 6E C0 CF 91 3F 0E 28 81 13 5B 8E 7F D5 5F 5F DE
 44 9F AA 40 67 D5 C1 92 BB 40 DF 5F 2A 52 39 06
 E1 D6 99 BC FB 1F 75 82 C9 A7 ED 81 E1 93 EF 56
 F2 C1 56 78 68 FE 86 E1 80 0F 48 95 8B 94 96 22
 21 19 FD F3 28 36 73 76 4D B1 4E 91 CA 26 B5 59
 F6 E8 E0 3F F4 E7 28 35 52 94 F4 04 19 0F C3 EA
 97 EF 6D 18 48 EF F7 09 8F F9 75 CC 57 27 D9 6A
 67 E0 41 AA 84 9E CD DC 86 8A 73 10 F0 8B 4B 7C
 38 35 7C D9 87 E6 95 9E 4C 78 A6 75 03 DE 7C 97
 00 A8 EA 88 1F DD E9 4D 24 8A 28 40 9A 95 B3 EB
 BC 61 BC 6B 3B E3 5A A0 B5 44 87 AC E6 A1 5D FC
 B5 18 15 80 B7 29 BF ED DC 52 23 15 51 D3 4F 18
 A6 89 03 77 36 A9 0B 82 DA 63 66 A4 EE A7 62 85
 8D 1D 34 44 70 87 A4 EE 62 44 D0 44 E3 F0 BB 4F
 09 15 CC DD F0 85 88 6C F7 E1 6E B1 4B 6E 78 23
 E1 C8 99 00 C9 84 22 DB F0 91 7E BF 4A 31 E4 A0
 83 44 A5 EC 33 20 7E 16 D9 1A A7 BB 6F 7D 6C 51
 C1 C4 20 19 7E 42 2D DA B6 1A B0 CE D7 E5 58 74
 DE 35 C6 CC 3A 4E EA D9 35 39 2D C1 EF 54 3F 93
 22 04 15 7F 71 CB 07 A0 49 82 56 BE 7F 18 B8 25
 5F 60 EA 2C D8 C9 7C 7C 19 B5 99 60 8A 82 74 E5
 AE A3 EA 10 5F 29 2F 2B 48 2C 29 84 05 3C 7B 64
 56 D7 9F E3 E0 5A 88 18 DD B6 F3 E4 41 B8 76 6D
 3D E5 E1 5A B0 F2 02 09 3B 6A 68 11 46 D2 C1 B6
 A2 FA 62 36 ED B8 50 0C F9 3B 8D 0B 29 A7 0A 26
 D5 71 32 51 FA 25 8F 0E B6 C8 6E C9 A9 F2 2D FD
 40 BE 8A 93 F5 1C 24 4D F3 E2 80 A2 F0 D9 F9 A1
 4E D8 03 04 62 4E CC AB 0C F7 FC 40 9F CE 09 C7
 69 52 6E 83 32 4F E6 35 3D 45 E9 10 33 05 EA 1A
 82 80 80 75 44 3A F3 66 77 A7 2D 2D D2 E3 F4 C4
 FC BE BA B4 18 E3 B4 E2 70 2F CC 41 2F 41 DB 44
 79 47 55 06 E3 24 33 68 09 F9 DD AB 81 00 52 9A
 C9 5B FF 54 2D 55 38 BC 3B 19 18 0E E2 30 F9 56
 DD BF D5 79 59 1C C6 5E 72 E3 D4 B8 35 2E 43 E9
 A7 27 B0 FB EE B9 EA 81 95 21 D4 F5 58 85 B1 2D
 B6 44 BE 68 78 F4 79 22 8C AC 56 0B 3D 74 8E ED
 E1 16 2F 3D 78 01 9C A3 09 B8 FF 0C E2 F6 3B BB
 49 F6 54 74 8E 24 6F C4 F4 FC 37 7E A1 C4 72 C0
 14 38 77 52 07 E5 56 61 10 00 19 7A 1C 4C FB D0
 E2 35 D0 5E B9 58 33 31 A8 BD D4 A0 7F AD 1E E2
 7C 3A E9 BC 32 80 42 75 B1 B7 2F F7 C7 30 BE 37
 7F 47 21 5E 22 D9 E5 55 57 79 2E B3 B3 67 5A 81
 6E BE A3 85 3D 28 7D 29 28 80 FC 3E 99 85 66 4D
 1D 92 20 12 E7 C2 39 A0 BE D3 04 AE 63 C5 99 AB
 DA 4E C8 F8 7D 84 47 E0 4E 89 9A CB 37 5B 03 74
 B2 11 BA 6C 1F ED 0E 92 6A 16 75 66 80 65 B7 F7
 E4 34 77 D5 2D 22 7C 83 23 A4 94 53 7C 48 29 C2
 03 14 7A 67 F4 82 58 83 03 C0 1E 9D 41 2B 78 22
 DC A4 93 C3 29 65 B7 C6 DB 2F B3 FC A8 FB 8A 7D
 D4 C0 CE 06 88 4D 8A AF 27 FB 83 21 22 20 0E 05
 E5 FC 31 EA A1 3A 61 B0 7D D6 E2 17 36 5E 81 4D
 7F 42 5E 65 21 1A 44 8F 2E DE 5D 7F 3C 62 FF 75
 58 D2 C5 6B CE 91 94 9A EE 25 9F C3 8C DD E6 1C
 A3 A1 78 80 00 92 3C 24 EF DA 6A 61 CB B6 6C 54
 95 34 FC CA 1F 8C 6F 8F 66 34 56 5F 30 00 A6 DE
 94 E2 CD C9 B3 C8 62 46 00 1E 61 52 4B F0 CD 0D
 DB FF BD 71 EF 2C 31 16 99 D3 1B 8E 41 2B AF 70
 7B FE F6 E1 93 24 91 90 34 73 E1 06 2F EB 2B 0B
 FE F7 38 6E 4E 93 1E 13 A0 95 CB AC 04 91 02 6E
 F7 4B 0B D7 F9 88 A2 96 52 11 77 DB FE 5C B9 28
 4B 6C 50 37 CE 18 5A FB EC 7B 61 83 5B 2A 72 44
 91 86 AC 7C 3C 5E F4 B1 72 6E 32 51 AF F7 CD C6
 A2 F7 B6 D3 AB F4 6D 8C 22 04 FE 58 C9 BA 9A 46
 45 3A E4 40 8F B5 19 95 3F 83 2C 41 0D B9 39 61
 60 B8 DD 9C 3D CC B4 63 A7 EA 5F C1 B5 FC 1B BD
 6A 79 6E BE 04 38 82 73 4F 68 3D 54 DC B1 EA 1C
 7F 33 53 55 AB 3A 0E 3C A1 5B F1 03 C8 B1 3F AA
 39 C9 0F 4C FA 5B 54 07 42 B1 91 85 25 FE 04 A4
 F2 61 7A 21 C2 24 12 D9 CC AF 4D CB D2 9C FA 61
 79 BC CD 97 B1 C2 DE 40 64 99 2A 5E CD 61 98 25
 93 EE 50 7C A6 D9 BB CC 56 5D D7 EF 1D 28 6B 7D
 F6 02 B8 3D 0A 3F 98 1E 55 0F 8C 8B 1A C9 46 92
 57 01 FE 99 5D 7D 2D 6F 0D E6 86 EB 43 B5 2A EB
 D4 DE DA FA C6 16 9F A1 4D 69 F5 B7 95 EB 54 59
 34 2B B2 D1 CC AD D6 AD 28 0A B6 45 91 F6 EC B6
 60 65 D4 EE F2 64 62 F1 FC 65 C3 34 5F B2 F6 E1
 CA 66 F8 30 D9 E5 11 39 17 27 72 00 48 14 1D 84
 34 95 D5 10 FA 9F AC EB B5 AE 71 36 69 E4 FA 2D
 16 64 52 F2 95 F1 26 05 71 41 95 A0 1C D0 B0 E4
 AB D3 FC B8 4A 45 00 13 1A 4D AC 59 C9 95 40 6A
 11 84 AF 36 43 A5 D9 3A 55 4E 9C 82 67 98 4A CD
 E8 05 6E 33 82 7C FE 9C 4B 45 00 B6 3D F1 0C 4D
 76 FD C7 6E 06 06 8E 22 39 B2 9C 35 0C 47 5B 89
 28 7A E7 4F 67 FB 3B EF 2B 16 C5 BA B0 04 0C 34
 32 5B D5 55 47 C2 82 0E D9 04 BC 05 62 17 15 5E
 55 93 EC 67 42 BB 4F 1D 09 E0 0F BD 61 25 57 90
 D7 D7 50 9F 8C CE 8F 28 CD 16 3B B5 69 3B 84 31
 B5 A6 F3 5D 79 EE F3 6C 4A 7F D7 02 41 05 CA 75
 DC 28 A9 4A 5A 0F 37 5F 99 F9 F3 5B 52 04 EE 10
 2E F7 BE 36 74 9C DA 09 08 23 91 32 1C BE F1 2A
 C4 B3 A4 BD 48 B2 22 54 F2 E8 58 08 21 BF 52 6D
 D0 44 95 87 ED 85 A0 2D AE DD 05 48 DE 78 FD BB
 9A F0 08 3A F5 26 C7 CC C8 5E 8F D2 50 01 33 3A
 E1 77 5E F1 3A FE 7C A5 C1 3E D7 7E 39 E6 37 96
 A7 4B 62 7E D2 15 E1 51 8F EE 7F C5 47 94 A8 48
 31 24 0B 35 0D 98 DE 00 51 1D D5 99 17 FD 09 18
 B6 73 A7 CD 93 A2 66 D4 2A 3E D2 29 49 03 84 AC
 9F 4A 62 2A F4 F8 B5 26 CE 55 A1 95 22 24 AC 44
 32 DA 37 59 5D B7 6F DF B1 17 DA 89 4D 53 F7 23
 C7 C9 C4 43 46 67 4F 03 1E BB 03 AE 76 D3 65 CB
 FA B7 F8 80 AC B3 48 00 CD FA 9D C2 E2 55 90 69
 2F A5 94 44 F6 72 37 0D 52 1C 50 AC 23 41 E3 88
 4C E1 C6 B8 1F 7B A9 B9 22 9C 00 F9 97 CA 43 6C
 40 0D 7A CB 31 35 1A B7 05 2D 22 F5 92 C6 20 D1
 25 C8 5D 94 9F 6B 67 12 FC 4B 69 05 44 F8 65 1F
 AB 38 1B 2C 45 88 1D B2 24 4F EA FC FB BB C5 C5
 78 21 47 D5 2B 39 2F AD 90 BC 7E 81 43 44 AD 59
 D6 4C 48 DB A1 DB DE 72 F1 3F C6 A1 40 34 4F 75
 B5 6D 92 1D 16 B1 EB C3 71 D8 3B 3D 47 84 76 72
 B4 AF 1D ED 97 0C 4B BB 67 3F A3 63 5D E9 8C B1
 3C C8 01 EC 97 B2 73 42 93 BB 1C 02 10 B9 70 92
 24 B6 B5 62 0F 78 20 6C F0 AF 63 97 A1 22 0E 59
 95 2D A2 AD 11 46 26 F1 8B 9D E9 C7 F9 65 8B DF
 19 8F 98 FA 50 8F 00 E3 A1 DE C2 DC 36 CC 2D FE
 17 BB 02 62 C5 1C B8 7C 81 24 B5 3C E7 8F A1 51
 B6 9C 6F CC 33 2C 4B C8 BC 84 5F D3 00 11 0A 2F
 4B 17 11 69 17 D6 01 E8 68 1E 3E FA 99 C1 E9 9D
 64 F3 14 A6 F8 B9 A2 40 E0 79 18 D6 87 31 FD 41
 3C A2 9E 45 7D D0 CE B7 D7 7F 82 45 89 06 46 6C
 EB AE BE B2 56 5A 72 4F 52 02 FC B5 14 BE 9D F9
 4D 5F A6 33 E2 4C 70 12 08 F9 A2 E4 F8 D3 22 63
 C7 27 A9 08 32 54 09 31 7C DB 76 B4 C8 5C 3B F6
 09 E5 D1 22 62 4B EF 4D F7 29 0C 1E FC E8 89 86
 3E 4F B2 B4 77 D4 65 EC 85 F0 8A 7E 21 41 D7 4C
 EE C6 FF 39 43 B9 BC 95 4A AB 2C 75 D1 9A 59 8D
 17 C3 C5 0B 66 E3 21 14 E7 49 56 B5 1F 14 3E D9
 5D 77 B1 0E 5E F0 2B 7E 5B BA 91 E3 C2 63 4B 8A
 24 67 4A 8C 0E 39 9D FE D9 37 97 D4 D1 4B 28 C9
 BE F2 49 9B BF 83 9B DC 23 F0 70 5E 40 5E 9B 5D
 60 DE 9D AE D3 80 D2 2F 67 B6 18 A4 08 13 10 25
 16 12 73 62 47 10 AD BC BC 13 35 93 E3 18 6D 7A
 CB EC 71 D1 19 DB 27 66 A6 95 F8 53 5B 6D 36 B2
 8F 9F DD B8 4E 2A 0E 25 30 56 E4 41 CC 56 9C C3
 45 06 F2 02 E3 90 E2 7B D0 B4 07 AF BC 2B 9C 14
 DF 27 61 2C D9 98 C3 A0 71 05 CD 41 21 F7 70 05
 57 8A 71 5C 58 94 A7 2D 49 F2 17 34 E7 E5 FF 71
 F5 BD 62 AC 72 5A FB 2B 20 12 B9 7B AF 70 46 FE
 42 91 78 1B BE 3B 92 5A 38 25 A8 A8 F1 D0 7E 76
 AE 01 74 79 65 E5 D6 0B 76 BC 7B E7 26 92 98 EF
 D1 72 BC 4A 69 0B 79 FE 8B FD 99 12 63 8B 57 3F
 78 12 DA 67 4E 57 28 FE 0F C7 9B 8B CC 41 36 FC
 01 DC 4E DB 96 5E 97 54 1D 09 12 8A 67 3E 28 E1
 88 FF 95 76 92 78 42 C8 25 34 F7 3E 8B 37 E8 06
 42 F4 F9 07 88 56 41 EB 90 73 8E EF 15 DC AF E3
 AC D9 1D EF 43 B2 BA 23 3C E7 A3 71 C6 A1 74 2B
 21 4E B3 F9 E8 ED 25 12 D2 06 AE F3 31 5D 01 42
 AE 18 E8 7C 57 A5 7F 3A F7 5C 42 BC CC 50 63 60
 BB 4E CB 9F AA 05 6B F0 24 5B D4 2E 92 08 BE D4
 4E 2A 2D 0B 9B 67 B4 CD 5D 5B 9B 71 67 8C 2D 7B
 FC B1 14 82 D4 1E 65 8C 75 F8 13 AE F2 7D 73 AB
 5A 41 42 7C ED F3 24 19 73 DF 3F 7E AF B2 EA 23
 C7 F3 3C BB FA 87 BD BE 5A E9 EE F6 0B 83 FF FF
 48 AA 75 C5 C0 C3 7F 5C 47 15 4F 20 EA 0E 51 E5
 1F 9B 00 AC A8 8B E9 06 B9 05 2B BA 94 26 8B E2
 E1 D5 53 3E 13 39 F2 1C 35 1A DC 4F 02 11 D4 94
 40 4A 02 C8 21 BC 1F 3C E8 8D 22 6C 8C 2C B4 94
 AF EF C5 87 6D C9 A5 DF DC 71 05 9F A8 2C 51 33
 71 7E 4C C7 67 FD F7 2C 77 CF 4D FD 78 71 82 73
 3A 77 71 03 5C ED 1C 01 1E EF 58 43 D5 30 46 62
 F4 11 FE EF BA 4F 18 C9 87 90 95 32 89 0D 61 45
 C6 73 A4 B5 6E 85 99 95 3F 26 04 42 9C 56 86 4F
 9E 43 07 F8 A0 50 29 48 5F B1 CF 29 6E A2 BA 16
 E3 56 CB 1C 6E D1 A4 51 B6 1B DF 51 64 F9 0F 73
 15 39 70 D7 74 06 04 2E E7 65 7A C0 BC 6A 43 CC
 45 A2 0A 65 98 C2 05 FB 66 E5 0B BE F2 6B B2 CC
 28 C3 F1 13 E5 A5 96 73 32 06 D9 CC E6 59 75 F4
 21 4B 2D 50 B4 ED 34 C8 3C 23 8F 14 2D AC 71 5B
 5F 17 8C 81 11 FB EF 52 44 69 81 A1 07 86 D1 0C
 20 21 39 75 D3 04 D9 AC 1A CE C1 36 04 0D A4 11
 6F 02 7C C8 A6 AE 6F 70 73 4D BE 89 84 99 BB D6
 3F 52 DF DB 5E 1A F6 DE 97 19 9D A1 2D 14 1E 62
 72 6E 9E 19 14 8F 0F 05 98 EC 36 8B F2 01 AD 28
 59 53 10 F6 F1 D1 FD 4F 0A 11 ED ED 4B 36 64 9B
 ED A3 2D 6D 3C FB D3 5C 7D 55 F2 56 78 67 3D 29
 B6 41 C3 68 62 8A 7B 32 11 79 1D 0F 0A C4 2E E9
 92 2F B6 C0 8F EC BD 00 F8 63 28 2B AE D7 08 C9
 39 B2 45 71 FB 30 54 63 FB 73 4E 55 8D 64 8D FE
 84 F3 F9 0A 16 A2 F7 2C 2D 9E 7A 88 DA 23 48 95
 77 3D F4 33 DB 03 71 F6 8A 77 14 24 1B C1 24 05
 F5 1C 41 85 C1 9F F0 04 2C 6A 7F A8 AE 15 DF CE
 0D 8B 2B DB CE 01 1E 31 DD 2B CB 37 3A 8D 5A EE
 23 F5 14 71 BB 60 F1 23 46 AF 61 62 43 88 46 95
 BD CC 99 7C 62 17 8B 12 4B 7A 8E B2 72 67 AB C6
 D5 C4 41 8E 19 DB 47 05 71 48 51 71 8B F4 4B AC
 E1 4C BC 24 BC 12 01 29 F8 37 32 80 1E 2C F0 64
 14 25 44 5B 72 49 7B 23 8B 3D 81 4C 70 21 60 3D
 86 6B 5F 90 44 19 C5 D1 46 82 F4 F1 06 79 43 5A
 E1 D3 2E A2 2A CA 3E DF 5A 06 51 69 E8 66 A2 72
 BC C7 81 91 F1 53 FA DA 64 66 D4 FB 86 DC 49 8B
 A3 D2 F3 70 5A 72 F1 69 55 10 C0 04 FE 36 2C B1
 B6 20 0D BB 60 37 DC 48 96 D4 B7 B9 FC CC 2D 1F
 A1 61 9F 70 B6 EA 27 C9 2B BA 40 CB B8 41 C8 AB
 30 A7 B0 EE 8E 03 68 D7 14 F0 0B C6 03 B8 46 CD
 50 2E AA 9A 9A 66 59 A1 B5 25 67 88 31 04 0E 28
 C4 94 38 93 4A 5A 80 F1 18 27 D1 F8 C8 6A E8 5B
 53 B6 57 FF DE 16 A2 40 2C 7D 6D 47 1B B3 BE 59
 62 10 09 A5 C8 77 B5 06 EE 03 DA 3B D0 A4 23 C0
 40 0B F5 15 FD D1 61 C7 14 BE 98 38 EC 06 DC A0
 E0 26 37 44 AF 7D A3 4A 97 22 5C 22 86 A0 28 88
 E1 C6 24 4B B3 B4 17 2F 80 49 4D B0 21 05 B5 98
 0A E4 CB EA 70 3B F0 4A 3A FE 9F CC 35 7B 3E 8B
 5A AF 04 91 AC B2 7A AD DF 48 B0 02 7A 14 F0 A2
 69 FF 98 31 FE 06 08 9B DB 49 54 78 AF FB 24 2F
 31 8F E8 FE CE D4 CA 55 EF 4F 8A A3 43 FD F5 BE
 8D 55 11 26 4C 69 6F 83 83 2E 64 A2 EA 7C 4C F4
 60 B5 66 BB F8 C1 39 B6 7A 34 64 A0 DC 7C 20 4D
 B6 90 B9 D9 F8 C7 36 0E 5D E6 F3 93 F7 75 90 6F
 73 D9 E3 45 DA 45 B1 BE 6C 28 9E 93 8C 43 EB EB
 EB 64 6E 48 F9 F3 7F E0 0E 35 86 5F AB DA 56 2B
 62 7F 0B A6 79 AB E2 81 E2 9A 90 81 50 D8 92 0D
 7E FB BA 9C 16 A2 B8 8E 97 D1 48 A6 B7 53 4D 7F
 7B 3E AD 44 4D A4 81 84 50 B2 FA F9 C6 5A 47 3D
 EC 39 FD 9E F1 E0 4E F5 6E 1B 98 CB E1 27 95 65
 2E 46 AD 9C C9 43 7F 0E D7 B3 00 87 DA 64 56 C1
 9E 7F 7F 93 8A 10 CF 12 C3 E9 52 73 17 13 6A 3C
 9D 7C 4F 96 1B 8A 2F 05 D3 9D C4 68 F9 DB 11 1D
 9A 65 02 FB 2C 82 B3 91 D7 5A 84 EB C7 B5 10 C1
 A7 67 15 08 E4 B4 04 45 02 A2 63 A8 92 CE F9 16
 EE D9 28 1A 28 F2 1F AB C6 5C DE 4E D5 39 65 19
 54 BE 6A C0 6D 62 B0 CE D4 46 26 CB 71 7A 5A 7B
 C7 1F 68 81 71 B0 9E 10 58 1B 30 CE 19 F2 3F C6
 EE B0 BE E7 BC 7B 66 74 A8 23 3E 2F 25 D0 89 AB
 89 D7 E9 AD D2 FA 68 B5 BD 13 A2 63 D7 C0 A9 22
 5F D3 16 EC 40 CC DD F5 41 CE B1 81 56 97 F6 3D
 05 BD 17 26 F0 D3 E5 F2 3D 90 5E 42 98 45 8B 06
 A5 B9 84 31 0E FB 1B 8A AD 00 86 7C 13 26 15 F5
 7B 4B BC 13 A2 93 3A 67 FA A5 44 49 8A 4C C9 C8
 84 F6 29 BE 0D C3 F7 A0 82 6E D0 05 2A 03 9B 45
 EA D0 DD 5A A3 C5 CF A6 DA 6E CF 94 60 1C F9 14
 C9 9A 8B 85 3E 3C 74 0E 73 B5 6C C9 5D 4F 47 F1
 1C 01 1D 6C 2D EB 63 A4 37 F4 09 CB 27 0F B4 53
 E4 0B C7 6A 85 9A 81 D2 CF 6F 08 51 A5 CE 73 4F
 2E 1F 63 E3 AD 59 A3 56 D1 4A 15 E3 DF 36 0A E2
 7E 83 E8 FF 09 7F D9 E9 6B 24 AC B3 5C 64 28 0A
 72 AE 26 73 C0 59 B7 BD 88 5C 47 98 CC D5 48 72
 98 BE B4 65 9D 63 A9 CD 13 C5 8A B7 94 AE B6 EC
 17 60 9F 04 79 44 69 D4 14 93 EE 44 29 C4 1E 33
 D2 46 A2 49 49 25 65 E2 35 7F 90 43 FC EF CC F5
 05 77 55 00 AD B4 AD 94 0F 72 0F 3F 8D 86 27 0E
 33 9E 83 8A C3 96 3B 50 A6 68 D8 7A 9D A9 9A 44
 15 55 51 B6 9D C7 39 9D 68 FC 9E F3 9B B9 61 88
 19 DE 17 25 95 EE C1 D1 58 07 47 44 77 B3 47 F6
 DC 58 41 4E 83 6E A2 E5 A4 98 46 57 02 03 6A 9B
 4B 06 47 80 7F F5 93 0E 6B 8E 28 42 8A AF 4C F4
 32 B5 6B 86 20 F2 09 19 84 8E 7E 1B 02 2E C3 27
 91 46 17 D3 A8 B6 83 A3 47 6E 71 11 37 91 B1 8C
 16 E2 CC 8B 2A 1B DC CC 55 FB DC 93 29 DB 3E 50
 09 DE 3E F6 1D 05 D2 DB E1 7D 0E E2 C4 FC CA 29
 F2 19 05 78 7B 0E EB 46 EA E5 15 29 86 49 C8 00
 E9 36 31 69 43 C1 17 E0 E8 1B 7A 52 B7 C4 58 8B
 F5 6E 42 9B 64 4C E2 8C 6B 2D 07 70 3D B1 D4 E2
 08 54 E7 23 27 E4 00 57 1F B0 17 68 6D 62 C1 B0
 6F 4F 91 7E 58 81 B8 94 6C E0 B7 9E 59 7E E6 32
 1E C1 ED BC 05 E8 C0 5A 22 ED 83 1D 71 0F D7 1B
 C6 BF 74 35 D4 FE 5D AE 4E EF 96 1B 48 27 AC 4D
 01 E5 C1 A3 CC DE 5E 33 A8 E0 36 1B 8B 8C EE D7
 96 43 7B 8C 8D D2 7F C8 F9 38 91 05 6A 9E 33 97
 88 BA 61 32 5F 2E 4A 01 69 60 51 4F E5 FB 21 B9
 AD F8 09 B3 64 0F 0D A3 91 5B 27 05 63 98 A8 43
 CE AF D3 87 0D B3 96 49 B5 7D 62 B6 1E 87 BA CA
 08 E5 43 48 EE B3 AB FB BB 23 E6 2F 22 C3 F3 AA
 42 D1 8C 50 0A AA 50 3B 6F 0C 56 5F E9 7C 5F 84
 D6 43 C2 96 14 AF 5C CA EE 6E 16 78 C7 9F D9 A5
 E3 E3 93 41 11 1E 37 CB 40 52 00 48 19 85 95 1A
 00 0A FB 72 05 F1 44 B3 90 87 D1 13 27 65 09 19
 26 C5 DA 31 A0 9D 99 30 AD 48 68 EA 8A 2F 25 4C
 CD DE D8 E6 5E 42 FD 04 C5 22 87 21 2A 5A 6F 6E
 65 88 DF 17 68 D3 CA 62 14 92 60 9E E7 3B 14 66
 F8 34 07 9C 8C 5B 8A 05 15 12 EB 81 67 D0 3C F4
 0F BF 56 1D 76 69 43 39 43 89 4F EF B3 AC CF 7D
 79 A9 10 29 84 A6 98 EB 84 50 1F E1 7F A0 7D E9
 7B 95 90 D3 CC E4 11 3D B7 11 48 11 81 B1 ED 3F
 66 B7 F3 98 05 26 B3 1E E2 33 22 1D AE E2 11 5D
 AD E3 EC 0E 99 EB F7 FE B5 42 A0 A5 0F 58 B9 1A
 DB 97 82 2E 09 71 5D 9F 7D 0A BF 7F 59 9C 77 FC
 8E 9D 90 04 DB F8 25 DB 09 2E 65 35 4B 87 D3 02
 0E E0 5B F8 38 F4 03 D3 3A 81 58 8C 8D 69 CC E0
 57 83 4B 6E 5C 7D FA 77 7A 25 10 AD 03 4D B6 61
 63 31 EE 70 F8 B4 C5 9B 78 A8 83 EA E1 B8 D0 A8
 DD 8B 48 C9 94 6A 74 75 25 DE 10 1A 12 D0 C9 CF
 1F 5F CE 29 AF A9 A0 A9 C5 7A 40 4B EB 9A D2 2B
 AF BB 54 C5 51 E7 E4 EB BD AD 71 56 98 93 5A FC
 68 DC 46 2C 01 32 AC 1B F5 96 72 F4 71 81 E6 8B
 6F 92 C1 B3 05 56 F8 BC 69 07 35 2A 1E 94 03 C6
 4C C0 CF 6D 5C C4 01 00 39 B8 73 46 E7 90 10 FC
 A1 0F 65 E7 37 10 58 03 4A D0 2E 3C 34 29 2A A2
 71 F6 27 D1 CB 5F 5F 05 70 1E 53 D7 11 22 AB 4B
 E1 16 D3 D7 9B 07 3F 7C FC C0 D7 73 E1 DB 4D EC
 D0 D9 79 C7 8A 26 46 20 75 36 DD 58 6B 0F 39 F3
 36 B1 BA 9B 58 F7 28 20 5C 3F CA 96 44 24 21 0F
 BA C6 2D A7 92 B2 3E 5E C5 2A E8 8B 77 4A 50 1B
 E7 B6 84 E5 8F E5 07 9F 54 EF 80 91 3D 94 26 A7
 7B 02 18 57 65 B6 E9 62 79 B6 D4 6A 66 89 D4 46
 60 98 A7 7E 5F 98 D3 1E 9B 41 30 2C 14 05 35 6F
 3D 5C FD 3F 20 E4 4A DF 93 7B B1 B7 56 0A 87 58
 48 84 FB 26 67 EA 5B E8 8C 15 6E 56 E7 4D 20 C3
 01 E1 0E 1D A2 89 36 15 D5 E5 60 E6 5F 05 47 F4
 4A 6F BD F3 89 5A 60 2A 15 45 9D 89 4D C4 CD 28
 1C 31 EE 49 8A 4A 34 FB 16 7F 30 9A BA 32 94 0B
 91 6F 54 2F 5D C6 64 57 F8 61 D9 48 24 AE 06 57
 B0 40 FD B0 AA CF 38 7D 74 E1 EA A5 1E B5 27 86
 27 7A 19 29 F5 D3 37 4F 99 D4 0D 37 A8 02 43 C1
 F3 B4 47 FA 6A 67 CC 34 D9 E1 4B 31 93 CC 4B 89
 9C 32 8F 42 B7 46 9F 6B 53 20 58 D1 93 87 CF 0A
 D0 31 57 19 7C B8 9D 01 9A CD 5E 99 23 1B 67 73
 38 45 20 C6 C0 6F CF 18 08 2A 96 77 52 69 B7 0A
 4B 2C 04 78 5B 49 6B C1 44 69 B0 20 42 F7 A2 04
 DB FD 62 30 5E CC D1 8F 4B C8 14 60 05 DE A7 DD
 D0 61 C4 C7 93 62 71 D6 E3 08 9F 09 85 1D 17 A8
 FA F1 46 89 DD 21 49 B6 00 42 8A 6D E1 3C C7 48
 BE 3E 4F DD 4E 0F 8D B6 B2 8B 05 9B 47 6D D7 4E
 CD 26 10 5B B0 24 24 8F 2B 9E 48 84 4F 20 32 A4
 1E 16 26 BA 1F 7E 7B 54 49 A8 A4 A0 E0 64 20 B7
 03 38 70 DE 36 92 B6 48 94 9E 56 E9 75 80 F5 01
 E2 9E 50 13 CD 12 2D 22 10 1C 73 BC 0C 51 14 61
 E5 DC B6 A5 17 46 08 08 D5 AB 58 7F C1 97 FB E1
 A4 FE 77 55 A3 71 3E 88 A0 2E BD A2 AA C8 BD 97
 69 A7 53 8E A7 41 A9 FA 65 38 C2 8A 82 F0 3F D5
 66 80 69 15 64 A1 02 FE D2 F7 64 6B 34 7A 87 35
 1B EC 25 3F 7C A3 99 E0 DD C3 68 CC 2A E3 4B 83
 FF 3B DD A8 8E 90 57 F8 8A 96 09 76 9D 58 12 3E
 FB 72 E2 A9 E4 C4 60 B6 B2 F5 57 FA 30 BA 08 E2
 18 73 5B FC 78 D6 93 DA 6E 1C CA 46 17 76 12 A9
 62 C1 C9 7A 89 1F 1E 5C 77 A7 69 AB 79 12 90 5A
 BC 79 F4 99 82 F7 93 91 F8 18 EA 37 F1 9B 7B 68
 33 C1 29 9B 37 A4 6D 21 8C 65 9B DA D8 A6 08 A8
 89 B4 04 22 63 F6 0C 66 0D 75 C7 18 2A DD 1D 63
 D6 61 DE BE 72 D0 8F A3 A7 13 50 35 BD A6 CF 2D
 7C F4 0E 08 3E FF 0E F5 6D 15 52 32 B6 65 83 F2
 11 99 9E 7E 3C 75 3D 13 30 D8 B4 F6 19 89 9A 8D
 6C D9 20 62 9B 5A 56 DA F7 5B 43 AF 1E 33 CB 14
 E4 50 CD 6F 9B F4 BC E0 5F 60 FD 4B 77 59 CD 0E
 F2 2D 26 A9 89 E2 B7 B7 BA 1F 25 8A 6E 83 03 62
 A1 A2 7E 58 48 4A B5 1D C0 8C D8 22 19 D5 D3 F8
 73 5F 86 F8 B2 25 BA 62 B6 84 55 33 63 D5 46 38
 FE CE E5 82 6C 6C B8 8E 27 A9 C0 8A 36 B5 27 9D
 12 8A E5 1C B2 79 45 42 41 A6 D9 65 EF E0 FE 74
 B4 3F EC AC 0A C4 1C F3 39 8E 6F 79 06 CF 35 54
 C9 6D 35 74 4A B9 82 0E CA 57 24 32 80 58 02 EF
 E0 62 8D 09 91 96 5B EC F9 09 18 A1 FE DF 5E 5E
 A6 67 1E B1 27 00 40 31 3C 22 B4 EC 17 B6 21 34
 20 1B D2 4E 19 FB 7A 91 64 30 8A B4 3C F9 35 C1
 DA 69 D5 11 30 4D 36 B3 10 C7 5A BC 9E 2F E0 65
 90 9C 83 3E 60 E5 F0 6E 02 6F AE ED 13 A0 DA 6F
 2A 6C 77 2E 36 8F 99 25 A2 23 7A 93 CC 19 6E B9
 1F 5A D9 6D F3 68 28 A1 D4 DF ED 28 3D DC 8E 5D
 D3 9D 52 50 00 3B 90 7A 37 A0 66 03 ED 15 A3 2A
 82 33 DC 8F AA 80 84 B6 D3 34 B7 7A 6B EA 3C CE
 CF F8 39 B5 58 8B 5C DE F2 A3 96 3C 30 40 68 13
 3A 41 71 1C AB C7 21 7A 47 F5 1E F5 55 5E B7 11
 46 D9 06 B6 C1 37 D4 43 63 D6 DF 9C FE D7 B3 1C
 B7 01 12 77 B8 44 5C 5D 79 75 46 E1 F4 DB A4 96
 7C 4A A4 EC A0 1D E9 41 1C 1C 32 3D FC 31 69 78
 94 0A 54 CB 21 29 98 51 B3 5A A8 4A 15 16 76 61
 BB A3 A5 1E 4F 4D C4 78 B4 78 08 F6 4B F1 92 AA
 4A C0 82 0E 33 37 21 6B 02 5F A3 BB 02 53 0D 39
 F5 1C CA 1B 26 48 33 B0 AE A8 DD 67 B4 CA 1C 93
 7C 47 B0 74 21 20 83 C4 3F CF 37 55 FC D3 84 9A
 04 75 6C B8 CF C2 5A 91 9E FE A6 E3 5D 71 04 25
 D0 E9 72 8D 14 99 F0 55 87 2F 0E 1D 17 39 D8 69
 ED CF FD 92 F6 99 23 84 B1 63 80 CD 81 2D F1 84
 35 83 D1 32 09 05 71 12 5C 8D 40 47 AF 44 5D 05
 18 2E BA F9 B8 64 EE E0 FC 3E EA 11 94 EC 3A D7
 8B D3 56 6E 2F 04 68 91 8B 2C 82 EE D6 A7 50 76
 28 43 5A 5E 6A D5 1A ED 15 AA 36 C5 7B 1D 1D 8A
 DF 98 A3 EB A9 30 EC 0B 66 51 7D 1F CD 83 4D 39
 55 A2 A6 03 6A BF 32 31 35 AA B9 A1 6D 60 DB 7D
 38 3A F4 70 3A 62 BF A7 76 41 63 68 54 25 E4 C7
 F4 C0 4E E0 56 FF AE E0 D3 8E FF 0A 36 05 3A A6
 CB D1 9C 15 A8 EE E0 88 40 F5 FB 1D AC 06 E2 63
 3A 0D 73 27 59 FB 41 33 69 14 D0 FB CE 11 51 1D
 B0 B4 73 93 20 86 98 EE 71 13 78 09 D7 88 CF 0A
 A2 99 D4 07 2B EE 20 06 45 36 67 B4 80 8D F5 6A
 F4 15 09 F6 77 0F E3 1B 92 28 65 1B 38 20 3D 1C
 29 C2 32 BB 5F C2 A5 D3 21 2E 63 A7 13 30 3E F8
 96 E8 A5 4A 08 1D EF CC AF 4D 01 BA F3 3E B6 8B
 AF 23 3F 67 15 1E E1 2F 3E 54 EF 21 74 92 CA 8D
 EF 28 F4 73 3C 7D FA 67 D1 44 2B EA 9A 48 9E E5
 CD 66 3F 68 D8 7A E7 E2 15 50 FF 07 40 37 62 49
 43 9C 1B 1A 0D F2 5F E6 03 A9 76 FF EE 7C 93 9A
 F0 31 9A FB 53 8B 5D 4F F8 28 65 BC DC 3D 31 34
 DA 9D 6F D0 53 82 1C 3D EC A5 E6 52 13 4B 95 E6
 AF 49 FB 5E E8 11 15 58 3B 3A D0 74 21 0D E2 70
 2D C0 E2 DF B7 93 7A 41 4B B0 5B C5 55 3E 39 3C
 86 97 69 5B 19 06 A3 43 2B 92 9A 1A 5E 29 B9 0A
 25 BC F4 83 9C 74 18 89 99 F4 9D A1 48 A0 78 8D
 BA 56 83 24 52 EB 1D 69 DC 29 C3 AD AF 23 8C 61
 3C D4 1C 12 64 C6 D9 7C 28 A0 DD D4 E5 6F D3 CB
 E5 90 FC F7 E4 F8 88 6E 24 E2 1D 52 8C B4 7E 66
 52 DF BA 61 34 CF 6D D8 37 4B F3 11 BE F2 E5 1B
 78 FE CF D5 12 C1 3D 98 BD C6 92 67 EB 5F D8 CC
 08 36 2C A6 DD 65 4E 5D 9E 00 6D E8 56 36 25 74
 93 25 09 83 B3 3E 4A 96 9E E5 57 1B 56 BF DC F7
 F2 15 34 6D BB 89 8B F4 1D C8 15 50 6C 10 3B C6
 9B 99 D8 4D D8 32 28 DB 74 0E 1C C2 F0 11 F5 7E
 64 17 6A 8F 0D CA C5 65 8D CD C9 D5 AE 54 06 E7
 36 04 5C 8E 0D 19 36 A5 29 19 23 AF 7A CB 47 D5
 9F 34 CB A2 20 7B 8C 35 60 D0 52 E8 7C CD 29 E3
 D6 A8 B2 1A 4B D7 22 DD 16 73 C4 6D 42 73 15 36
 6C 35 B3 E1 EA 95 94 75 62 95 88 70 FA CC 11 14
 14 C1 75 D8 C5 D4 74 4F 9A 9D 72 BD 6D FB AB 6C
 36 E6 FA 33 65 28 19 7E 30 2D F7 6A E0 E8 30 9D
 A2 C0 B9 8D BF 1F 1C EF 67 76 78 CF C0 6E D8 B3
 F0 5E 3F 72 76 70 94 A1 55 01 BE 5A FE F9 8F DA
 77 8A 73 7D E1 C3 AE 23 4B 56 38 93 6A 3E BE 6E
 99 1A 6C 34 37 0F 0F 38 ED E3 CB B7 E1 1D 43 B7
 5A 78 89 F8 4A B8 A7 CC 2B F0 1C E8 0A F9 61 45
 C7 A3 9D E9 81 89 29 1A 2D 4E 61 A4 52 6D 87 91
 07 3F 3A 05 A2 07 A5 CA FD FD 8B D2 FA 14 A4 8F
 17 5F 2C 1D 0A DB 72 35 9B 1C 91 FD 1E 6E 5D 8F
 45 56 04 C1 15 14 E1 2A 42 45 E5 26 80 E6 7D 52
 33 8F 0D BF 63 FA 97 C1 7C F0 A6 9E 9D 04 B7 F0
 2D DB 7E 9D 12 CF EF D6 80 4B C8 FA 08 AA 69 4B
 7F 93 2E F7 E3 69 D6 9D B2 50 41 D8 BD 65 28 21
 8A 86 72 16 05 71 7E B9 95 56 B3 1F E7 AD 5D 28
 D9 AF DC CC 85 43 F1 A1 41 E6 F6 1E 1C 40 33 6C
 05 80 94 36 C3 AF 0A F4 F3 72 BE 59 6B E4 C4 81
 BB A7 16 6D A4 F4 62 04 61 E7 80 08 CB A5 32 DC
 FB 05 17 48 CD 4A CD B2 6A CA D4 E6 65 D0 F4 43
 2C 4C BA 40 08 9C 5F 8E A3 7E 32 A8 23 C5 05 06
 48 9E 59 40 6D 8E 90 A3 D9 64 59 22 07 21 53 A3
 E7 16 D9 5B 81 A7 20 6C 71 EB AB DD 17 4B 83 B3
 46 76 E5 8C F3 3B B8 01 72 22 E3 29 49 2C FD 8F
 F1 8F D5 75 04 39 AC 99 86 D1 A1 49 4C CF C1 4F
 28 39 0C 0A 30 E6 78 A5 7C C8 97 FE F8 F6 9B 7E
 BC 8C 57 34 C3 6F 4C 66 09 A9 78 09 C7 A6 0B B6
 60 57 13 52 71 16 1C 39 AF BD 07 4E 6D 9B 63 A7
 0A 54 C6 B6 50 D8 D1 02 90 DC 5F A5 58 E6 6A 00
 87 8F A9 0F DA 64 03 C7 6F 92 08 28 4B B5 A3 99
 BA 67 CB 18 D0 9F C5 FD 18 D3 B6 C3 5E 11 4B 95
 5D 21 FE F9 71 B5 2C 76 6C E0 7F 1E 71 71 2E 5E
 2F C9 1E 9E C3 A9 93 CF ED A9 84 C9 06 6E E1 89
 8E 43 9A D7 92 8C 90 61 A6 4F D8 98 B0 C9 DE BA
 00 C1 0C 91 4D 89 22 ED 14 A7 8D 92 D4 FB 6F 0E
 74 27 59 7E F2 D9 F9 75 C7 B4 FC C2 FB 85 D2 0B
 13 0A 57 A4 C5 2F D7 B2 FE BF D2 91 37 1D A7 78
 C8 D6 ED 16 8B A8 32 A4 3B C4 8B 6F CE 4A 49 FF
 DD E4 A1 30 DB 50 47 70 2F 35 DD C0 E0 20 9C ED
 92 32 9C A8 DF 5A 35 AC D3 7B 07 D3 22 07 37 C6
 42 CC 9E AA FC 53 31 E9 6F 7A DF 4F 1E C1 16 52
 97 6E AD B7 5E D4 1D 88 9F 84 D0 EB C2 AD 6A DA
 78 93 71 FC 6D 73 85 86 BE 3F 6D D6 D7 5A 45 B0
 0D 02 B1 F7 20 7A 1A 71 FE 92 B2 AA 56 F3 26 2C
 95 9F 06 90 94 E7 28 54 B1 77 4C 98 6A 1D 2E 29
 24 A3 92 81 01 F5 D1 9F 8A D0 C8 45 89 D0 15 9D
 7B 66 80 15 2A AE B7 CD 01 6B 41 91 BF AC 7E 24
 E4 41 F4 08 28 55 ED FE CA 85 50 8D A6 E4 63 5D
 2C EE 72 06 17 C3 FA BF 77 B0 9E 07 02 AC AB 9B
 E7 E5 8F D9 02 18 D2 66 E4 B4 CB A9 9F 55 1E 58
 F6 F7 01 6C 75 2D C0 08 20 C8 B6 21 BF 46 39 97
 20 F3 C5 6F 06 C4 2F 60 11 43 C3 B7 43 CB A5 74
 54 69 B2 4C 73 C7 0F 7C 6B 3D CF 4E 43 63 D4 E4
 C6 77 ED DA 21 3B EB C7 37 02 E1 32 D8 5A 62 09
 EA 60 91 01 E3 70 63 89 04 4C A4 D3 1E 87 96 D5
 67 82 1C 6A 79 EA FE 45 84 C8 67 4C 34 64 D4 02
 CE AB 9C 59 09 FB D8 23 B1 03 09 E2 2B 92 CD 6A
 F3 0D 47 90 9D CB 09 30 9A C0 A3 22 8E 2E 25 53
 9A 35 F6 28 A8 AA 03 E4 83 46 49 95 AD A8 17 E3
 2B 36 82 70 00 98 8A 0E B9 42 E4 86 4D B8 55 A5
 D8 A4 5D 8B BA B7 D9 F9 F7 8A 4A FF 53 5A 26 97
 0B 09 C8 A5 6D CE 93 33 4D 69 4B 7F 0A 22 56 F3
 3D B3 18 B7 35 C5 DB D2 5E 83 5A 7E 25 B1 5E F2
 17 CB 85 92 80 2A DD 0A C1 E3 72 DF CF EC 41 0A
 5D 03 11 39 1D 75 C2 72 03 9D 9E 34 10 A6 5B FB
 57 A3 15 EE 09 9F 8E A2 B5 B5 F3 1E 77 07 4C 97
 8C E5 FB 61 BA F5 BC C1 3A 2A AF 71 73 92 E5 43
 94 A8 AB 91 80 19 D8 A5 BE 32 95 C3 CD CB F7 51
 B3 42 33 59 CF 81 1C 53 75 83 65 4F 99 1C E9 03
 F4 33 25 43 18 EB B0 B2 21 2B 99 AB 63 E4 31 35
 78 47 56 A5 66 9F E4 26 35 94 C2 EE 78 1F 88 21
 6A 54 A4 06 48 93 A9 DC 10 27 7E 8E 47 06 ED 3C
 0E B0 8C 85 29 31 84 37 23 A5 54 5E 03 7A DA B3
 F2 92 32 79 71 64 C2 6E 4C 4C 34 DD 95 92 8D 61
 B3 CA 26 4E 93 C3 07 43 1B FF DF C2 6B B1 D5 2A
 F0 09 DC 3C A5 44 C0 26 BD BD 78 AF 84 C1 22 E2
 5C 07 47 01 C9 F8 81 4B 5D 47 03 C2 B9 19 D3 6A
 8D 3B 3C 88 04 36 DD 2F 1F B2 EE C1 1C 34 8F 83
 3E 96 8A B2 9E 51 70 59 7D 48 2A 0B 37 60 22 A8
 0F DC 6A 45 58 0B AF B8 02 71 7A 54 89 49 E9 AC
 33 CA AC B4 B7 00 F6 B2 AA 0E 5E BD DE 58 51 2E
 83 B8 D2 9F 49 6A 7D 7B 40 C4 42 6C BE 52 6B 08
 78 1B 02 43 A3 D1 A7 5A B5 B4 29 7B 82 27 E3 B0
 D0 C1 59 9F 6A 55 B9 EC 4D 80 C4 CA 66 8D F0 07
 B3 2B 4B A1 A2 90 18 CF 2A 18 68 3F 0F AC D1 62
 18 0D 4F 35 9C 14 8F 34 13 52 15 7E F1 75 5A 7D
 32 F8 BD E8 F6 C9 0B 00 38 DB B5 9A 4C B2 7F B0
 8A 0B 73 F3 4C 97 16 D7 67 DC 03 E4 CA 4C 62 A0
 42 01 12 37 2A 61 B7 99 1C 81 5B 16 A2 4E 6D F3
 D4 C1 FF 39 80 06 58 5F 8E 31 79 97 1C 6E AF CB
 CE DF 83 7B 81 D5 BE 0C 7E D4 47 B1 D8 EB C7 2B
 BF 09 8C FB 48 20 4B 9B 19 73 FC 39 5A 0B D5 80
 01 DB 4F 6D 1A 66 0D F2 4E 96 A8 D7 7F 8A 10 22
 BF 1D A0 68 18 A0 E3 62 F0 77 56 37 A5 5B 7C 1D
 5A F4 F1 37 F0 BA 6E F6 6F E2 DA DC 5F 81 83 EF
 A1 73 67 39 94 CC 23 04 2B 37 EF 52 7F D4 F2 5D
 04 6E AD 73 FE 09 8F 4B 5E 25 90 2B 4F 4A 88 45
 F3 FD 0F E9 9F 9F E3 95 45 A7 9A C6 C3 0F 1B F7
 23 0C 63 B0 F4 DB 5E 90 BF CE B6 46 F8 4B B8 5D
 58 19 48 0B 3D 29 0D C2 D2 67 4E 7E 6A 45 40 C0
 E9 46 80 EC 53 E3 FF 6F 81 C8 9F 55 D8 93 82 2B
 83 3B 0F 22 7C DF 5C 19 3E 28 BD 91 0B 8E 6B 9D
 B9 59 8B 72 9C 17 6E 4C 33 68 3E 37 4B 8E AC C5
 F7 90 FC 04 52 90 1C 34 46 C5 25 C6 84 6F AD 09
 FF EC C6 9C 7D 26 C7 EF 37 7C EE 44 A3 22 8C FC
 BA ED B5 55 48 70 03 9D 99 70 57 E8 10 C8 6A A0
 B0 D6 B1 3F A1 E6 B4 92 D2 AA F2 CB 3C 9B 9D 82
 B4 DB 19 18 32 D9 58 9F 55 39 09 08 C7 57 36 59
 71 39 50 EB 8B F7 5D 09 86 0D 59 C2 49 03 29 4F
 FB 92 A1 6F 7F 43 CC 0A 06 FB 6D 04 15 E5 BE 87
 9F DA 35 E0 E2 A2 15 9E 2C BC CB 62 C1 68 53 38
 18 81 30 9F 1C 63 A1 30 40 24 99 B4 9E 83 3B A6
 D2 EE 22 2F 13 EA 86 C4 FF 3E 9A DE B4 7E B6 30
 AB 27 A7 33 1C 0F F3 A6 10 74 7F D6 64 AD 37 9A
 B1 C2 80 BB D5 30 5E 1A 9C 65 B9 B8 13 8C EE 83
 BC 8A 84 BE A7 5F 15 9F D3 2E 3E 48 97 06 E0 52
 1E 48 F1 02 F9 F5 D9 B6 29 0F 74 76 9B 1F E3 37
 96 C2 16 79 A6 80 E7 BE 6C D0 40 95 D3 9E 0D 0B
 7A 7E A5 E0 34 4A 2E 5D D9 4B 14 14 79 13 BE FD
 E6 1A B0 11 D2 E5 5B A5 33 2B 13 0E D9 1B 56 A1
 B1 81 53 72 82 CB E5 91 1D 6A 1D 2D 3A ED 2D D8
 85 35 C1 9B 47 60 21 37 8E 3F 0B A1 24 94 46 D7
 17 B0 FD 80 74 9F 27 AB 26 8D FC 4B 02 F6 42 1F
 63 D4 3E 72 C3 6E E0 34 24 1B BA FD 7B 02 5E 7B
 92 4B E7 70 9D A1 B6 02 EF 00 28 D1 59 03 3F C1
 0E ED A7 6A 5C 8F 78 45 7B 83 A5 4A 7E 0C 7D 5E
 A2 2D FB 8C BE B6 AA 8C 51 6E FB A1 6B 79 80 0A
 96 6E 96 54 98 D1 E4 09 62 77 39 0D 3A 0C AA 6B
 1D D7 72 6B 60 DD 72 E9 3B DD 46 39 C8 A0 57 D1
 07 0E 15 61 26 D5 96 75 54 63 FD E6 C2 C0 7F E5
 03 D9 19 50 80 D8 24 F0 98 4F B6 43 8A 58 D6 94
 BC FD 56 A6 3A AE 02 BB C5 2C BE 36 F6 58 42 CE
 23 C9 85 25 ED CD 60 0B 44 05 3F 71 96 A8 19 B7
 82 CB 27 45 74 02 4F 63 60 56 70 F7 55 0C FB 45
 EC 93 61 F6 90 E3 F8 24 D3 22 66 09 15 97 F1 39
 1F DE E2 6B A1 65 C0 10 B3 7B 31 31 B8 A7 FE E7
 CB C2 A1 2F 40 63 D8 AD EF 6E 0B 47 43 10 DD 06
 10 57 29 41 F5 07 11 F4 46 8D 7D 37 CE 98 98 9D
 CE EA 31 AA 6B 6F 7E 44 F4 E0 6B F0 DB 93 A7 FC
 72 26 6A D0 E4 82 81 05 D2 50 1D 56 EC F9 5E 1D
 20 96 DF 42 46 3D 61 3B AE 87 D8 25 45 6B 87 83
 38 3F F4 9F 41 1D F5 DC 00 78 17 FD 0A BF 4F 49
 41 79 FB 69 6F 46 9D 51 D1 A9 80 53 A1 0D 67 59
 9D 2A 2E C6 34 A9 8D BD 67 BB AF 3E 40 52 D1 2A
 92 5C 10 E9 BE 34 6A B1 08 C2 96 A9 09 BB 23 32
 8E 12 EE 27 02 3B DE E8 57 DE 78 E5 EC D5 0D D5
 70 03 C7 E1 19 71 64 0B B8 35 96 2F 82 BA D4 6D
 AD A4 F5 ED C4 81 04 A7 46 FF A7 70 6B 6A D9 72
 4B 82 11 22 C3 B3 1C 14 7C 36 A9 72 96 0D 13 3D
 A5 A9 BF A9 FF D5 CA CD 48 AC CC 98 92 DD FD 68
 B4 8A 1F 5C 06 C7 12 30 60 54 AB 57 BB 69 3B 84
 AC C4 F4 63 68 23 EF 12 BE 1F 86 46 9B C9 E8 24
 F6 F9 66 D3 95 BA 90 E4 56 18 05 8B 23 9C AC AB
 5A 97 BD 36 44 16 C0 FB C9 09 BA E7 A2 6D 56 A7
 31 42 08 9A 69 59 A8 E5 2D D7 1C E9 77 10 F6 EF
 EB A6 64 BF 3D AF B5 FD 4C 20 1F DB EC E0 6A CE
 E7 2C B8 5D FD A6 DF 07 FD 6A B6 93 71 DE 73 2C
 7E 87 77 CD 5E 99 12 1C 18 71 FD 7D 5D DD 4A FC
 68 6A 33 3A 12 74 49 98 AD 80 D1 9F 49 D9 91 F7
 F0 99 30 25 87 C0 9E EB C2 E1 99 65 26 F5 D7 5C
 93 EE 4B 36 F9 2B 59 76 FE 71 C9 CF E2 75 F5 5F
 03 3C 2B 66 02 E2 2D 21 CE DF 6A 49 7C C5 40 1C
 EF 94 A7 3E A0 43 63 70 73 4B 4E A0 47 81 7E 21
 2B 9F 14 FA 82 B8 CD EB 22 1A 2A CA 33 3D C6 FE
 E6 28 41 D8 3F 43 39 FA 2C 32 AB 75 EA EE A8 29
 D5 EB F7 D3 4B 04 2D 69 AA AC 5E D9 AE 71 E2 91
 5B 8C B2 B3 46 AA 8E 37 ED E2 9C C6 8F FF 04 81
 FC 9E FA 62 16 78 23 FB 62 B7 E6 45 AF 28 EB 75
 99 52 B6 C0 A2 C3 29 88 50 22 F3 52 B4 74 62 C2
 08 F9 E1 29 42 E4 CB 66 20 5A 44 17 48 91 5E 43
 71 62 10 76 AF DA 1D 72 EF 3A 91 76 14 A9 B7 0C
 90 87 15 A6 2A 9C CB E0 A6 12 1E C9 69 06 7D FA
 2D A2 F0 28 4D F3 14 0D 3C CE 05 A3 BB F3 10 1E
 04 91 3C FA 5A 4B DC 94 7E 7C 68 46 A5 76 2C 64
 AE BA 17 A6 D3 01 E7 99 82 CC 82 7F 0D 03 D5 89
 6D CC 46 89 E6 7E 6A 80 43 7F CC C9 2A 56 BE 0D
 52 A4 EB 1F 5E 5C 1C 38 D0 DE 64 9E 11 2D 65 2A
 39 75 6B 17 73 6B DD 43 BF 1F A8 ED B3 99 03 02
 43 AE E8 4F 99 49 79 A5 9D A1 F3 0F A9 DD 7B E2
 01 FC 3B B9 9F E0 D2 98 FC F4 92 21 BB 92 C0 F9
 A0 02 3C 33 7B FE BC A6 F2 4F EE EE 2C FF FE D3
 BF 7A 3C A4 8B CA 8C A3 02 46 07 7D 9C 1E 73 E9
 BD 62 43 ED 92 CC 53 A6 5A F9 F5 5F 19 23 6F F5
 9E FA 33 86 5E 8A 49 A9 97 93 EE 9F F9 0E C0 B4
 18 00 FF 72 D2 42 6D 40 6F F2 8A ED 49 38 F0 AC
 A6 99 E6 3A 4C E2 19 74 27 24 53 BB 06 76 CC BF
 24 6C C9 42 9B 83 BA 32 B4 3E 05 62 E4 E4 92 B8
 5F 2B AB 2B F9 29 DE FF F5 AC 0F AA 7B B3 C6 01
 5E 2C 7E 4D 7F CA 2A 1E 23 81 5D EA 6F 32 09 A0
 B5 BF 5B 33 59 5A 7F 52 3F 4B B4 AC C2 0C 1C 67
 C2 46 F6 85 88 38 8B 1A BF 6B D4 8F 40 15 C6 9A
 CA 5C B9 42 62 C9 5E E6 71 04 19 A0 84 68 E2 E0
 F2 C6 3D C2 63 21 4E 21 F7 15 E6 99 AF 8B CC D9
 0F C7 6B 38 F8 6D 16 F8 07 16 72 FE CE 4D F1 DE
 4D AD 01 56 6A E7 7C BD 12 E7 AA BC 76 E8 0A 0C
 27 6B 9D 48 46 2E 74 E8 9D 50 E0 09 61 45 06 B6
 EE FF 35 EA 0C BE 81 03 D4 61 EE 41 76 C4 AB 1E
 41 A4 41 B8 AE C5 33 AB BA 16 8E 5B 49 9E 40 6E
 1E B8 3F 7D 25 75 06 F6 67 0F 03 50 7B 01 E9 F1
 C5 5A 36 CC A9 9A 70 20 C0 CA 34 A3 57 D3 47 17
 3C 41 4E 27 F0 9D BD F9 61 33 B7 50 B5 A1 74 F5
 2C D6 11 92 80 2E 7E 31 EB 05 9B EA 44 DC 5D 98
 42 75 AC A5 DC 2A FC 4C BA 0C E9 EC C9 A4 5C F9
 EE 5B 34 BF 8A E4 3C B1 D4 36 A1 8E 39 3F 99 25
 CA 90 24 E5 82 C4 C2 56 02 23 42 89 ED E8 6B D5
 24 6A 0A 2F 7A FF 5D 07 ED 2E BD 9C AB E1 5A 07
 7A 69 20 A7 42 A8 88 89 08 4D EB 14 50 24 54 AA
 A0 3B 74 8E 64 83 4A D2 F2 58 A9 F1 EE 70 EF 21
 43 5B 4B 70 5A 09 86 9F 39 20 C9 E6 AA F9 F8 1F
 C8 B6 5D 5E 43 9E 65 02 94 3A BB 2E 2D 9D FD B5
 27 F8 71 5A B2 11 B7 00 2D F4 C5 55 13 86 60 66
 A0 89 63 1F F6 5C B6 30 66 1B 22 9F CF 56 8E AC
 DC B7 95 51 3D 99 4E 58 8C 1A A8 42 8B FF 50 1D
 0A E1 6F BC 42 40 35 01 B7 3A 05 F8 A5 D6 69 D9
 FC ED 83 CC F7 BF 14 50 7E A3 5F F7 67 EB F1 E3
 EA 34 D5 BD D9 3B F0 EC 05 CA 18 C2 76 21 53 CB
 A5 D0 4D 7F C5 A0 D2 2B A9 EA 4B 63 10 6C 64 00
 72 62 F5 1F 5D 91 B6 12 E7 DD C4 BF 92 4C E9 B2
 09 66 4A AF E4 88 9B B0 9F D7 5D 48 46 18 F8 27
 CF FE 06 05 74 87 3D C0 EF D4 86 78 B1 DF 10 39
 B1 4B 38 CF A2 D2 3D 72 02 37 76 B5 58 48 CF 90
 10 E4 6E 6E 20 60 44 D7 B1 12 6C EE 22 D2 C7 4E
 73 DB 7D EA 60 7B 6A 81 FD 6A 50 88 4C B7 53 10
 E7 7B DA 48 A0 03 50 D1 6D A4 D1 4E 1B 27 C9 F7
 D9 1C 20 58 DD AC 5C BA 54 30 23 67 4F BB 94 AD
 1B 07 3D BB B7 46 1F 6C B7 C5 97 4F 96 5B 0B AB
 BC 06 C1 3A F7 62 76 7F 69 6C 80 AF 58 38 75 C7
 5E 65 16 21 FD B4 E0 D7 3F 77 8C D1 79 4D 45 3B
 8B 74 8E 8B B3 03 D4 74 34 27 F8 EC CC A4 E2 15
 9C DC C3 85 B8 01 43 EC 7B 56 8C B4 2F 0C 0F 79
 8B 2A BC 33 0C 86 DC 5C ED 30 AB 87 E6 36 FD C8
 5C 41 5E B7 C3 03 7A 69 8F 10 9A 06 C1 E0 C2 29
 AB F1 3C B2 62 91 82 FA 14 C8 8D FD 78 78 D8 E4
 23 01 12 F7 5B 11 04 F8 CC 6B 3E 99 65 A3 7F 27
 7C E2 9A 7F 67 6E 87 75 00 30 4E D4 90 19 7F D3
 A6 66 3C CE 37 FF 8D 86 4E 9C 68 05 3F 88 9C CB
 1F 15 70 B5 E5 6F 26 8F 39 DF D6 A1 C7 B8 65 0F
 FA 24 68 2C 72 8D 47 DF 24 93 06 1D 7B C3 16 55
 5E 22 DB A5 0E DB 0D DE E0 0E B8 1E 7F 7D C4 83
 92 BA 1B 45 40 BC 8B 02 DD EE 96 EA B2 FB 0E 29
 AF 2B 36 7A E5 96 0B 3C EF 11 DE 08 2D 13 60 C9
 65 76 A1 E1 29 72 6A 42 8F C7 85 CF 15 BE 6E 30
 3C 71 DB 7D 7E 4E A4 F3 9A 7F 6D AB 18 B8 C2 69
 85 EE 1D C9 02 47 7B 0A 59 43 7A A0 04 AA 8B C2
 C0 CE 67 AE A6 98 F8 1D 6A 9B 5E EB F8 19 7A 6E
 61 29 FE 9D C9 CA 37 1A 8B 7E 3E F0 2E AD EE 8F
 3D 23 32 B7 B2 25 2C E1 C5 39 CD 61 15 96 9A 74
 CC 79 1A 80 A8 16 E2 E9 4A F5 1D C6 38 2F 8A 45
 8E 54 A0 5D 28 CA A2 1C 70 5D FB 46 73 58 BE 59
 6D E2 89 0F 11 8D 56 B3 F8 17 54 31 B0 70 11 D5
 42 C5 78 8F 8F DD 8E E8 13 FE FB 5F 1C 55 22 8E
 5B 68 58 66 6E 78 BA AE D8 76 90 D7 C1 F5 6C 84
 B0 1C 28 7A 22 19 CE 28 9C FF F7 7C 4A 98 DB C6
 F2 82 FE CD AB ED 7F 77 7B 0F 33 FC 5A 89 82 FD
 EC 37 BC B8 CB D0 37 41 3B 1B A2 E7 1B EF B1 3E
 5D 0F F5 A0 21 3C C2 F4 7C 75 82 C3 D1 2E E3 BA
 4E 94 C5 B9 5B 31 9C 2B 06 A8 8F 2C D0 E2 56 BD
 1C 6D 61 65 B2 D1 84 C3 2F 3A EB 4F AB 99 FB 10
 6E 68 65 6E 50 C3 F4 71 CB C6 1C 83 9D EB 9A 70
 A5 E1 63 FA 91 61 CA 9D FD 8D FB 26 B6 20 15 03
 80 5E F2 93 66 DE 70 B4 F0 E8 9B 77 0E 92 30 D2
 B7 82 8B 43 B9 18 BA 31 7F 47 0B 19 25 C6 9C 54
 26 42 10 FD 57 1E A7 DE A6 6B 6A 55 31 8D B2 7D
 FD 39 A7 B2 04 7B E3 9F D6 4F 50 64 7D 53 BB CC
 9F 94 33 37 7A 73 C7 94 03 3F 23 C1 11 23 11 D7
 6E FE 01 FF F5 D6 23 B4 A4 3A 59 43 F6 BD CC A0
 3A 5B 70 C1 28 FE 90 6A BD 78 D3 70 C5 57 B3 9B
 90 CB 6F 03 7D 5B 82 8E 4F 67 D7 5A 53 86 02 7B
 BA 98 21 F3 F4 66 0F 59 6F 75 F3 BD 68 6D 60 DF
 CD C2 1C A2 99 1D 27 25 EB FF CA C2 D3 14 B4 D5
 C9 8A 81 3F 4D 3B 5E B9 DB F5 67 0F 2A 10 87 E0
 02 06 AE 5E ED CF E3 8C BA 63 E7 C6 8C CC 3B A1
 C2 37 E5 CF AC BE 9B 57 EA 60 10 1F D9 D0 11 A3
 D4 81 8B FF 61 A4 BB 73 A8 B8 A1 E1 5C 28 0C E9
 3A FE 3A 53 81 C2 17 C3 16 49 38 B3 24 14 53 8A
 B1 8B 28 D2 E0 3C 5F 8B 1D 83 EF 09 7A 0B C6 07
 2C D3 CA 78 79 5D 44 0B B2 2E 10 15 E2 CF 0B F2
 BB 2D EE BC C6 4C 45 22 81 E8 F5 31 BB 3F DC 41
 6A 83 97 8A 91 41 FA D6 8B 10 F4 95 5C 32 98 75
 64 37 3D 1D C8 AE 04 84 0B 94 BE 76 D2 A6 50 9E
 7B 23 F2 B2 17 4D 4A 12 9E F6 A0 27 BA 1F C4 B8
 12 AB 17 DB 55 26 68 57 A6 9B 82 1D 6F BB 08 E5
 E5 A6 AF C6 73 88 8A 53 29 23 98 61 F5 B4 8A 0C
 CD 3F 24 62 AD D1 0C 4A 48 69 F9 C3 6D 36 15 6D
 CA 96 D6 2E 6D 15 B8 10 1F 10 1F C8 25 04 3E 23
 A8 F4 72 29 72 57 BD 05 6E F2 B3 3C E7 00 DF 8E
 65 50 0B 53 86 08 E2 57 32 4A A1 68 5E 5E CF 25
 24 7E FA 64 45 FC 6B AB 1D 42 43 5E 48 75 FB 49
 98 6F D6 FD D9 C0 6E 3C CB 44 31 39 96 84 05 78
 30 E1 50 16 2C 8A 69 74 5A 65 E3 52 03 B4 56 D1
 15 97 DA 5A 3F 9E 78 44 F5 BC B1 01 75 68 A2 0C
 E7 5B 1B CE FE 82 54 44 27 8A D2 F1 C9 AF 5E 48
 B1 A8 BE 97 00 2C 28 BD A6 94 3B A4 09 1D E0 9F
 1E 34 3F 74 3B 9B 73 DD D2 51 C9 47 BD E5 B8 7C
 75 C2 74 1B 10 A3 C8 FF 3B 7B BC 3B 95 12 71 A1
 CF B3 9C BD 85 A0 0E 66 4D 00 A8 92 0D A2 C7 E1
 6F 27 5D FB 04 F5 86 18 61 96 8D 05 17 02 CE E6
 CA 9A EF 08 4A 3D AB 9E 0D DA D6 86 E8 77 C7 0B
 84 A2 60 04 B3 AF 3B 55 B6 9D ED A8 A8 B8 9C 28
 D6 8F C0 61 CC 25 ED E3 B4 F9 85 C1 73 36 36 7D
 DF 27 D9 AE 5A 89 60 CB B4 EA 1D FE CC B7 6D E5
 97 65 10 7F 8E 12 C8 4E CF EB 64 2C EA 74 82 76
 A9 32 21 7F 36 26 15 F1 3F E8 E5 6A 8A 6E C4 57
 F0 43 93 72 E0 7D 41 48 90 24 4B 57 F6 C4 36 7C
 E7 9E 7C 49 88 67 8A 81 34 B5 27 E6 2E C5 7A AA
 1B 9F A6 63 9B 2E 80 BA 94 51 87 C6 39 96 8B 66
 C3 64 9D DE 55 68 AF 7F 42 96 70 AE 5D EE 5D DF
 CB 6A AB 30 BF 0F 6B F3 85 C7 2B 1E 24 2E F9 54
 D3 15 71 76 8F 9B B4 53 E0 53 81 72 F0 6D E2 14
 5F C7 EB 1A 14 C3 38 B0 63 D5 55 4D 91 5F 0D F4
 E6 71 A1 87 0F 34 AF FD 80 41 6C 91 F9 40 D8 C8
 9B C5 B2 E8 1C 5A 50 44 17 47 41 B0 81 D5 6B C1
 CE CF FC D0 E4 2B F6 CF 47 8E F5 49 24 72 23 6E
 93 CC 67 47 B2 BA 3F CE FA 62 5F 99 D7 67 11 6D
 F7 A8 BC B7 88 C8 1A CF CB 72 8D 8A CF E7 92 17
 B8 EC 85 24 FD 05 3C 27 DF 58 D5 73 81 56 C7 0B
 D8 2A A7 7F 43 35 BE B1 AE D3 26 10 92 9D 2A E2
 1D D3 D9 11 DE D2 A1 6E D1 AA E7 1C 81 B0 48 8F
 55 C7 86 CE 9A 6D 25 D5 27 DA FF 07 7B 23 3A A0
 83 01 66 F8 56 A1 95 5A 16 64 E1 E8 7E 92 B5 DE
 29 D8 9E 50 93 60 4C E6 4F F5 EA 8D 5A 23 4D 09
 F8 AA 15 45 64 0B 76 5A EB 39 1B 9C 21 B5 1A 19
 52 43 9A 2A A9 20 71 5F 88 65 40 2F 31 CC 4D 98
 54 8C 13 2E 4D 5C 8A DC A7 BA 11 A6 DF F9 0A 94
 A5 8E 1F 1C 5A 57 8F 87 2C 8B A7 37 68 B9 62 50
 5C 2B 9A 04 FB 57 3F BB 5F 3C 8E 76 9D 9A E0 ED
 AD 0A 9A FA E6 C8 0C EA 47 35 37 59 7E B1 7A 55
 8C A2 0D FF B8 A8 93 4E 30 82 85 BF A9 F3 EE DE
 F4 17 A5 5C FB 8F 53 9F E0 69 69 2B 82 32 EE 98
 10 E4 77 13 05 CC C1 2C DE E0 DB B0 91 4A F7 8C
 FB C0 18 02 28 66 66 29 84 50 2E 50 84 D3 54 62
 74 8B 6E 38 E0 60 65 25 66 B5 D3 1A 25 B4 67 07
 0B B9 CB 43 FC B7 35 D4 BC DD F4 0D 30 0D 80 1A
 A2 CD 41 56 99 C1 EA EC D9 B9 2D 9C 4C A9 2A 56
 D6 24 65 B7 25 36 BF 61 13 D9 12 0A EA B8 5F F0
 90 51 62 BB 1C 7D 4E 7E DE 6F D6 F9 77 F9 7F ED
 DD BB 8D 15 90 E4 E2 0B 12 FF AA CA A9 64 4B F0
 30 0C 5C EA 35 E0 CD 5F 2D 0E 3E B2 1C 60 22 17
 30 26 DD D0 3C C5 78 19 CD 46 21 52 10 A4 5E D4
 62 A8 7B B9 E7 67 19 C4 8E B7 67 A1 03 C7 96 7B
 F0 21 91 C3 F4 19 5D D7 A7 EA 13 8B BD 4A 28 AF
 CC 40 91 2C 50 8C 48 D2 E3 3F F5 42 D0 5B 89 12
 79 F8 AF C9 95 FD 79 25 2C 3A 32 1C 27 AF CE 96
 C6 26 DB 57 E9 74 95 62 D0 57 2F 75 E6 DA 2B 3A
 34 00 E2 AE 59 20 CE CD F6 FC 48 E4 A5 C0 09 EE
 35 B1 1C 2B 8A 2B 06 EE 2B B2 A8 D8 8C E6 BC 30
 83 0C 2B 2C C0 6E 52 6E A4 94 DF 2C 7B AF 1C 14
 62 50 46 BE 41 0A A3 4E 6B E7 24 63 76 51 22 32
 8D 30 6F F9 95 CA 35 14 7A 57 9D EA DF A3 54 90
 61 E1 3C 99 45 FA 13 EE A0 F9 A4 DB 70 57 6A E0
 66 D4 88 72 19 8D E0 08 BE 10 F7 58 16 87 58 1E
 EE 4A B5 BF 67 19 B3 05 93 24 BD 4A B4 F0 47 3A
 AE 26 44 4A 8C A3 72 2F CC 92 73 95 C8 D3 B3 D1
 C4 9C 36 9E 3E E7 CA 65 11 73 D2 C3 A8 4F 46 E6
 E2 33 09 DC E0 36 7A 21 CA 47 56 14 A1 FC EB 4E
 23 71 99 63 DD 1C CE 9B 10 85 BE 70 1B AA B9 68
 5F 07 80 2B 5D C2 13 CA 3D 3B ED E1 D1 0D 23 AC
 29 E3 53 3A 9E 32 DB 64 26 C4 B0 82 54 72 6A EE
 47 9B 8C C4 A2 07 D9 F7 34 2D FE DF 0D 3F E3 76
 A5 55 56 A3 6D 88 BB 8A DF 3B 02 AF 6C FF EF 5E
 81 19 15 CC AF A7 43 9F 81 FE 47 A2 24 F7 9D 10
 12 E7 80 B8 FA 25 43 54 F4 00 D3 CC D8 85 5D 6D
 93 65 69 63 34 EF EE 4C 3F A4 56 82 80 10 CB E1
 06 31 7B EE C1 33 7E DA BE 58 47 C7 1C 4A 51 AE
 B6 C6 12 6B 23 82 20 85 B7 89 57 98 44 A6 B9 54
 ED 38 16 78 DB F2 61 3C 28 BF 08 CD 46 DD 11 9E
 37 DF 0F AE 43 7F 7F 0E 90 C3 84 77 F5 F4 5B 48
 CC 07 E0 9B A2 1B 6F DF 66 22 C3 56 A1 AA 69 AD
 A4 4A CC 03 9E 5B 70 30 37 13 4D F2 E3 4A C8 B2
 F9 32 C2 C6 CF A7 11 D4 DB A5 90 BB 51 67 6A A2
 E7 BB 23 03 D0 1D D7 A8 A3 C6 AA 34 9E 1A C2 40
 70 59 8A 4C 40 0B 5E F7 6F E7 B6 24 4E C2 FE 4C
 F5 62 DE DB DA 94 86 BB 5B C2 4C 67 9E 5E 2C D6
 FD CF 3E 3A F4 B9 32 4D 0A BB 08 7B 02 69 2F B5
 7E 06 DA 91 84 58 8A 0F D9 51 3A 5E D7 CF 4A 33
 A8 EB CF 15 61 16 16 18 2F 46 EF 01 24 C7 5C A7
 1F C6 D7 CB 87 D7 34 43 FF 2F F6 BD 95 9D AD A7
 A0 60 F7 85 8F 1C 9F AF A4 15 FD 91 C3 F2 8A BE
 D9 7E AE B4 70 26 20 80 5B 94 EC EF FD 92 65 4E
 6E 3B 56 48 21 96 CF AA 03 74 E6 AC AC 42 63 4C
 22 47 E0 2D 05 B0 F6 18 E5 92 A3 46 69 4F 40 7C
 7F 83 06 2D F5 44 F1 40 2A DB 4D CE 98 CF 25 19
 F8 9C 97 CF 86 C2 50 FD 4F 18 70 75 DF 2A 0F BD
 AA 16 F1 7D A4 71 FF CC A9 7F BB 95 04 76 B9 9A
 82 41 F3 37 3D 3E 8F 67 FF F5 5D 70 10 B3 DE CA
 A3 4A 47 61 86 B7 E1 B1 52 BA 46 D4 FB 2B 3D 53
 BC 2E 44 06 CC 30 E2 8E 9F 91 18 1A 6D AC 53 32
 74 E5 A9 A6 BB 37 69 E3 23 E6 23 D1 06 E4 C1 14
 D3 9D F6 0F 93 74 F8 FF 93 31 3B 6E 9A FF 32 80
 74 D0 89 A1 C8 33 E4 EA AC A3 0D 13 2A 7E 9B 3F
 96 DA 9E 6D 65 C7 19 F6 8E 95 A9 39 B4 43 7A 12
 94 AD 32 F6 24 5D 37 3F F0 EB C8 47 3A A0 A7 AE
 C5 9E 0C 62 91 61 20 C3 FB 65 C8 DB 01 44 60 7A
 C6 5D DC E6 D2 88 23 2D 58 50 80 50 49 9A E0 6C
 56 4D 1C F4 C9 C1 E6 17 35 8D 6E 48 6E A2 30 C2
 30 AA 68 F7 73 B1 B0 A5 AA 25 E8 41 22 F0 AA 32
 5C 6F 2F 9A 87 1B BC B7 EC 1E 6F DD 23 C4 B9 54
 CC 1A A4 F2 25 E3 2C AE 5B 1F B2 DC AF 8D 71 BF
 25 16 F2 16 00 96 48 A6 B0 A7 37 80 33 5C B3 20
 41 72 26 B4 CF 6E AE 4C B2 6C 2B 71 A3 EE 84 C0
 CB F4 45 E0 D6 1B 31 A4 F2 C2 16 00 5A 59 A8 7E
 BA DE 64 A9 0A 21 FE 46 F9 04 0E 12 42 C8 22 64
 C5 2D B6 EF 3D 55 B6 E8 E1 99 59 D6 0D D9 F9 AA
 53 E0 E0 0E E9 6E 6B B9 6A 6C 61 AD CA 00 01 08
 B9 65 BD 08 53 C0 24 E0 6F C0 54 73 34 82 0E AD
 88 FE 0A B0 2B EC AA 4B 40 CA 11 01 6A A9 59 A9
 E2 FC 14 9F 14 55 51 3D 72 A9 11 6A 55 8F F0 77
 1E 97 89 D8 8F 6E 20 DE 7A 29 C3 C3 22 1E 4A 73
 A4 52 EE 1F F7 C9 12 85 AD 3A C1 20 B0 6F CF C8
 EB CF FE B5 6B 8A CE A6 61 08 CE 76 3E 61 87 11
 47 8D 50 90 D8 0F 8F F6 33 BB E2 C6 EC 57 6E 26
 4C 98 A2 AB 64 7B 65 32 C6 53 00 66 D1 79 2B 1E
 D2 B4 0B 42 EA 9A 12 36 1F 36 4E 67 07 CC 94 9A
 73 4F 8E 18 0C 29 16 46 D2 EE D7 12 3D C7 B3 C1
 EF 99 50 42 6F 1C 47 35 73 EA 0E 19 44 AE 3C 32
 74 8D FC 32 A4 0D 3C E3 51 4A 46 17 57 64 E0 1A
 2A 4D 9F C6 20 1E 94 16 1C 5D C6 86 16 F9 11 F9
 19 8C B5 EA 30 EE 44 77 1B CD B1 FB DF C9 EA EE
 9B 2F 2A 56 DC 18 F7 D5 27 0E 9C 61 66 0C 25 03
 96 38 1A 18 E4 31 D5 E1 29 96 F0 4A F7 56 A4 36
 10 3D DE 26 8D 29 73 2F FC B2 4A 0E B1 19 BE 53
 F5 5B 13 42 58 E4 02 D2 A4 DA B9 B9 9B B5 C5 54
 42 47 F1 A4 10 DA 1B E0 15 A4 88 E1 9A D4 BA FD
 B2 1E 15 82 F8 26 A9 35 48 E0 C8 A5 1D 87 63 34
 10 F9 04 79 44 39 57 8E FF D1 2F 45 4F B1 05 11
 F2 9F 93 8D 74 A1 5F 90 07 A8 80 46 C4 EC BB 6F
 C5 07 2F 8E 1D 8E C2 FC CE E7 3A B9 03 07 4D 54
 42 73 9D AC 4F 23 8B 10 66 AF D6 1C 2D 67 15 91
 43 99 63 33 42 CE C3 3B A0 27 04 E5 DC 69 91 EA
 3E 69 BD 90 EA 99 20 A5 89 5C B2 07 D6 F3 ED D9
 10 D5 4E 5B 60 1D C8 12 21 20 0E 56 58 50 23 27
 F5 69 5D BA 11 B8 C0 0B BE 0B 74 1D 03 B9 CC E7
 8F 99 C8 91 FE 5F 4E B1 14 A4 87 E4 7D FD 4F 65
 F8 94 2F 90 9E F9 90 15 F5 04 C1 05 A1 EB 87 89
 75 45 0B 12 11 D2 B5 E3 E8 29 53 8A FC 40 9F 5C
 F1 DA 01 28 A7 57 C0 F9 52 75 D6 01 AB B0 B4 93
 01 01 7E DC 2C 69 E3 B1 64 62 58 C0 AD 7E 0E DF
 41 6C D4 B1 64 53 56 83 65 B6 10 56 79 F1 FB 7A
 0A CF 87 8F 8D D7 49 68 E5 AD 09 EE 7F 89 4D 2D
 C7 BE 92 B0 48 7A 21 67 A6 0B CA 3E 60 27 A7 4F
 CB EE 8F 0C 07 EA A6 BC 35 D4 21 46 B9 4E 08 43
 D3 70 6B F6 B8 1C 88 01 56 9C 05 2A 8A B2 F4 5B
 C5 83 E9 25 E8 BA 7C C9 E5 87 79 0D 4E 0A D4 04
 5C DE 09 36 67 0E E6 31 D9 E2 65 AE BC 52 30 4F
 F7 67 67 95 56 53 49 50 4D 30 F8 A3 6F 48 C5 66
 96 A0 06 AF B3 ED 02 A7 EB 0E 9F 1C 03 48 72 60
 7A 61 B3 26 33 F6 3F 78 8C 0B 9D 8C EA 72 99 6B
 F3 34 0D E8 B2 06 34 11 95 9F 2E 44 9A 44 42 75
 5A 95 9F F2 36 F6 6B 8A AB C3 37 16 81 EA FB D9
 5F 2F 04 61 1D 79 ED F3 7D 68 F9 29 1D 19 50 B9
 45 7E FC FD 4E 5F 44 DF 4C 64 FC 9A A1 DE BE 47
 C1 13 AE AE D9 96 B2 77 BA 05 74 CC 70 7A 07 69
 EF 57 E8 92 29 75 68 E0 6D E7 F2 75 DB 5C F3 2A
 46 11 91 37 35 91 70 62 69 62 56 C3 D1 A3 27 D1
 57 6E A9 EA ED 37 42 8F 51 4F 7A 6B 5F 38 81 D0
 86 1A 01 D2 D2 69 C6 B1 1E E1 8C FA 4C 5B B6 A8
 BB 2C 9E 76 0C AB 19 B8 89 AC 20 0F 4D 74 3F ED
 2F 74 12 58 1F 93 77 C7 70 DA BE C4 3A 48 1D 5F
 6B 43 1E 1F 99 79 C2 A3 40 EB 03 14 C2 08 5F 2D
 67 52 37 88 5C E0 78 27 81 2F 14 76 25 BC 49 76
 69 E0 C0 DA BB 1C 98 4D 46 D5 9F 33 35 F6 EB 9B
 2F 57 51 74 7A 28 6F 6B CD DC AD 04 B0 CA 24 74
 97 21 10 ED E9 30 96 F2 F3 F0 12 68 6D ED FD 3D
 18 49 C7 14 46 39 2C E9 91 9E 81 35 6E 2C A6 85
 B7 43 22 27 BB 83 88 6A 5C 42 AD 7E DD 9A FE FD
 06 25 00 E2 C4 48 A8 DC 3B 3A 59 11 EC 6B C0 79
 89 E7 9C E9 80 AB DE 40 9C 11 83 7D 93 70 E6 9C
 4B 01 60 50 D6 4A 97 25 20 BD 94 B7 F5 7B B5 FE
 6D F7 2F F6 4A 90 CE 03 4E 05 DA 25 C3 2A 4F B2
 B5 C4 E5 A2 07 CC 3B 94 E9 75 F1 00 AD 0D B1 56
 32 B6 48 CF 02 4C E1 2D B7 31 9B B1 56 65 30 D2
 15 EC B0 19 88 22 06 60 65 C1 43 6C 67 6F 38 5F
 AF C3 BF CE 43 A6 5C AB 5A 32 32 A6 D0 08 2A DD
 D5 0E 43 3C 90 CE 4F 14 33 B9 22 DE 22 9E DC 4E
 7D 31 EB 88 34 D5 E4 1F 64 D0 F3 98 FB 9E F5 D1
 9C A9 F5 AF 68 10 96 0B B8 5D C6 1E 5A BF 59 B9
 71 13 88 E6 B5 84 D5 D8 4F 75 A0 AE 47 4B AC 20
 FE 88 5A AC F5 DD B6 37 67 39 69 8A 4C 07 3D 29
 4D 34 F5 41 29 DE 3A C3 33 3B AB 7A E9 88 EE 45
 66 BA C2 FC 83 61 2B 3F EC 1F 4A D4 74 72 54 95
 91 6D F6 53 F6 29 9E DA 2D 12 EF 94 87 01 6C C3
 D1 5B 18 E1 86 62 FF 0F 44 B4 72 55 9A C6 8F BD
 18 09 FD 3D 0D E3 F7 30 28 B8 53 99 20 E4 09 C9
 D4 D1 17 C4 20 6C 84 FD BA BD C3 9F 25 DA 2A 69
 0D 1D A5 49 FB A9 71 08 6C 8A DE 68 9B EB 3C 51
 06 35 CF E4 A1 D6 92 74 1D E7 81 B6 B9 D8 AF ED
 15 EA 83 84 38 B7 12 03 88 36 0E 9D 1C D0 EF 47
 C9 45 6F 5B 24 84 5C 21 F3 9D 21 5B 6F A0 89 B0
 C7 7A 2C CA A1 D0 80 1B 64 4C 84 3D 5E B9 D4 E2
 C5 80 BD D4 0A 71 99 E4 55 6E 33 2F D1 DC 6F 2C
 DA 76 0C 13 1C B8 D4 BC FC 79 C7 42 31 C5 4A C6
 D3 A3 26 CD B2 41 F0 89 14 CD B3 72 CF A6 BB E2
 AB 35 F6 F9 D2 98 87 C2 46 F4 D1 5B D0 EB 74 62
 99 9E 5D 06 0A 45 33 A0 0A 46 0F 4D DC CB DF 5E
 9C F4 36 67 04 69 FF 8D A0 97 B5 1F 42 E7 37 CF
 B1 1C BE C9 75 8A 98 08 9A 87 9A 2E 18 DD 21 B7
 27 30 0D 00 08 A5 59 6B 0D D3 BE 01 32 27 34 A5
 70 90 B1 CE 94 7B 9E 81 40 45 D7 E5 8B 6B 19 94
 19 1E 91 87 2E 87 D4 3D F4 56 C7 3E 25 1F 07 65
 4E 95 0D B5 E6 71 67 81 B8 E3 50 18 69 23 22 6D
 39 CB E8 2C 62 D2 A9 B9 EE B5 41 17 92 B5 D3 FE
 58 9D F1 EE 31 9F 97 62 DD E4 67 2E EC 97 EE 5D
 A3 17 67 BE 48 F0 05 1A 33 90 C8 6C C2 13 FB 71
 27 F1 8E 3F 44 A0 0E A8 84 28 9B 90 52 D8 CC 31
 F0 76 D2 25 FD BB A2 18 D5 52 3D 96 72 1F 18 D5
 BB 3B 5D 0A 34 70 F8 FE BB 03 29 F2 5B 33 3B C2
 C4 76 A5 45 85 16 A4 FB 5B 32 AD 0E 16 60 2A FB
 57 7A EE BC DB 0A 7C 9D D8 8C 65 F3 6E 7D E3 04
 6B 6B 0E 83 2E AB 1B 74 C0 F5 B5 05 65 79 1D 1C
 75 53 77 95 CE 28 FF 0A 94 4E 93 A3 75 FB 37 C1
 16 44 4D C1 C0 C7 33 40 69 77 EA CF 73 A9 A0 C6
 6D D0 85 B0 85 CB 43 43 BC 8F D7 E1 C4 04 34 30
 50 CC 73 71 7C 1F 41 C0 97 2A C8 E8 82 A6 08 21
 87 FD D5 6E 98 7E AB 40 C3 84 63 B0 49 70 2E E7
 6A 05 E5 7B 68 27 B5 BA B0 B5 E9 31 5D 97 6C 21
 09 DC C4 CE DA 83 21 AF 1B 6D 19 4A 69 8F AA A8
 CB 4E D3 A7 75 99 5D 50 74 E5 6A B6 A5 A1 E8 19
 9E AD 6F BD 37 45 E5 69 D7 B3 7B 76 94 05 9A 5C
 86 1E 0B BC 4B 93 DF 56 1D B4 CF AD B9 ED EA 63
 82 E3 F4 D0 A9 71 DD BD C8 30 3A 8B A6 37 B2 4F
 FD 0E 66 99 30 C5 04 DD 2E 9A 26 30 1B 97 D8 7A
 48 80 F4 9F A7 6D B6 F3 6B F4 61 45 00 F8 42 C1
 C6 F6 45 9A C8 10 7A 05 41 CB 1F F1 0C 68 DF 21
 7D 9C D0 71 2C BE 33 50 77 3E FD 02 C9 CD 9B 7B
 F7 24 E2 61 A8 29 85 3A DF 3E A0 76 EC C7 C1 B4
 A9 23 52 8D F0 01 53 46 9B 83 49 99 20 98 08 21
 08 E3 82 B0 66 3F CA 0D E8 44 27 57 F1 F0 63 B7
 B9 AC B7 E6 93 7A E4 E9 EC 4F E1 EC 41 83 8B EB
 49 3A 36 8C BB 0A 21 C1 84 20 33 BF 02 C9 BE 9C
 54 08 27 C4 B5 D2 AF 46 29 ED 04 AB 55 B8 41 CE
 95 31 14 6B FD 76 98 51 A8 A3 D2 D4 53 6D 78 44
 A5 B7 C9 81 DC 00 A6 4F B7 E2 66 D4 2E 32 3E 25
 3B 2C 9B 43 AF CB 07 45 9B 0F F9 68 BE 23 5E 86
 FE AC B2 02 E6 15 78 7A 56 7B 6D C8 5D C2 D0 BD
 96 3B 46 68 34 EB EA F0 F2 FA 99 39 27 4A 09 89
 E8 0B DD F0 36 C5 F3 CD 4A 90 4C FF F9 09 7F 87
 4C C8 8A F5 16 01 65 61 CC A4 E8 C3 70 EF 18 EF
 7E 1A B1 73 FA CC 69 DA 92 14 9D DD EF 28 0A 44
 5F 80 CD 3A 63 22 88 75 C5 90 DE 8C ED EC AB EF
 1A 79 70 4E 29 E4 15 FF AA 91 8D 8C D5 82 BD 5C
 F1 E0 DC 92 83 9A 38 B7 8F 86 97 42 14 0E C4 EA
 48 90 61 44 9E B4 22 46 7A 1F 45 9A 1B 30 D9 57
 42 E0 A2 E9 B8 50 F9 3F 3D 80 50 57 62 EA 79 B6
 D1 31 19 54 C4 D3 57 3A 85 3B 78 1D 2A DA D3 1E
 A0 FB 56 00 D2 F6 56 44 33 F4 4F 51 28 67 D2 32
 4F AD 66 83 88 68 6D 28 17 E7 FD A3 93 D1 75 F4
 5C 34 0A 53 8E 39 B3 38 89 FE B5 D2 89 FF 59 FD
 B1 81 B3 65 83 9A 44 AA A0 3E 69 E4 76 E7 0D 26
 EF 64 EE 08 91 18 E8 D2 EE E1 B6 70 2C 30 82 BB
 FF 98 3F 93 D0 08 C1 8E 87 78 F8 BA DF 60 5A 0A
 BC 63 53 FF E9 9B 06 E9 55 61 3D 1E 17 68 AF DB
 90 D7 89 1D B8 16 1F C3 A2 85 59 B3 1C 29 68 28
 A0 47 99 D1 B3 27 C3 7D B1 2B F6 48 25 8F D0 D4
 2D 41 CB 27 39 79 88 2E 6C E3 C7 30 48 F2 0D E2
 7C 16 EC 91 49 F4 0D 3A F3 2B 49 5E F4 D4 06 DB
 08 EE 26 4C 1E 8A D9 23 F6 A4 E9 84 D8 C9 96 E2
 88 4B F2 8C 79 0B 6D C4 70 71 97 8F 2B 15 B3 86
 F4 31 EF 8D 10 10 15 03 F0 A2 02 A0 3F 8A D2 44
 EC 92 A6 08 E1 51 99 C3 70 B6 3D 62 9F C5 63 A2
 0A 89 8E 6F DC 1D D7 6E B2 2A DE 7F 2F 4A CB D4
 83 60 83 B0 AC A2 AF 64 85 B7 89 FF 44 A3 E8 5E
 A8 91 87 65 1C 39 A4 54 AD 2E 35 EB DE F7 5C 12
 9C 27 B6 5B A6 A5 C8 C3 00 5D E8 DA 19 CD 1C C6
 F1 D9 3B 32 65 E1 09 1A 19 47 BE 25 06 4A C2 62
 BA 44 F4 74 C9 4C 22 18 20 1A F0 9A FB C8 7E 03
 09 FF 74 AB 1C 0B 90 74 FD 54 99 DE 67 64 39 CD
 66 D4 ED E4 89 BC D1 45 87 1D 82 BE 64 9C EB BB
 D0 DC 47 B9 2A AC E7 B2 A1 39 EB E3 6F C1 1A 0D
 56 3F AB 89 A5 DD 56 87 71 30 07 1E 1C FA 94 BD
 72 1A 0F 49 C7 EE 90 10 6B 94 EA 48 4A E1 84 41
 AB F0 20 74 F4 FA EE 9E 5B 6B BE D1 8C 58 CC 61
 F1 E5 F3 7A 25 0C B6 23 F5 E2 39 FC CB 9C 77 15
 B8 92 C9 3C 08 B4 9C 70 16 98 94 96 62 7A 13 0E
 6F BB 68 61 A7 24 A7 5C 86 57 59 E4 BE 89 21 ED
 3E 96 5F E1 93 07 18 30 97 BF A9 28 B3 9E B2 C3
 2E 3C C8 81 A6 0B CE FB 66 80 E3 C1 6D 18 06 C6
 5F CD D5 17 4B 09 F8 E9 96 64 35 31 C6 4B 77 27
 88 66 BB 98 63 D5 F9 97 93 0C 48 CF 98 0F 82 3D
 07 BB 8C 19 4E AC 80 23 E3 93 8A BC 8F 41 0F CB
 74 D0 9B 3E 27 C0 09 F9 EB F2 FA B3 28 09 AC 2A
 1C FF 86 9B CC 8A 32 FA C6 05 21 9B D1 5C A9 CF
 FC 9C 4F 68 75 31 6C CF B2 01 61 5A 18 6B D2 9C
 78 A6 F0 F8 8B BD 5D CB AE AB F7 B8 3C E5 56 6B
 6A A5 0A 24 7E D7 28 34 0C 15 15 BB 55 7E 31 CB
 FF 03 C2 EC 25 F9 12 27 28 59 24 40 C8 9D AD 2B
 58 A6 26 1E 0E 3A 71 E6 28 54 AB 43 C9 FB 86 3A
 42 50 5D D6 D6 26 60 A3 36 93 7E D1 4E DA 4F 16
 61 DC 11 4D 48 67 56 1A 26 0C E3 07 B9 86 0B DA
 CE F8 1A 47 69 34 E5 CD 16 F4 C4 19 2D 23 1C B5
 25 72 AA 42 15 99 24 71 0E 3F 07 70 37 E7 46 A3
 42 CF B4 5C D6 CC 7C 49 4F 53 7F CD 83 B6 66 29
 FE 51 A9 3E 9A 3C 10 8D 81 B9 90 D7 4A A6 73 EB
 26 5A 95 23 04 2A 86 6D A4 6E 58 CD C1 8D E5 32
 C1 C6 C0 05 36 53 98 16 56 22 D7 82 FA B2 D9 56
 E6 EE 6E 88 8A 27 6B BC 92 86 B0 AF 84 72 7C 52
 A5 72 04 76 C5 36 F8 12 62 AD 35 EB 7A C0 42 10
 BD D2 40 6F BF 0B D5 4B 1D D0 B6 FA 04 36 69 C3
 AF B8 AD 30 70 BD DF 31 A2 01 5A EE E2 0F 0C C3
 26 AB FB E2 9E 5A 28 99 36 BE 2C F0 FA E1 5A 3E
 68 5A 9A F5 5D AF C6 56 D5 A9 8D 57 97 68 00 6C
 9D 8D F1 C7 5B E7 D9 A2 71 9B F0 97 D4 8A B0 48
 D8 8B 70 DA 7F F0 34 3A CB CC 6D 4F 76 EE C7 8C
 18 19 38 35 F6 47 CC 97 D5 03 A5 04 B3 DB CE 55
 A2 BB 63 F2 6D 10 BC 8F 24 6A 8A E3 04 BB A9 38
 83 EC DA 1B E3 A1 FF E2 ED B1 69 5A BD 48 5B 01
 5E 23 38 F5 A7 EE E3 06 0F 22 BC 25 F4 E8 E8 85
 7F 93 B0 36 50 0D 8F 62 9A 9D 4F B2 DC 3C FD CC
 9C B3 C5 2C 7D E0 2B B1 5A E0 98 13 CD 08 45 14
 8B B5 71 F9 E4 75 A7 40 B5 A4 DA 9F 46 0E 00 0C
 CF C9 BA A2 ED 31 44 5F 21 C0 5D 26 D4 9B FF B0
 D5 97 2D 2D F4 44 0E 3D 42 4F EC 71 54 E9 B1 24
 73 79 ED 01 0E 0F AC 49 BC D2 AA 18 88 5F B8 CF
 25 72 60 51 1A A4 2A 3D FF 0B 9D 70 AC 46 D2 2B
 FB 89 27 A7 66 74 76 C6 02 96 CF E6 B3 23 6C 65
 F9 FF 7C 3C 52 DB BD 46 54 74 16 59 5C 7E 94 10
 A5 CC 4D 2A CE 3B 94 DB 34 6F 97 36 76 29 D8 43
 EB 02 6B 71 16 71 F0 C5 4A C0 EE 34 82 AD 2A 36
 20 0B 5A CE 33 85 D0 E6 F3 FA 14 F9 7F D8 1A 7C
 14 4E F2 A7 FF 4B A6 A1 DE B4 EF 80 78 53 BD E5
 0D 49 9A A1 28 50 73 90 6C A2 9A 3C DC 60 92 5C
 92 D3 E6 B8 50 D7 3E 49 82 AD 3C BE 4D 67 4C 2E
 BE F0 A3 2A E5 77 EB D7 ED 17 88 F0 EB B6 D0 BC
 AD 5B 67 FD 5D E7 33 83 71 47 15 0D 09 0D 92 F2
 A8 7F 0C 70 8E 01 95 DD E6 92 82 35 8B B9 2E 3B
 4A 32 BF F1 56 04 51 53 A5 54 9C 44 51 AD C9 90
 DB 0D A6 9C EA 32 ED BC FD CE B6 20 C9 E9 F8 F2
 F8 49 16 4F 6E 4C 98 19 0A 93 C9 BC 37 C9 D6 A5
 83 0A BC 57 7B C2 69 84 FB DA 88 69 75 1D 7C 2F
 F1 79 6F AB FF 20 0A C4 D4 EE 8B 7E AE ED 0B 02
 6D 9E 15 4F 96 02 EF B4 BF 47 70 E2 CE 85 E1 F1
 E2 F0 A6 30 20 2B FA 18 30 A9 A8 A7 75 2F 04 65
 5B F0 BD 7C C7 13 C1 EF 38 28 25 AB 33 09 F4 A7
 AD 85 B3 E3 DD 05 73 B9 D3 10 C6 EA EF AD F2 F6
 CD 8B 5A 50 DB C5 E9 96 BF C3 72 EA 40 7D 56 27
 67 39 2C 68 0E 16 80 1B 50 3F 67 A7 A7 78 D0 4A
 1F A9 77 5A 7D 77 6A D4 E4 35 D5 7A BA 7F A2 21
 DB 77 D7 D1 A0 A0 7E 71 37 2F 7D 4B E7 77 A6 1D
 BD 10 55 90 45 28 8E 8C 8D 40 52 22 36 21 56 F2
 22 F3 A0 F8 57 AC 47 A7 AD A4 8B 54 32 7A 8C 51
 81 C0 22 47 DA FF 14 87 51 9C DA 92 A9 E8 7E 15
 51 1E 40 04 A5 71 3C 20 BC 78 C1 F8 59 2E 6A D0
 B5 91 9C 59 84 76 08 49 61 C9 6A C6 93 99 E6 6A
 24 94 38 8F AA 22 C8 CA 7C A4 EF 94 7B 36 99 D4
 0C 9F D3 68 EA 7B 33 8D 3A 94 76 22 8A 54 5D BC
 1D F8 45 BD 77 EC C8 30 14 BE 23 96 FE C6 63 2F
 CF FF D7 41 1C C4 FB 91 CC BB 0B 8E 6A 1B A1 4E
 1D EF AC 58 56 9A 07 B7 F5 51 B7 75 20 F9 85 82
 15 AD 1B 3B FD 8D CF 6C E8 67 FC 21 F4 2A 32 DC
 E6 51 09 EF DA 06 F0 D6 1C 65 F8 26 3B E7 CC 6A
 44 C6 A9 8E 24 24 45 E1 AC 0F F9 C4 32 2B D2 DD
 11 04 BF 81 FA 04 EB 6A 75 CE E0 E9 F4 8E 01 AF
 18 6E E5 13 D7 57 DE F3 6B 4E F3 3A C8 6B 3D 61
 CF 5C 0A FF CC D5 28 73 E8 F3 59 DB 7B 3C 21 6D
 F0 AF B6 7B C8 24 F2 CC 31 25 2B 44 A3 FF 8E AD
 53 40 AE A9 A9 52 DD 17 15 B1 73 A8 58 40 47 50
 75 3E CC B9 C1 59 91 14 DB BF 07 3E 96 E0 18 32
 A5 49 E4 23 B7 55 10 90 C8 32 76 70 7E 72 CA 14
 42 D9 B8 A3 C4 62 10 E5 5C 53 CC 03 6F AA 95 C4
 DF E9 39 14 C0 51 61 B3 17 5B 56 E0 BA 8C 5B A1
 F9 D4 F3 A9 15 77 69 92 75 F4 19 A6 AB 1F AA F6
 13 E8 B3 BA 08 05 3E 70 66 B0 D4 F7 B3 E4 58 3C
 D7 53 83 78 B2 9E F3 98 D6 14 37 77 44 4C 8A BB
 70 C8 B0 79 AE B1 44 7A 2B D4 8A 58 45 35 78 90
 B3 30 A4 6D 9B 83 4B 0A EC 4F F0 D5 5F 20 18 E5
 EE 8C 92 EF 64 CC 60 5F 2B 94 4F 3B 69 15 33 83
 B1 16 F2 66 40 C5 C3 99 C9 87 64 54 84 23 90 9F
 CF 86 0D 6D 9D 0B FF B1 5F 7D D4 D3 31 31 22 8C
 80 C5 E1 52 6D A3 F1 58 EC E3 DA 67 8F 20 12 19
 17 01 8B 96 07 7F 0F 32 56 5E BC 5E 93 6F F7 87
 E0 A5 88 AC D1 96 13 67 CE B1 01 3A 7F 28 3D E1
 0A 27 CC B4 30 0B 9A 50 CF B1 A9 9C DC 20 38 D6
 DB 61 7A 5A ED D8 7B EB 04 2D CE 79 FF 0A FB 63
 95 A8 3A 4F FB B1 33 8B B0 0F 4E 9D 7F FD 5B C6
 DC A5 FD 5F D5 C5 23 5D 14 F8 C2 AB E6 AB 9C 7C
 1A B9 DC DB CA D9 50 68 E8 08 0B 17 B1 30 31 4A
 D4 EC F5 74 08 DB 68 8B 96 BC D2 78 36 54 7A 4F
 C7 AB 2B C6 71 3E EF D4 0C 4C 87 55 DA E3 8A 64
 88 2C 7B 02 76 29 24 1E 28 C9 AD DB 67 F5 D5 56
 A8 81 FD 6D DF 19 E4 9E BF FC D6 DA 7A 79 6C 44
 34 FE 8A 83 75 54 73 C8 4D 85 AE 15 85 A5 B6 81
 56 9B 1F 53 C4 79 E5 DC 26 13 FE 45 D3 E1 94 4C
 5C 70 6A E9 37 ED 35 25 B7 31 C1 5F 53 95 5D 58
 10 E1 76 9A 25 1F BE 55 FC FB 7B B2 07 58 36 F1
 CE 3F 8D F0 34 55 04 62 6C 41 06 49 CF 7D AF EE
 2C 81 F3 63 B3 5D E8 4C 77 0C 2F 9B 0E D2 23 84
 09 BC 0D F3 17 81 AD 68 77 DE B6 4F 36 4C A8 97
 A3 4A 73 29 90 B2 BC 9A CD 26 F8 D4 7E 62 57 7B
 9D 30 A9 3F 9B BC 34 44 DD C1 09 B6 8A 52 1F F4
 DC 8A 9E 6D AD 5F DA 19 BE 5D 5D A7 5C FE 40 A9
 B1 76 9C 61 AB 50 41 63 BA C0 54 BF 6B A7 76 AE
 86 D9 E7 15 3A 3E 0F CA 05 42 AB 7E 25 36 54 03
 F9 80 7F F2 67 78 7A E9 A7 F5 EF 79 D2 4E 0B 85
 D6 A1 D2 94 37 99 E7 F6 48 5E 39 12 00 89 31 21
 15 8F C5 C3 E0 7D 49 3C 78 3F C5 71 76 2D D3 A8
 2C B3 21 24 7C 49 EB 38 03 79 CA FE 15 E7 6C 2B
 2C 4E 7A 31 20 04 57 51 D2 4B 15 54 9E 5C B6 EB
 06 79 80 34 87 39 0A 6C 97 01 D5 85 79 8A 0C 47
 26 D7 6E 24 B6 35 C3 D1 F5 F8 64 B2 91 1A 09 6C
 95 58 67 5C 45 3C F4 50 3E 2F 45 06 1F FB 80 86
 B9 05 A0 41 1C AC 31 36 04 0B E2 99 52 F3 97 84
 08 04 22 F6 17 6B B0 3E 70 0E 0F D8 1C 37 EB C3
 20 A9 75 78 0F 81 AD DB D5 D4 47 38 BF 01 97 B9
 67 F9 6C 80 F2 10 2A 0B 7A 2D 10 05 A9 23 F1 B4
 53 71 85 FF CF 10 F3 21 92 58 D4 BB 3B 8A E5 64
 22 49 3F B0 52 66 29 B8 7F D6 5D 82 1A FB 63 8F
 7B E7 E4 82 0A 7B 3C BC 55 88 E3 39 04 19 7E D2
 0C 05 92 1E 9A B4 30 A3 77 BB CE 91 D1 C1 42 C0
 EE 10 30 48 C0 30 19 10 CD B1 C7 AB 29 BF BF 91
 51 A7 F3 F7 AF FD 06 BD 0E A5 97 80 68 89 1A AF
 F3 64 76 04 49 1A 92 8B AA 20 9F 49 CA D3 35 FB
 CC D9 A1 02 84 A5 E9 F0 D5 C5 D9 D3 32 9E 9C 87
 2C 28 6B 29 48 F1 F8 93 58 86 4F 82 EF 28 B1 DF
 7E 39 52 79 DC 63 B2 AF 83 75 7F E3 42 4C 7B EB
 C9 3D AC 05 86 E8 4A 54 DE A4 0D 6A 95 93 56 3A
 A9 06 52 05 65 DA BC 89 BF C9 40 0B E2 47 12 34
 B5 36 65 7C 63 73 1D D0 94 C7 1F D9 5C AF 37 44
 A9 B4 0D FB 58 F3 3C 0D 0C 87 71 DE F3 1F A1 A8
 E0 71 07 6F B9 10 C7 F0 28 95 21 67 EB 21 56 23
 66 C5 16 5C F5 3E 5D 65 98 32 17 5A 98 E9 36 6E
 70 24 50 76 91 B1 90 B5 82 D1 A9 DF 36 54 1B 3E
 08 07 02 5E E3 13 E0 D2 D1 F1 5E AE 3A 98 A2 9E
 22 6B 76 20 EA 0E B3 3B 95 B1 7E 59 C7 E4 1E 89
 95 C5 D9 B9 FF 61 79 E2 D0 F8 43 23 BE CC C0 83
 0E 6C 6C 86 C7 91 F4 91 9F A5 1E 67 4A 81 35 3F
 88 E5 B8 DB 3F 07 4A A6 F5 B1 B9 E0 7D FA CF 37
 E9 31 35 39 38 E5 8E 33 A2 16 8C 10 2F 56 B0 B1
 AB 47 FD 8C 8C A5 52 78 F2 23 1E 1D 4F B1 D2 08
 B0 3D 70 23 AC AD 02 63 CE D5 C0 B7 BB 78 E2 C8
 A4 C3 ED E2 03 46 EB 54 CD 6C 7C A8 C2 31 69 3A
 A9 85 45 42 13 87 D7 95 43 83 2A 28 A1 25 64 9E
 88 DE 8D BB B1 F7 71 D2 AB A4 72 0D 7E E2 2D BB
 E1 03 76 A1 DB 02 A2 89 6E 41 D6 3C A3 F1 C0 EB
 6C 28 74 C4 43 83 ED 28 C2 DA 12 3D EB 22 93 A4
 28 F9 8B D3 E1 E6 CD 8F F4 A0 F6 01 E2 01 2A 21
 DA C7 B0 F0 8C 62 65 7A 40 D5 5F BD 03 B6 9F 59
 C9 12 E3 93 54 30 D9 F9 FC C1 1D 4A FE 36 68 23
 47 4D 34 2E FF 88 67 EE FF 28 66 B8 39 9C F9 0B
 A0 CF 19 BD 8C 2E E1 70 2D F2 92 D3 ED 8F EA 3B
 14 FF 5A 8E 37 FD 95 9B 96 9C 6D 0C CB 01 1C F4
 D5 16 68 13 08 06 F7 3C 50 86 3A 43 1A 5B E8 92
 D0 C5 C8 EF 90 97 E7 D1 19 A5 72 B7 6E FC 12 E8
 28 02 7B F5 D0 83 6A F6 62 B3 17 DC 08 D9 4C 7B
 30 2B 20 39 6E 3C F9 41 8D F7 DC 40 05 FF FC E5
 18 06 66 66 90 78 3B 1E DB 9A 0A A0 DA AE E0 E9
 F1 F3 00 C2 98 FA CA 93 47 BE 38 B8 0C 0D 3D CE
 88 45 92 DC C1 8E 13 FF AB 78 FD 0D 20 FB 06 1C
 F4 57 BF 6A A6 E1 BB DE A2 73 05 AB A8 22 B2 AB
 9D BC C5 27 79 62 D0 D4 66 6F 64 B7 42 AA 60 CD
 81 97 20 46 A8 FA FD BE D8 B9 61 1F 5B A9 31 93
 95 75 12 70 57 A4 9E 1F B1 A6 D3 8A 7C FD 24 E0
 1F 9F A1 6E 9E BB 47 70 29 10 14 7E 12 CE F2 BF
 A5 1F 42 2B 98 39 01 F1 CD FD A0 7D 3C 06 D7 AA
 A1 F9 EC 0F 28 71 87 ED 88 BE 59 C8 28 23 D7 B6
 4C 56 82 F8 6D 96 4B 65 17 F5 E5 FF E0 6C C3 C7
 8A D0 AA 43 B2 7F A3 6E EB 0B 67 DC AB E2 95 06
 6A 79 0D E9 2F F4 AD 96 5C D4 EC 6A 88 EA 9A 9C
 64 32 D1 53 CE D5 69 DD FF 68 76 E0 EA 15 09 39
 F1 0F 2A 38 2D 1A FF 33 64 24 31 BD EB FA 49 68
 7D E1 F8 2F EB 0C ED E9 52 C6 AB 47 6F 5F EB D1
 D8 C0 14 A8 85 83 3C 4C 86 EA 29 CC 6A E7 1A 6F
 1C 8A 7E B1 59 AA 21 08 2C 04 F3 9D 15 14 33 59
 A0 9B D5 F6 FC EA 00 BF D5 97 D5 33 AF 2D FC 7D
 90 36 EA 3D 25 8B AB CF FF B4 E6 FF 9B B9 ED 14
 6F C2 E9 EC 32 E5 EC 5D AC 63 49 97 1D F1 8A 74
 26 C1 D0 AB FB D8 30 84 41 3E 67 E6 EB 0E A3 CE
 50 D4 7C F2 FF 8A 9C 14 14 19 24 0F BB 42 83 60
 57 B9 C7 F7 05 6D A6 10 14 05 C5 48 4A 44 F6 55
 6D C6 35 E7 65 C2 0E 02 C9 2E D5 4F 38 0B 7A 5D
 45 98 27 8C 96 59 9C 33 4E 58 6F 8B 9C E6 60 71
 40 40 88 59 9E 43 AD E1 D6 FB 3E 5A 87 4C CB B1
 9E 9F C8 04 1D 97 8A 70 CB 6F B5 8D 27 A7 59 E0
 5E 90 A4 EB 4B 9A E0 34 3E B4 75 4B 6A 87 E4 9B
 86 ED 44 6E CA D0 36 D5 63 BB C2 8F 93 44 CD D5
 59 72 DF DA 5C 26 48 FB 9A 12 61 DD 91 94 9F 37
 31 32 BB A6 DC 54 9B CE 76 9C E8 0C 7D 9A 92 BE
 F0 D9 FC BB D2 6D F5 73 06 14 81 D5 36 F6 A8 E9
 49 65 FD 9E EB ED 5E 49 B4 2B 91 8E E1 9A 52 9E
 7C 7F AF A9 A0 69 E3 2F 13 3A 90 3E B2 33 20 42
 D3 1B A7 9E 19 7F DB 92 E7 B6 DA FC E3 57 15 2D
 EE 55 AF 52 A3 CF ED DC 1D 22 60 9F 8C 6B A0 73
 E2 BD C2 BE 73 3A ED 8B 32 C3 BE 00 16 D6 C0 57
 71 A1 CB D7 C1 06 BE B2 5F 1A 48 0A A2 8A A1 C7
 0A 82 0D 9A 19 04 AF A8 28 54 45 ED 2C E6 45 4A
 65 F1 6E 58 C8 18 23 5C C8 82 57 15 65 C6 40 A2
 32 89 E0 34 15 B6 6B A8 66 19 BF 2E 34 C3 5D 7B
 D1 F8 EC 65 DC 39 0D 36 5A A6 C4 16 6C 32 35 43
 E7 F9 1E 03 18 95 07 B0 84 FB 65 AB 8B 06 9C CA
 E0 A3 18 16 5F E8 7E 59 C1 49 46 2D D4 7B CC 94
 47 9D F1 99 11 94 F2 C1 AF 0B 43 C6 4A FF F2 E5
 0C 0E 91 F7 D8 B6 65 2A F6 8B BF D7 EC 87 E7 A1
 62 09 A3 0E 92 17 16 1F 01 21 72 78 F7 98 20 88
 7A 1B 5D 36 45 F9 D6 96 A9 F4 E5 55 8B 4D 3C 16
 F8 50 91 31 B8 29 77 1A 96 D6 C5 16 A3 97 09 BE
 DC 18 E0 3A 84 52 97 8A A6 B1 CB D2 D6 43 E9 34
 EA D4 72 90 8B 98 32 59 3F C5 A5 19 AF 3F A4 D3
 C2 6D 0B B6 C4 30 F1 A6 F2 F9 1A 63 49 A0 C2 37
 25 7F 9F 74 5B 2B AA D2 F9 76 5B D8 C2 02 2F 8E
 B4 86 91 3C 21 ED 47 1C 75 70 A7 45 2D F3 50 5D
 6D AA B1 70 46 67 10 5C E2 2F 2C F8 3F 0C A2 95
 1C 62 E4 D8 F1 DF 62 26 5F FB 95 9D 76 EF 76 06
 29 DB 1F 6D 29 44 07 DA 5D 94 4C F2 C6 61 6A 03
 71 2A 24 A5 C6 4F 53 E6 16 C5 6E 4C 37 1E B6 8B
 22 94 FF F5 0B C8 0A D4 7F D6 9B DF 61 B5 75 7A
 24 4F 16 A6 ED D9 11 27 53 D2 6E 5B 52 98 09 C9
 52 AF 25 3D 86 63 E8 F6 7A 47 33 16 00 76 67 C8
 FE C7 81 13 A7 B9 CE BB B9 A6 65 52 67 2F 6F 15
 00 3A 59 DA 91 70 D3 97 C2 FE A3 9B 9C C9 A6 D8
 AD 19 DA 2E 65 BE 66 C4 08 FD BA 09 84 3B 62 B5
 09 64 2C E1 2B B6 1D 5F 8C 76 18 14 06 13 6B 9B
 6B 1A 8B 34 A3 8F 57 58 DC 20 8F 27 4C B6 56 7E
 B4 CF 5A DC B4 4A A3 76 8E 18 70 80 8E D5 F4 13
 B3 32 53 55 05 6C 27 57 E2 42 F2 FC 3A C9 E3 9D
 50 25 1A 56 50 2E 9C 88 8E 7D 01 5B CB 02 78 E4
 3B B7 8B 12 83 02 EF 39 DC D9 50 FD CD C8 20 9E
 7C 52 93 4F A2 9F 3D A8 94 AF 88 7D 8D CF 8A 06
 BB FB 8A 20 C5 9F F8 63 EE 8E 4C 17 0F DE F1 81
 A4 94 32 4E 74 3E 36 D7 54 AA A2 82 8B F7 75 39
 47 89 93 CE 77 53 E8 30 43 CD 99 50 A8 4F 67 94
 1D 5E 34 77 FB 88 08 99 93 20 55 9B 77 86 7B F9
 BC BE EA 9B FE 0D E7 31 27 36 4F 98 12 5B 74 7A
 8F E1 A0 FF B8 D3 A1 1A CB 0B 2C 79 50 41 71 B0
 4E 62 C6 7B D9 8D 01 E8 FE 7B 76 11 92 14 BE 6E
 2E 8A 7D BD 27 0C 6E 0D C6 C7 CC 60 4F 7F 4D C0
 EB 16 B2 56 21 88 AF 2C E6 E0 82 F1 CC C4 96 7D
 34 38 FC 01 3C 14 91 96 39 EA 30 65 77 7D CB 60
 F8 D5 36 B7 7F 96 75 DD 34 36 93 7F C7 FA 88 21
 3B C3 E5 BA 22 4A C2 F3 74 69 D9 5B 99 E3 EF 3D
 04 4D 47 A1 2C 5C 48 2C 6B 56 FE 4F A3 E0 58 C2
 4C 32 36 3F E5 38 F7 5A 8E 07 BB 64 0B D7 A2 60
 75 70 5C 79 29 44 45 F9 F1 24 1D 7F 52 A5 AA D2
 35 71 E6 21 50 8C FB 74 17 44 3E 64 DE 88 1F D8
 40 BF 8C 77 23 29 1C D0 CC 96 AA 38 8B C3 A0 32
 5B 8D F2 E7 20 D4 74 B3 E0 74 D1 69 3F F0 9A E4
 25 9E 7E 3B 98 6A DE 5E 65 F9 88 87 B0 48 D5 B2
 91 87 D8 BE 50 DD 23 CF D3 17 B2 D7 99 7F 10 7E
 B4 BF E6 9F 6E 67 A8 B8 FF 9A 3B 04 3E 9E C3 62
 E5 9C 97 0D DA AE E0 8E DC FB DF 1B 57 1D D3 2F
 4A 4F D9 37 25 6D B0 D8 55 0E B4 D1 83 FB 7F DA
 48 CE EC EE 3B 8A 12 DF 9F DC 97 66 08 FC FB 5F
 02 6E 9C DA D6 15 31 FE 6E 96 AB C7 74 2F 98 92
 56 11 9E D0 B5 15 32 D5 43 D1 41 4C 3F 11 04 AE
 63 DB 55 67 3A A9 09 31 C7 E7 BA 56 E4 34 D1 E9
 8E A4 F1 24 03 41 25 E6 7E AF 9F FF C2 5E 1E 9F
 5E 33 8D F8 F6 89 95 87 D9 DA 69 44 4C CA A8 24
 8A 3D 28 D9 45 49 D2 32 BE 70 F8 B6 6E 98 E6 10
 D8 0B 4B F2 78 16 8B E0 D0 B8 AF 09 B8 28 A2 C8
 E2 71 F3 C2 09 03 D6 F7 D7 8A 9F E4 90 83 C1 02
 8C E0 B7 EF A1 84 B6 C5 AA 69 79 73 40 4B 2D 7B
 04 37 D3 97 E6 E2 18 2A ED 09 CB A7 E0 DD 10 1C
 4B F5 16 DA F6 EF 7D 3C 75 3B E2 C7 36 50 82 F5
 F2 0E 30 05 79 FC E6 F6 F1 93 9B 34 42 42 BE E4
 38 22 FD B0 15 FD 03 00 1D D4 D6 AE 7F 15 B5 E6
 36 C7 53 BF 7B 86 2F D6 28 58 C0 85 26 D1 8D 4A
 F4 A9 51 FC 94 44 F3 80 68 1C E6 59 C3 1A 76 5D
 6E 2C 6C B1 C8 09 A9 70 12 80 17 5B 7B 94 C8 CE
 D7 A5 40 40 0E 9C 4A A3 70 55 95 9D 59 33 95 E3
 63 CA F3 33 32 8D DB 2F 5B AC 08 2B 13 26 1B 7A
 32 DD FC 1E 45 0E E6 72 BE 35 92 0C B8 A2 42 8F
 C3 8A A8 EE 7D B9 11 94 F2 C2 A0 3C 77 DB F8 A5
 50 F8 FF 63 6A 21 F2 67 5E E6 6B 28 C2 C1 6F 74
 66 8D 15 8B 39 E0 D3 1B 6F D0 83 D1 3F 2B C9 3F
 E1 77 5D 58 5B 8D BA E3 33 F5 87 02 3F FB 39 D1
 E9 99 A9 3A B1 4D B0 F0 B8 B8 D6 04 66 D8 09 1E
 19 77 C2 AE 68 72 57 0A BA DF 3A DA 16 5A 79 7F
 9B A7 19 7F 3C DF 8A 12 A8 85 A9 8F 76 9A 09 64
 7F C0 6E 4D 52 8A C2 0F B8 4B BE A3 DC E1 52 C2
 98 1E 22 5F 7C 03 41 17 FD 90 38 A8 29 D4 CF 60
 E8 E6 F5 11 82 8A 69 FE 85 A9 88 B0 EE A6 3F 45
 78 6F A3 A1 EA 9C 8E 54 F8 D5 37 0C 06 5B 49 72
 AC AF 2D 07 18 0B 02 57 C4 47 E4 13 96 46 ED D6
 86 87 F0 E5 E6 22 88 15 23 44 3B F3 3C 66 42 DB
 69 47 F4 9E 53 7D 08 78 2A 0D 29 03 97 3B C4 25
 DC C5 C0 E3 C0 75 FF 57 52 38 2F E2 8E 24 3F B1
 43 56 D0 2D 28 B4 92 C8 7A BA 57 8C 5E 50 B2 9A
 AA 91 78 51 8A 4F B6 C8 3A F9 1F F8 2D 34 FA D4
 B4 69 BC 98 F8 22 7D 5C 01 6B D7 0D 37 A3 23 77
 33 6F FD FC CC 5A BA 84 9F 67 35 3D D6 93 8F 19
 99 D9 97 B0 06 A2 54 62 3A 78 5B 74 F1 0F E2 CD
 FD F3 05 7F EA 7D 12 05 38 47 FF E9 88 2F FA 45
 34 E8 9B BC 0C 36 ED E7 0A 63 B2 99 61 68 B4 97
 15 BC 27 6D 22 F0 78 53 9E AB 8B 79 8B CC 11 70
 8C 89 F2 04 D6 BB 7A C8 46 0E 1A 9A 32 BD 34 C6
 6B A4 09 16 42 52 45 BA 6C 09 E8 1E 86 4A DE 20
 63 E2 19 40 65 79 C5 22 C8 28 97 40 43 E7 8D DE
 E4 EC 69 E1 53 5F 35 90 8D 89 49 19 26 61 BB DE
 F3 52 D5 8A C6 14 3E 6D F8 2A 3D DB A3 E1 CE E9
 1F 10 AA 29 88 66 B5 B2 96 D5 34 50 B7 6A F0 0A
 58 80 93 FA 30 D2 14 04 36 CC 67 7A CF 34 37 06
 99 09 73 62 23 07 D2 47 53 56 D5 34 CB 56 86 30
 77 A6 EF FC B9 D8 D4 8B 9E 24 D9 D3 E9 EC 05 1A
 DB B4 36 1D 6E 93 4E C9 F6 C3 4C 6F A7 A2 E7 B7
 E6 52 88 AF 75 E0 87 82 AD EA D7 55 15 F9 32 C3
 DA 13 62 BB A8 C0 E3 14 97 6F 31 11 9F FF 2B 86
 65 9E 90 33 0E 42 20 84 45 08 7C 1A 4D C9 FC 9D
 1D 4C E2 D5 96 9B 6C C9 82 2A 34 11 80 C9 FF A4
 33 DD DC 23 29 F6 C3 C0 FF D8 4C 82 17 A2 AC E1
 93 84 D8 BF 8E AC 67 00 36 DA B6 44 88 97 61 4F
 55 F0 EC E2 F5 05 ED 57 68 CC 2D F0 BF BD 16 10
 0B 55 69 96 DD FC 25 90 24 BE 0E 28 71 58 8A F6
 74 7F 78 93 41 EA 2F 2E B0 6D 16 89 51 7D 88 87
 92 3E C4 AF B4 2F 2E 41 F0 AD 06 F7 A3 34 33 2E
 45 68 BC 15 83 2E 88 E2 12 73 CD C5 0C 89 C0 15
 5E F5 CE 0A D6 7F 65 BB F1 8D EA 29 94 69 3F D7
 42 62 6B 2F 89 47 E8 BF 31 A1 57 9B D3 F9 EE 57
 F0 8B 54 72 EC 34 B8 06 6A A5 7C 48 DE CC 46 93
 CC 9E 2C 43 1D 28 EE C0 B5 17 4C A3 FD 0F DF 29
 9B 67 CA 6F 0E FD 48 0F AF 86 6B 34 40 17 B5 5A
 17 3E D1 05 F4 49 09 3C 17 96 8A 3F 38 8C C7 38
 4C 1F 6E 40 B1 7D E2 07 5B 2E 32 92 25 13 9C 36
 CB 89 8D 52 7B 2E 1C FD 5E 8B E7 64 AC 72 07 6F
 B5 53 AB 37 8C 90 DA 64 39 B8 0E C7 29 F6 AC 43
 24 FA D0 2E 6A 0A 35 49 FB EC 13 0B 34 7A 9E A3
 89 46 60 FE A2 F8 C0 9B 86 14 77 D7 31 26 EA D8
 1E 4D E1 49 6F F7 B2 91 EA D6 09 92 01 CE 0A 98
 77 50 F0 CA 0B 45 26 C8 7F 45 3A C5 73 44 A0 01
 27 58 A8 3D DD 92 94 A9 3A 63 69 DC BB 84 C6 B5
 EE D5 E0 D8 6C 58 53 3B D2 CA 43 D7 15 D1 42 C3
 6A 45 07 FE 94 BB AE 79 58 90 02 D7 72 A2 5F E4
 2C 27 BC 82 DC 68 07 37 89 8A 9B 41 A0 EA EE D3
 F2 7E 99 39 AA E6 B8 4C CB C5 D8 97 8B AE 03 70
 8B AE BF C6 EF 0B 76 C6 2F FC 95 2A FE 46 22 0B
 C8 FE 61 81 C9 A1 5E D4 6D 7F 91 FB 3C 1F 4F 55
 EA 17 39 B0 E0 69 EF 77 F3 A0 6F 19 3A 19 8B 60
 04 90 76 23 F5 9D F3 77 94 16 30 21 18 89 92 36
 E2 27 25 C1 C4 02 D0 12 C0 7F 03 5C F4 4E AE F1
 F4 4A 5A 1D 43 05 51 C2 75 24 4F FB 0F 82 D4 88
 37 10 C2 D6 EC 99 71 35 4A AF B2 BA 64 64 C6 DB
 D6 80 3C C0 A4 8A D5 50 11 A9 0D 5B 40 35 0C 90
 38 47 B2 AD 82 42 41 40 34 D6 04 00 D6 6B E3 B2
 F0 23 BD 20 C2 63 37 52 5E 44 F4 BB C6 D6 A5 32
 89 3F D5 F8 19 B2 2C 11 4C 77 80 04 2A 2A B7 4A
 29 FA EB 3A B5 32 DD B2 B0 2F 6D E2 76 E5 43 E9
 95 CC 1F DE D9 3F D0 73 08 18 03 06 27 9A 7C 46
 98 21 DE 8A 82 F2 03 D9 63 FA 6D 49 B5 BE 23 73
 DC C9 7C C2 A9 F0 DA AA 21 79 51 58 6E 86 F6 B0
 87 E3 3C 69 D9 93 D0 DC 00 E7 69 2B 3B A9 DA 45
 C1 C5 71 36 FD F3 42 94 C6 98 0C B8 20 24 C9 4B
 7E 80 87 BD 3E AC FD 9A E8 17 E7 19 B1 36 55 95
 9C 28 FB 11 23 87 EB 4A D2 AE F4 7F 57 E6 EE 02
 F8 99 E7 3D D1 A6 E2 0D 85 28 67 22 18 88 62 87
 8A 38 09 1F 62 E4 42 FE 9F 23 57 E9 35 57 40 3F
 A6 5C D6 69 A4 8F 46 DB AE 4E FA 1F 48 5A 4E 75
 45 B1 DB 5D BE 48 51 C6 2B DE 2F 79 43 A8 F4 25
 74 6F DB D8 AC 88 F6 39 B1 DA 6A A6 88 DA 66 F1
 33 B1 60 A9 62 66 4F 53 51 4B CF A4 F3 3E 40 DE
 6A AB FE 92 1D 8E A6 82 32 82 E8 6B E0 CF AF 73
 99 60 9C B1 4D D8 3E F9 C3 97 B4 D1 97 D9 68 FF
 70 72 68 BC D7 A8 C3 9D 24 98 B4 06 E7 01 7C B8
 3B 0B 83 48 2E A9 F8 D4 A0 64 7A 54 AE 0B E5 FF
 14 B4 53 33 AD 18 D2 93 E4 74 2A 55 FC 6E 55 1A
 76 A9 43 3D A4 76 65 FE 57 46 29 33 E3 13 A4 D3
 E1 DC CD 25 9B D5 11 C5 A1 82 F4 69 18 47 CA 08
 3B DE E9 38 95 4E C5 4B B0 D8 68 9A 3C EE E2 0D
 C3 E0 9C E5 52 44 7C F3 82 83 66 EE D8 CD F0 35
 3D 5A EB F6 14 59 89 67 E2 0F 19 34 9C A2 D1 D8
 29 6E 53 64 96 95 31 D5 AB 9E 2D F0 52 08 F9 8E
 2D 50 C5 2F 36 BB 02 16 BC B1 65 21 45 C4 4C 35
 71 B0 4D 4D 58 42 E0 28 B4 A5 7F B3 1A 70 70 C6
 C7 DC 92 7B 94 F9 3B 68 02 49 A0 27 B6 E2 DE 17
 C6 BC 5E 46 C0 A8 88 6C 02 22 DF BE 3A 8D 38 F7
 3C D2 94 5B 68 F9 44 56 38 EC 8A 8C CB 2D 74 A8
 A4 52 1C 20 3E A1 19 50 63 CF D8 42 C7 8C EB F7
 68 77 3A DC FC DC 3A 94 CD 63 C7 D1 C1 44 40 62
 83 22 93 5D 0D 49 A9 5B 4A B2 A9 2C 79 AA 10 7C
 FF BC 53 DB 36 08 38 9B 38 3D DC DA 0B 23 24 C0
 02 A0 17 9D 8D 43 8F 86 4D AA D4 D1 FE D7 90 D4
 DF 0D C4 96 24 88 4A 90 37 15 3F 98 F6 40 3B AA
 D6 B1 CB 2C F5 ED FA 54 7B 0E 18 A6 BC 4F 61 DD
 E8 32 18 86 60 D9 53 41 9B 96 66 57 43 F2 FD F8
 BA 48 C1 DB 17 4E CD A6 48 85 BB E5 C4 B8 E0 31
 53 FB 95 CA BD 35 DB E7 EE 21 15 58 8F 18 C6 27
 35 ED B1 55 C4 57 10 71 86 20 FF 1A AA F7 0D 89
 56 B3 2A D5 43 5A BC 0B 25 E1 03 57 B2 09 E8 F0
 30 ED 1D 75 80 85 DE E5 DB FB 98 3D EE D8 05 A5
 A2 2D 75 81 D5 9B 90 5E 8C 13 5B 47 CA 54 4D E5
 54 9C 31 40 15 4D 65 C0 AB 3B D4 C2 8E DD F1 9C
 18 2E CF 93 C8 5E 61 09 E4 83 EA D1 A4 44 34 7E
 16 B7 75 EB B8 5C 48 04 3B 7E 06 82 01 C3 9D E8
 E2 68 0B 58 80 FA BC F8 BB B6 B7 90 06 34 B8 AE
 EB 7E 00 34 99 0F 4C AD B1 3E FE 55 A8 DC 4A 3F
 95 08 A9 13 86 EA FB C1 30 01 E6 48 8E BC 29 48
 51 1B 73 7C 64 4F C8 13 3D CE 7A A8 45 A8 04 99
 BA C7 92 E4 95 38 07 39 52 C8 DC 38 AD 54 12 53
 41 63 65 6C 82 B3 9C 87 B6 0B 5E 15 EC BF 97 FF
 92 59 7D B1 8E 01 A2 6D 8C 3E E9 1C 9B 5B FF 51
 23 23 2A 55 13 48 5E FF 83 29 FC 4A 45 52 53 BA
 AD 13 DE 98 14 84 CC 21 8E 8E 8E 53 EF 4C 4C 97
 E8 84 3C E0 71 1C 22 DB E3 C1 54 36 AB 5A DE FE
 B4 81 FA F1 2A FC CB 31 82 F1 B1 F7 30 83 3D 3D
 10 B8 7F E0 83 0A 02 65 0B 1E 99 F2 A3 87 DF CD
 45 67 E8 F3 D4 3D F1 94 80 F0 D7 B7 7C DC 1C E3
 86 6A F7 14 13 29 B6 EC 74 8D 64 A8 9F 0E 01 1B
 A3 EF 9D 43 CA EF 9A C0 F7 5E E1 5C 79 51 87 33
 37 B9 F7 89 5B F0 6A 53 F2 FF 50 19 3D 80 66 2C
 56 65 01 8D FD 5B 0E F1 B3 5D 3A E0 38 F7 F0 F3
 99 D9 B1 0C F8 E8 5C F1 A6 AE D2 0F B9 61 93 6F
 51 CF F8 FC B2 61 FA 22 AE 59 F2 64 58 D6 21 08
 46 24 EE 64 61 1F 50 77 69 ED BB D7 EC 09 5A A4
 20 28 13 EF 5D C6 46 10 35 24 F4 30 90 BA 73 74
 75 AF CB 49 8C 21 B8 60 14 27 3D 58 72 3B 42 14
 91 C1 B5 10 CC 88 AE B1 37 14 CE 5A 29 DC F2 76
 A9 DA D7 9B AD CC 2A 42 EC B4 A1 62 16 74 3F 70
 0A 9C 50 D0 F8 51 F1 2E DF E1 97 76 9A AE D0 D7
 54 C5 01 E5 A1 99 30 03 79 BC C2 A4 82 51 E9 01
 7B B8 D4 93 F2 9E 7F 0E F2 8A 32 A5 C0 5F C5 EB
 A3 7C D1 29 98 B8 D7 29 7F 38 E5 9F A4 2B DB 1C
 DB 1B 97 0E C6 68 E7 02 9B 6F DE 7F 56 53 70 FF
 FB FF DA C6 24 BD 9D CC 81 F5 E9 B8 CD 98 85 B4
 FA 8E 14 25 F7 E3 55 BB CB 44 C2 EC C0 96 3A C8
 70 D3 E0 5A 45 1C 23 5F 0C A9 4B 0A F1 00 F0 D4
 47 4B C4 37 1E 8A C4 3B D7 3A F6 2D 0E 71 30 A2
 9D 58 72 6F D4 1A 72 02 E3 38 3B 81 7E 73 DF D8
 E1 A6 07 B2 3A F2 61 9F F3 CA 1D 88 04 26 8C C3
 D4 09 1A 1C 40 2E 87 39 5C A2 B7 C9 9B E7 3E 2C
 4F 3D 07 53 14 D5 22 6F 9B 3A 54 57 71 97 09 89
 C6 59 E2 DA 60 DD BA EB FA E3 60 3A C8 50 A3 03
 FA 1C 1C 14 B0 85 48 E0 E2 FC 88 00 27 1E 78 0A
 D5 1F 2E 14 F6 6C 12 6E D0 AB 40 28 ED 35 7E 9F
 86 56 F6 CF 6B E5 19 56 3A AD 52 50 63 0D 11 D6
 82 9B 31 66 09 07 EA 31 A5 B4 34 DC 6C 09 6E 97
 F6 6A 30 9D EC B4 14 65 8D 23 CB 5A 89 31 E9 97
 46 B4 1C 49 F5 92 1C 57 A9 2D 53 CA 05 0A AF D1
 F0 B8 C2 2A 44 34 5B 23 D5 F4 F1 10 E4 F7 F5 EA
 32 CB AF 52 11 11 2D 4E FD F1 25 86 7E 63 0B 6A
 86 3A E8 D2 59 21 BE 31 1E 44 69 FA B6 62 55 44
 14 44 33 49 11 FA 23 0A 79 DF 10 7B B1 36 D1 4C
 59 D2 B3 9B E0 3A 06 F5 97 E6 93 89 1B BF D6 F1
 D4 3E 1B ED B2 39 E1 C1 64 6B E8 6A 35 F5 61 29
 99 36 E6 6D 22 58 8B 5B 50 87 9A 93 26 01 6E F9
 AC 15 EB 53 1C 3F 6A EA C8 56 19 AB CD D6 DF 8E
 27 29 BB A4 77 68 18 2A 82 05 51 22 C8 60 B6 E8
 03 83 D0 7D 28 47 B1 89 9E A9 90 75 DA FE 8A C8
 00 0A 7E 31 82 84 77 7F 98 F3 D0 81 46 73 87 66
 F2 D5 A4 2D 6B 97 D9 5F 53 51 25 C8 F2 B8 A2 78
 B4 35 EB 6F D8 B6 31 CD 0C E0 AC E1 FA 34 AD 09
 47 7F 2B 6C A3 7E 6C 28 E1 BD BD AA 16 D1 23 1D
 C2 1E FA 88 15 9D D0 63 BD 80 B8 37 AE 27 0D 9E
 78 E2 E0 C7 FF C5 E1 38 BA 55 37 66 6D C3 90 B2
 C5 D8 A0 60 A7 8A 8F D4 59 21 82 37 15 50 21 AF
 50 54 11 8F C6 CF 9C 5D FE BF 92 0F DF E2 1E 99
 36 90 A6 F4 15 4D 63 DD E3 8E 87 35 17 53 CA 1B
 BE ED 19 D4 F7 D0 AF E7 F5 9D 91 08 D7 C9 7E 44
 68 59 8D 41 22 56 88 4E 1A 71 95 2B BD 7D CC 45
 F2 63 E8 BD DC EC 84 76 EB 4E C0 E2 F1 3F C5 D9
 E9 44 A4 71 FF 69 ED 0C 34 B9 FE 5B F5 94 6C 55
 FA 4F 7A CD B0 AD 37 35 AD C0 54 9E C3 3B A7 C8
 98 9C 58 2F FB 8E B1 80 9B 93 7F 4E 11 0A FE 95
 4B C5 1B 85 CE 0C 60 77 88 51 A3 F8 64 89 B7 3A
 EE 95 5F 60 7E E6 25 9D DB 09 0A 59 05 0A 7C 59
 83 53 B1 7E CA 19 9D 53 AE D4 09 49 39 0A 23 53
 DB BC 3A B6 82 03 0E A1 8F AC F2 1F C1 2D B8 49
 88 5E 20 84 26 C4 35 00 F7 2C 59 27 4A CA A6 2C
 4F 7E 88 14 83 48 27 58 DE B2 AE F4 70 B9 68 B1
 7E 2C 54 58 23 A5 02 06 17 76 CC A2 3B 5E 8B C6
 5B DD E1 9C 88 6D 02 0C 9A DC 81 FE 19 9E C3 15
 83 42 6E 14 BD 92 F4 61 A6 39 EC F5 00 6C E5 1C
 B7 10 9B 43 71 A4 45 22 AD D2 B3 2F 48 BF 90 99
 89 B5 7D 76 75 A5 CB 6D E3 C2 C8 BB 73 9B 25 AB
 D1 9C C1 AF 06 4E 78 E1 12 6E FE 29 AF 82 6A 99
 6B 4F 86 63 F4 4D A7 7D 81 86 6D 67 81 36 79 3E
 76 60 42 2B 0B ED 09 9D BA AD 78 E2 D8 74 A4 5B
 61 0F 55 11 39 C5 08 33 8B 0F 70 8C C4 DC 9D 34
 9B 40 13 C7 2E 21 49 52 C2 FD 02 46 4F 4A B4 5B
 F6 09 A6 03 AF 8D 56 C7 59 FE 66 35 E9 F1 DA B4
 C5 88 C1 59 71 98 1D 56 FA 86 E2 A5 E7 28 28 23
 88 D0 3A D8 B9 CA 71 A7 D1 BD 18 89 91 0E D5 0B
 6F 4F 3C 94 96 B4 2A BF DB 6E DA 43 AC 7C 54 33
 BC 57 3F A8 48 88 A0 8E 82 B0 39 D9 D8 C3 A4 AF
 50 FD FA 79 FF AE DE B2 CD 38 E2 E8 97 93 D8 14
 C3 8F 0C D0 C9 73 79 28 AC E3 CB C5 6F 0A B9 95
 54 46 DF 86 95 AA 2A 78 B0 06 AF 7A 9E 1C 0F E3
 56 94 96 BF CA 99 A3 2D FB 2C 51 7D 75 73 1F 43
 6E 53 73 8E 03 D5 C7 D4 39 D7 2E 31 A3 1A 40 79
 07 11 4E 0C 0A BC 2C 2C 37 7C 69 5E 21 56 92 24
 7C 56 04 97 63 E9 F6 6C AB 56 6C AD F8 FA 1C EC
 B0 CF 32 15 36 A5 99 6D EA D5 8F 86 62 6E C6 16
 38 65 5B 09 10 EF DC 82 5D B3 32 9B 23 F9 5C 1B
 F2 C7 89 68 D6 66 8A AF 2D 4E CE A1 3E D6 73 48
 0B 33 8E 2D 78 72 4A 8A B1 B9 C3 03 81 D1 34 65
 CE E2 7E 91 6D 51 2D 79 9C 8F BF 2A 82 AE CB 0F
 19 04 51 BD C9 03 17 8A 40 77 9B C4 57 8A DA 70
 E4 9C E3 8C C6 CE EC FC 5B 8C 4C E9 AC A9 A6 DE
 0B 02 5B 3C 27 08 2D 11 20 2D B3 3B FE 5A D6 BE
 EB E2 BE BA 9A EE EA 18 57 B1 26 E2 CE 02 AE C4
 5F 41 45 36 52 6C 10 F8 B7 7A 7D 61 D2 F6 78 CF
 6E 4B CB 3B F5 83 D6 10 8D 47 08 1F 47 11 01 7A
 39 4C 67 90 08 B9 08 6F D4 A6 A7 BF 7B D3 26 23
 FB FB 96 B5 44 E2 47 25 8D 94 9D 19 EE C3 8D 5A
 51 88 C9 96 38 74 ED 09 58 30 AE 03 7F 9F 20 21
 CB 0E 01 51 09 C7 23 7E 38 0A 2B 23 F2 6D 17 E3
 88 F3 55 16 68 E2 6D EE 28 13 A1 15 8A D1 9A 04
 A7 DD 3E 0A 96 1E 36 7D 6F 70 8F 41 B5 41 1C 19
 D0 24 3D 3D 23 00 62 F4 FE AA 4F 04 8C C0 CA 3C
 8C AA 4B 02 3B C8 D0 47 5E D7 12 84 0A ED 5A 97
 6E 81 29 26 D8 59 2D DC 4C D4 0E 75 F8 52 08 11
 C6 4F 88 AA 8B B5 36 67 E4 C4 8D 26 16 57 57 E3
 E3 1E FF 77 4C B7 1E 99 82 3D AA A8 50 BF 69 22
 BE C9 2E 1D 12 34 B3 A4 67 B1 B2 5B 7A 01 81 6A
 56 6D AC 91 F3 44 FE F6 93 5A 46 B7 1A 3A BA 2C
 B2 8D D1 6C A9 C3 1E 10 F7 86 26 FF EC AC 2C 57
 02 CB FD 54 A8 63 D1 C2 34 FE 9D 4B 57 7C 74 24
 2E B7 4E 16 05 CF D6 80 19 10 8C 05 43 7A F0 2F
 13 B9 9D B9 41 16 45 F5 FF E3 3A AC 90 0D D0 17
 03 C0 09 15 5B 57 BD D2 DA 22 D3 1A D5 CD CF 0B
 3D A6 30 0C 75 C9 8B D9 E5 58 AB 64 05 07 3D 4F
 EF 61 68 15 F4 54 1E 52 07 B9 DE 6F 61 4A 58 A4
 C4 92 4A 78 BB 9D CC 48 80 31 10 8C FB 1F C2 61
 53 2D 67 B5 79 F5 4E DC 75 D0 C3 BF 80 01 E1 D0
 6F 27 68 6D D6 66 1D EC A2 A0 29 20 52 DE 2F 02
 DF 7C 7B 0D 38 02 F2 18 18 19 C8 36 CD 9A EA 07
 B9 38 08 28 E4 FC E4 FE D0 71 88 87 90 F6 AC E5
 0A E1 FB 68 3D A1 03 84 74 2F CB ED 93 27 3E D5
 C7 F1 78 FD 41 AC 6A 58 70 F3 76 E5 C3 74 EA C0
 0F DA BF 1D 29 01 0F EE 02 35 8F B2 62 30 88 77
 94 60 FE 93 E6 C0 8D 5C 9C D7 59 94 34 9D 90 E3
 AE 3F 0D 15 C7 12 B6 F5 06 67 47 9E DB 74 FB 85
 FE 72 F5 13 4A 4C F6 AB EB DB 9D 33 36 1C F9 41
 7A 4D E6 08 2A 08 67 62 F2 C0 71 71 44 A4 33 89
 9F 26 F6 B3 97 6D BE 6E 43 01 59 77 B8 1F 7A 9A
 86 9F 86 65 B7 A7 FE DE 28 5C 09 97 F2 2C E2 20
 37 AF C4 C1 6C 98 5C 19 AE AC 87 31 FD 7F E1 D6
 B8 83 98 17 30 3A A0 AA C1 4C DA 7D F6 29 22 E3
 64 18 0B 15 57 88 94 C1 F2 31 9F 73 68 49 37 38
 67 B3 2A DD B1 37 23 79 4D 24 64 19 95 B9 FD 88
 DB 5A 5E DB 44 6E 1D F2 6D 80 5A 16 58 12 00 45
 F3 8A 78 A8 0C 7B AC 96 32 39 7B D1 2A 6B FA 1B
 8D 9F 81 B4 0D 89 44 3F 7F 58 B6 25 D4 84 CF B1
 BD 65 F3 D8 47 E5 81 79 95 EA 0A C0 0E 9F BF 41
 CC 3B 74 28 F1 D2 57 45 B3 A1 A7 F0 68 EB 65 B3
 52 92 F7 E0 94 FD 2E 0F 65 36 95 A5 CA 0B B3 01
 74 19 ED 81 55 A8 BC 90 80 43 6B 7F F2 60 4A B6
 01 E5 99 43 58 60 E5 6D 66 49 F1 B1 F2 56 F7 18
 F3 4B 3F 01 D7 36 33 B9 9F 97 B3 B6 2C 8A 22 1C
 5F 4C E6 F8 A2 A7 AA E2 97 B1 7E 91 31 EC D7 FD
 FD 23 7F 2B 31 E7 D9 56 F0 7D BC 59 2D F7 55 C7
 25 C1 C6 F7 F6 64 09 1D 68 B7 21 2A 06 87 E0 25
 C7 ED 47 FF 6E F0 DF B1 F6 63 98 14 18 72 D3 C5
 34 8F 4E D0 F5 22 13 75 9E B7 09 E5 82 21 22 D9
 91 4E F1 CB B4 B0 DA 69 9E 6D 54 F4 21 A8 63 A7
 A0 ED D3 76 3E 00 01 B1 5B B4 1D B2 29 3D EB 84
 32 84 92 21 50 E0 EA 2E 68 84 BD 73 2D 48 52 18
 F1 1B 7F 75 2D 76 C6 E8 96 93 58 B3 AA 00 65 00
 2C 09 C3 A6 54 74 7D 19 15 55 A5 5D 43 3B B3 6C
 DA B5 BE 69 7C 75 29 D7 FF 51 F9 7B A0 6A 57 D6
 1E 69 D5 FC EC 93 2C BD AE 73 2F 19 95 5E 96 92
 2A 0C 18 83 89 B8 08 56 F7 E6 66 B8 21 57 45 22
 2E 04 22 B0 9C A4 89 4B B0 B1 4D 11 87 E7 22 16
 9E DA 2A 3C 36 FD E1 6D 5F 3B 6F EA F1 5B FD 35
 47 90 CF 9D 81 F8 E2 B2 67 67 98 DA BD 4B 5C 30
 F1 B8 DB 80 F0 35 A5 26 40 AC EB 20 20 F9 5E 12
 06 A4 23 22 A9 97 44 A4 84 C2 3A FB 86 14 56 B4
 ED 3F 74 0B D0 E1 E3 64 00 85 65 9A 0C 8A 18 92
 67 F3 3A A9 3A 4E 73 30 0D 73 AB 4C 66 97 0C B5
 E0 F1 83 23 68 D3 20 62 5C 22 75 AB B9 7F 55 12
 35 78 9D A1 50 A4 6C 0C BC 38 96 55 F0 76 72 88
 9F 50 8A 05 CA CD C2 8D DC 99 C4 FA 2C AB AA 00
 FB C9 62 52 27 B2 7B A8 D9 EB 34 17 F3 80 78 45
 17 E6 33 3A 2C 15 B2 8C 73 2B C6 64 C7 3E 46 FF
 CB 8A F1 D5 01 72 B7 0E 05 27 36 F0 B8 86 FF 29
 85 73 90 51 9C AD E3 9A B8 89 63 FD B9 99 65 C1
 09 52 23 EC C7 F9 19 85 F4 69 F8 5C 6C 32 A8 25
 7E 08 EF 9F A7 D3 C3 9B 6F B7 8B C0 62 49 4A 31
 A9 B1 51 26 83 AB 58 22 23 4B 42 37 39 75 FA DC
 1E 4F 79 39 5A 49 88 E3 D2 12 3E B6 EB B6 30 FE
 22 C6 69 9A 22 40 8F 70 11 13 ED 6F 4C B1 D5 AD
 63 A4 50 E8 5B AA F4 80 B2 FB B9 F4 D0 2C 45 47
 42 1E EC F0 0C 6F 2D C1 2F 70 C5 41 70 15 85 55
 73 CD 16 67 89 0A 5C 58 88 BB 75 4B 5A 13 FF 77
 D8 D0 76 8E 96 6A 24 6B 05 C0 C6 EB 0A 06 7D 47
 6D 23 87 7D B9 1D 53 6B C7 32 51 38 BE D5 1A 2E
 75 68 DA B4 EF E0 6E 08 33 1A 89 29 87 E9 ED DC
 A0 CE 81 FF 95 4C 02 00 66 33 20 31 E0 27 51 1E
 EC FD CB 0E 58 E1 19 D0 6F D7 04 AB 8A 9D A9 E6
 E1 42 05 AC 82 4C 7B 24 1B 10 22 0C CC F2 4A 29
 63 E5 8D A7 86 4E B0 1D EA E8 59 53 7E EF 34 B1
 1F 1B A3 BE AB 34 8B 56 8B F1 4D 90 11 04 75 EF
 5C B4 B6 FF E7 81 36 45 85 6E E0 7A DC AC 31 43
 3D AF 62 87 FB 06 26 E8 C7 A5 A9 8F 2D DB F1 53
 5A 20 7D 13 B9 0C 1A E7 6E 2C BD B1 86 BE 42 9A
 6B FB 5C 67 71 01 C8 D8 CB 17 F8 42 3B DD 27 12
 A4 5B 11 DB DF C3 3C F5 A5 BE C7 E4 E9 0D 6D 90
 2A F0 44 B8 4B 19 EC 13 F3 C3 4D 13 F8 79 3B 7C
 19 3C 84 5B 26 5C 15 7B 4C 62 35 85 B3 6F 01 56
 4A C9 2D FD 5F E3 22 53 FE 53 F0 A6 2F 2A FB E9
 55 F4 D5 79 BA 55 A1 5C DC 06 1E 65 07 1D ED 82
 39 5A 69 55 03 F0 7E 81 3A F1 59 A7 AB 86 13 1C
 4F EA 8B E1 63 27 5C 4E 6F 58 0A CD 58 AD 20 85
 7D 46 A7 15 C9 E2 84 2B A4 50 69 BB 7B 48 59 A3
 BB 9B D6 87 F9 95 FA 0C BA 54 D6 7E B9 F6 31 2A
 56 E6 7C 3E C6 24 70 C4 48 24 7C E9 4B 01 57 AD
 00 4B 6B B6 78 ED E7 8B 73 95 BB EC 4E E9 C2 AF
 F7 E2 2E 4D CA CF AA B6 D4 4E 09 F1 26 C4 77 D5
 87 2D 1E A7 EE 45 34 F8 36 D2 C4 D2 4D 93 5F AE
 8E BC 5C ED D7 77 6C E1 6A 39 22 AD 6B 8A 5C 88
 8F 91 D5 34 ED 83 61 D4 8B A4 2F 2A DE 32 B5 35
 23 97 87 46 C4 A6 72 BA 77 AC 54 32 91 F9 C5 E8
 51 0A 0C 95 DA A1 90 20 00 11 A2 6F 31 71 61 BD
 79 91 83 8C D5 B5 18 E8 6E E3 DB 96 23 0D CC B5
 C1 3F A8 B8 EA B9 D4 F1 45 6F E4 E2 4F E5 0A 8E
 81 59 01 E2 DF 44 54 38 FF 9F 37 2A 20 47 96 65
 02 02 CD 8A 14 28 2D A7 D0 98 74 38 CA E3 67 35
 FC 88 21 C2 E1 8D 5B C8 E5 E1 D0 03 63 05 7F 3E
 1C 2A AF 8D AF C2 EF 9E 4C 45 BD D2 6D B9 6B 69
 4D A6 5C 7E F2 73 D6 76 C7 94 DF 55 3C A7 B6 C2
 6C 9D C2 4F 8B 6F 01 3C DA 45 73 A2 9E DD 1A CE
 C4 07 C4 4C 1E CC F9 FA 1B 1C 8A 25 13 D4 E9 CC
 5E 39 E2 82 CA 03 FB 42 03 90 D3 74 17 74 AF 6F
 3A 28 F9 33 B1 42 0C 3B 6A 87 B1 48 6E 46 C7 D6
 2A BF FE 45 28 62 E5 79 07 AE E5 0A 8A 6D AD 06
 2C 20 04 43 42 BA 4F F2 2D F5 7F 13 B8 61 47 7C
 99 95 17 94 4F 2D 99 10 78 C4 A1 87 D5 A9 A7 96
 DD 7D 32 EB B6 8E 08 B5 8C A1 BD AB 8E 8D A8 50
 CB 3A 4E 74 5A 1D 99 27 60 43 AE B8 36 1A 0B 05
 E3 DA 90 D4 7F 24 5B AD C7 64 85 09 0D D9 71 9F
 14 8E B1 E2 F2 22 62 55 37 57 F8 8D DE B3 38 EC
 07 CB C2 26 8E 0D 85 94 62 A6 5B 19 C1 14 F6 E7
 DD C8 8A E1 BF DB 47 1A 71 93 E7 98 11 11 80 E6
 38 98 4B 60 C5 A8 D4 2B 68 17 98 40 1E C2 AF 15
 0E E3 5E FD D9 97 08 FB A9 23 5C 53 2A FA B1 6F
 C6 BF FC 8E A2 72 BF A0 BE 53 ED F0 9F D3 4E A6
 6B 78 DB 56 29 ED B6 08 15 FA C1 E3 7E 2F 3A B1
 8A 17 AE 02 F6 8F 37 DE 3F 0B D5 41 61 A9 B9 22
 58 A5 72 54 E4 AD B9 C9 83 5D 4F 1B 2D C7 FF 08
 B3 6A 16 FE 6C A8 B8 40 66 44 96 7B 59 01 60 25
 2E 22 C8 B6 31 64 10 43 89 7A 1C 2E 2B CC 00 AB
 8F 3A AB EB F3 0C D9 08 8A BB EB 8F 10 71 8E 34
 6D FC 2F 73 55 E0 16 65 36 48 50 9A 00 71 25 66
 BD 0D E1 7C CC 28 61 7D EF 18 A7 1C E5 3A 7F A3
 13 39 63 63 68 25 91 FF 13 79 75 17 56 8D 27 2F
 7B 19 C7 88 4E 5F 75 64 52 7F 80 7E 49 90 00 B1
 5B 57 F0 3B CB DC 2E 4C 44 A2 8C 23 A6 A2 C1 BC
 8D 63 BD EA 99 97 C0 04 4E 3A 69 8C 7C BC 41 1A
 5E 4D 09 8D DE F9 CC A5 79 0F 97 57 7C 5B 88 91
 41 D0 F3 D7 84 14 3D A5 C7 79 58 D0 73 3E 67 23
 16 D0 D5 1A A2 EB D2 1D 31 E7 B3 F7 36 A9 75 29
 1A D3 CB 44 06 20 A4 99 1A 86 77 13 B9 F8 A4 B4
 DD BE B7 69 B8 81 73 15 10 D3 B5 C1 8C 81 25 A2
 DA 62 DD 02 E3 4C 31 E0 3C F2 99 1B B3 5D AE AE
 BF 2A 91 33 F3 0A 6F 95 CA 1E 66 97 1A 7C 88 94
 18 DC EF C9 B0 E5 FD 4E 16 0F 6A 67 9A 51 D8 88
 2F E4 22 0B 16 43 43 C3 C6 B1 12 51 D5 E2 16 47
 6B 10 E0 1E A2 4E D3 F6 46 CD F8 1F A2 DA 11 CC
 53 BA 12 D6 F8 CD 69 86 51 04 FA 45 C5 17 F9 A9
 CE F0 9B F9 0D FC B0 45 06 87 79 D6 54 D9 43 CD
 1C 96 BB 15 33 8B BA 8E B3 00 12 54 B0 2A 19 A5
 0E 93 A8 FF 3B BF 0C BA 65 DA 0B 64 5F 0B CA 3D
 FF ED AC 30 DF 89 EE A2 DD 28 18 04 E6 E7 F0 46
 B6 D0 C6 5C 19 46 96 82 49 CA 27 ED AF 6F 13 0A
 DB CE C0 98 81 06 6D 7D 07 BD 7F B9 0B 02 6A DC
 F0 C8 74 8E 4B 08 0E A6 F9 14 82 65 4C 5C 25 4C
 36 1F B2 FD 00 81 AB D5 0F 11 97 71 39 F2 13 8D
 70 7C 9A F7 F8 6F ED 20 6C C6 27 F5 64 C2 4C 70
 BB D4 AB C2 79 ED ED 4E C0 C1 95 BC 11 4E 9E 89
 7A E6 4B 42 AC DE 86 E9 46 18 27 02 DD D0 EE A8
 8E 75 6E E2 8E FC B7 3D B0 10 FC A6 5A 7F C5 60
 E2 3F 86 30 A0 83 72 C0 06 97 5C 5C B9 FA 5B 10
 B8 D2 26 A4 44 10 BB 75 81 8F 48 AC 87 69 86 CE
 F1 8C 2E 87 07 EC 9A 37 D4 88 E2 FF 67 3A 85 5A
 70 E8 00 32 73 DB 06 AC FC CD 0A B3 57 F5 83 FA
 70 F4 EA 92 29 BF C9 FF 81 A0 56 FD 0A 9B DB CB
 FA 54 19 C6 F6 86 EC 34 20 3D 15 70 9D 53 55 FF
 8A 35 84 76 A0 82 C4 6E 5F BA F7 41 7F A2 03 9A
 62 B8 9B 5B CB 06 2C 1F CE 16 ED EE 63 5A CD 44
 39 85 3D F1 4B 87 18 8A D9 AF CD F4 02 5D 6E 77
 73 1A 4F 77 1A E6 DF 48 D9 A4 8D D0 32 31 7D FA
 CB C5 D1 02 85 78 BE 35 8D D4 BA F2 A3 84 BF EE
 D7 37 FE 76 7F 17 32 A7 79 D3 97 33 55 A3 7A 89
 92 18 2E 84 C1 6B A7 39 F9 49 24 8B 2E 2C ED 63
 A3 06 67 B8 10 5E DA 3F 14 02 47 90 41 82 71 30
 4E AA E9 FC 9F 45 7E BC 05 66 08 A4 A9 B3 49 69
 86 3E 3C B3 8D 71 1F 2C A6 48 49 EC EA B3 D0 86
 8C 2A 40 78 D7 90 80 ED 4B 99 87 AE CF 4F B5 95
 68 A6 31 2F A3 B5 08 CB 76 45 44 C1 9B 6F 5B B1
 AA 41 16 20 97 EE 6F D3 6C 88 83 92 77 21 B5 7A
 C8 EF 6C 03 DC DB 45 8E 6C D2 67 2B 7E 47 AF EF
 13 ED D8 2B CC 62 AC FE 18 2A 1D 1B 98 42 A4 7F
 3D 8E C7 48 31 C4 1B BD 97 FA F0 55 67 54 4E 9D
 48 FD D3 20 04 66 BA 96 DF 95 A7 43 07 9B 22 65
 C4 C9 33 74 B5 04 6B 43 21 AD EA DE EA D7 19 B8
 0C 71 EF 4D D1 15 F0 2E 65 F1 36 63 79 16 A7 49
 66 35 B6 A4 E1 C7 1F 3D 35 11 3C 2A EB E1 69 7A
 0B F0 E2 FA 85 10 2C FF D3 F8 42 3A 37 E1 0B B2
 28 6A F3 BB 89 AA EC FC 89 34 83 B9 FF 4A 20 02
 C6 8B DC 69 70 67 63 49 44 6F 55 33 F1 EB 94 7B
 69 8B D9 AF 9B BE 35 6C 14 CC 29 BB 1E 0F 8A 82
 CF 2A 32 CA 16 DC 04 81 1D 90 CD 1D B5 1F 92 8D
 FF 00 34 6F 26 36 6C DC A1 3B 66 47 8B B0 A4 41
 79 8F 0A 50 08 5D 80 E4 9C 82 93 2C 8E C9 F4 64
 8C F2 CF 36 BF 06 4F 2F 6B 51 A5 FF 18 C2 2D F3
 13 ED 7D 72 B7 1B C4 39 81 2C 45 7F D4 EC 90 71
 33 5D 86 34 E2 65 91 CA A4 FE 61 C8 39 7A 7A 60
 20 A0 9C E9 D4 88 6F 1D 74 CF 33 B0 D6 48 E7 5B
 FA 64 9D AB 50 92 75 01 28 BB A3 36 FE 04 A9 2B
 CC CF 43 48 E9 B3 A1 EC C2 D8 58 64 FD 56 91 D4
 42 A8 4B A9 88 29 E7 50 7E FB ED F0 AD BB A2 BA
 D1 CE AB 5B 5F B4 C1 9C DA FB AA 1B FE 2E 06 26
 BC 6E 6D 88 6B 58 6D 7C 84 97 BA FB C4 1B D5 7F
 C0 85 51 21 FB 83 F1 1F 6D A3 08 41 C6 68 12 5E
 CB D6 8B AA 20 DA 75 CF 4B 9C E1 A0 F9 D1 80 54
 7D 37 83 6F 01 DC F3 4E 8F BD 0B 74 24 30 2D 75
 EF 30 B7 E9 3B E8 EC 8C 6D EE FB 8D 97 F6 D2 2F
 31 30 8E BA 2F 43 29 59 8C 51 77 07 BE 85 7C F9
 35 71 41 4D 4C 32 07 A1 3F 96 3B E8 C2 0A 9D 71
 2D 78 52 E1 1A 5D 4F BE 1F 8A AC 83 6D FD CE 9E
 64 C1 A3 6B 19 3E D6 F4 71 7C B2 E6 E2 3A 5F 82
 3C 9A B1 F9 1F 4F 40 61 34 56 E5 CB 16 98 D2 0B
 4D 53 04 3C F0 71 F6 42 83 4D A2 8E 30 A7 3F B1
 5B 7F E3 CF 44 0E 57 4E AF 62 F9 88 0D 5A 2D 44
 F7 A9 E2 4B 4A 06 AC 93 EA 12 A0 12 C9 28 C9 56
 96 9F 7C FB 1C 77 61 EC 15 B0 6A 62 FB DF E4 30
 C8 32 57 CD 31 82 7D CD C9 2D F1 DE 45 63 88 A3
 3E 20 E5 6F 68 5B D1 33 67 A2 E3 6A CF B1 AF 86
 98 17 FF 79 0E 18 29 19 CA A3 30 77 6D BF F8 64
 B0 F2 4A 69 FD 72 BB A5 51 65 A5 34 EF 33 D8 E5
 05 8F B4 35 71 F2 12 CD 87 D7 AB 8F 74 B8 C2 B4
 2B DE 28 7D 8A 66 99 8B 95 19 77 37 A0 65 92 A9
 22 80 2E 6A ED C1 3D BB B4 FE DF B3 5F BA 96 D5
 7D 1D FF 1A 28 AF 57 26 07 80 48 4E 40 5B E7 DB
 1A 4D 26 7A E0 AB 8B 22 DC 6A CB E1 F0 D9 17 34
 13 A7 E8 F5 AA 4F E0 DD F6 DC FF 5F 78 CD 99 A0
 44 8D 77 6A 3D B3 81 6F C7 D6 3D D6 12 EF 0E F3
 3C 89 80 69 F2 4E CA AF 79 0F C1 55 09 69 63 CD
 92 E1 96 E7 AD 51 89 00 20 A1 7E 8B 35 3E 0C FA
 A2 A1 0A 4D 1C EF EC C0 D3 8E CD FB 40 86 1C 7F
 1F 64 32 D3 5B 7C F3 D4 13 74 FD 05 75 AC FF C7
 77 04 B1 A3 95 A2 AC 0B CD F2 7F 46 81 5B B2 CB
 FB 6F 92 C0 AE 68 7A 7E 10 88 FC 48 8C 15 F0 36
 32 20 40 A9 98 3C 0B 42 D4 8D 92 F2 88 01 04 65
 7D 7E 9D D4 C2 30 04 38 99 29 A1 F6 C0 91 0C AB
 D2 6F C3 71 35 60 F9 F5 83 A1 71 83 8B C2 5C CB
 F6 D5 A7 9C 98 3D FA 45 A6 8C F6 D5 62 22 45 13
 3E 53 60 EB EF EF F3 30 F9 50 23 E8 52 EE B9 C9
 FD 2C E5 86 C6 7B FC 73 F0 DD 8F ED 27 A1 0B DB
 C8 2D 8F 16 64 D8 DB 8E 18 7D 57 B8 EC 93 46 F5
 36 88 94 28 77 AD 34 46 E3 5D E3 B6 30 8E 6A BD
 F3 46 60 4C 99 76 01 2C 68 D7 D2 B1 28 6F A6 05
 C0 C4 32 2E 41 6D 42 76 2E 88 D1 CB E6 A5 BA FF
 56 D4 EC 5B 30 05 92 50 93 D0 9D CC 4F 8E 08 1C
 67 9E D0 DB 3C 27 E2 9C 3D 3B 78 74 7F C4 05 54
 38 9D 14 E5 67 82 69 7B 3A 4A 34 33 33 C6 FC A6
 99 2C 8F C1 B5 2A 2B 27 4B 98 F7 17 95 4D 9F CA
 2A F1 6B BE 98 17 47 09 D8 F3 A1 AC 02 D8 8D 10
 04 60 00 27 01 E1 E4 BF E5 6B 80 E1 20 57 F8 1E
 A6 74 46 08 E1 2B 05 CA B6 B4 C8 CA 10 CE 84 BE
 2F 2A 29 42 A6 62 CE A3 51 7D 3D 84 41 70 2C 7B
 D4 AB 3B 66 5B 75 AC AA B2 FB 4E DB B6 46 1E B6
 8D C7 29 02 48 45 32 DE 40 01 CC 75 A8 D5 98 89
 16 4E 74 3F B0 C9 D5 0C 81 AA 62 FC F1 00 08 43
 C0 BA 4D 43 FF DA 31 9A 6B 4B 17 87 CA FD 09 4F
 7E ED D7 23 59 E7 12 D2 C0 F6 77 EF 6A D7 5E DF
 CC 97 36 56 44 F9 9C 57 F0 80 67 3C 40 E0 8D 72
 CB BC 1C AF A8 11 32 2B 30 92 E2 1A 25 26 29 B4
 05 40 02 75 12 13 B0 B9 B9 3F 44 28 83 F7 4F 42
 48 86 8B 72 A9 A0 63 25 B6 46 C5 24 7E 5D 2D 90
 B6 96 AA 08 79 FD BD E2 D6 6D C8 2B 79 C6 BD 54
 1D F5 50 ED 26 C7 61 58 6A 0A 0E E5 69 E1 62 98
 50 D7 C4 0C 6C C0 9A 66 29 9D F7 10 57 FA DC 38
 35 A7 F7 1C 44 E1 99 35 09 1F 95 89 FD 2A FB 5B
 EF 4E 04 BB 8B FC FE 1B 45 7F B2 DA A0 D0 28 85
 3B 54 75 25 59 59 17 41 B1 94 0D 86 19 11 87 8B
 E0 60 C1 68 6F 72 5B 6F 7D FA E9 F1 4E A4 13 CA
 73 8D CF D5 D2 93 A0 9F 29 0A 52 AC 0F CF F9 ED
 96 E1 67 77 9A 2A 99 B8 A9 5D 98 A0 25 75 EE 02
 12 E2 37 EB 50 B4 E6 91 2B DA B8 A9 49 36 2F C6
 2A 5B 96 2B EF C8 89 FC D6 8D 25 53 F7 C5 B9 B0
 82 FC AA F9 AC D9 F8 B3 7A 0C 1C AA 77 9E 06 CC
 C2 B0 14 C3 97 E0 BF C3 2F 20 B8 51 C7 17 F4 0B
 B4 77 60 8F 3B FF CA 3E D9 25 7B 67 8C 7D 0C 07
 53 21 18 AD D8 61 A5 D0 E5 00 79 82 95 70 1A DB
 06 F4 52 5C A6 E4 80 61 01 CA 18 C6 BD AD 80 75
 33 A1 28 D7 2A 34 B3 C2 B3 A2 E9 08 AB EF 28 47
 D7 CB 85 00 4F 5D F4 A7 CC 37 0A CD 3F 53 EF B7
 8D EF 28 43 93 0E FE 48 15 C8 B8 F6 07 6C 1A 57
 6E 07 82 AB 32 F8 63 EA FA 0B 15 DC EA 55 F6 48
 B5 73 0F 13 B1 1B 78 E4 03 22 75 EB B4 A5 D8 F1
 8D C2 66 F6 99 D7 0D 32 6D 2C 2A F8 54 C9 7D A8
 BF 49 18 E6 FD E7 8D A2 31 A6 83 9F 89 BA B5 E0
 0B D1 1E 88 88 59 C1 D5 E6 D7 8B 61 CE C2 9D 3A
 FE 74 9B EE 20 C4 3A 34 9F 68 D2 2D C4 1F 0B 53
 C5 AE 67 26 C6 7F E7 B4 22 51 9A 69 2B FA 4D BD
 2E 0F DE 44 09 1C 93 92 40 56 34 6E B2 3D 11 20
 92 6C 5A 25 A7 2A 20 9C 14 10 4B 4B ED 3D 30 39
 36 49 F9 28 F9 ED 6D FB 85 EC 62 17 38 A6 B4 24
 08 9E 6A 07 97 47 D1 2E 48 AB 12 B4 EE 3F D6 15
 3D 1F C1 E4 C1 3D 25 0B 5B DE D4 3A 90 DF BF 16
 A2 04 EF 34 34 D1 A1 2D AC C5 0F FE F3 8D C5 4B
 1A 29 46 A3 43 21 60 32 6E 22 AE FB 98 2B F7 65
 FB D4 90 89 54 7D DA CE 1B 0D 8F 78 78 03 63 F7
 35 F8 46 E2 87 13 06 71 9F 65 CC 44 5D 88 66 FA
 13 2B AF A0 38 53 8E 75 D2 EA DC 0E 9C 22 07 A7
 7A B6 98 4F 46 29 0D 91 5F B7 05 D6 F0 B5 E6 3E
 A4 82 F8 3F 5D BF 92 80 CC 78 86 72 F7 92 39 34
 33 C6 30 16 99 A4 07 79 24 F2 67 1D ED 61 99 EF
 2D 16 93 DA 2D 67 B3 00 CC 25 4F 07 FA 1C 85 8E
 DD B5 C1 F7 88 08 BA 93 10 03 F3 56 E1 CD 3C CE
 5B 15 C1 44 4D 6C A5 57 44 47 AF 4C 36 B1 A0 95
 E8 C4 FE 94 C5 03 A8 BF 51 36 2A A2 E6 02 E0 62
 75 E4 10 BC A2 2F 0F 5C B5 01 5A C9 4D 7A 2D 0A
 08 65 F0 D9 54 30 0A 8A 21 09 23 AF C2 81 80 73
 4A B2 90 DF FE C0 11 3C 10 4D 11 67 3D B1 1F 45
 2F 52 87 88 26 0C 73 61 C3 41 4C 34 4E 11 C3 BF
 ED 21 FF 1A B7 48 79 C8 7F 3C B2 E9 6D AF 06 83
 61 05 DA 98 35 0A 49 21 50 29 3C 03 0A D1 B4 C7
 9B 80 98 62 AD F9 86 54 FF 23 0E D3 17 9C C4 20
 82 DA 98 5C C8 B3 36 A6 A7 F9 04 BC FF 6A DC F1
 09 4B 8A 9B 5E 4C BC C2 2E EB BC 4F 1C F7 CD 71
 12 B7 BF 2D 3C 50 6B 37 4F 5B BC FC 1F 90 51 BE
 74 8D 93 38 54 E1 F2 ED 04 F7 CA E0 D5 75 C8 5A
 44 42 E1 84 3A D6 DD C4 0B 89 FC A8 35 ED 48 43
 9D C2 9A BF C2 50 0C 89 E8 11 CC 78 20 72 19 87
 CA CE 17 5F BE 35 EB 1A EA C1 E8 D4 0E 7F F5 90
 07 F2 35 77 B4 52 5C 9B F7 44 24 26 FE 63 18 C3
 18 5D 09 45 70 43 6C AE 68 A7 93 CB BD 33 EB 75
 FC EC D0 8A 82 B2 97 A3 08 28 48 A1 53 E4 DF 8A
 8A 39 03 8A D2 02 DB 99 B4 B4 04 84 69 19 AE EB
 2A D3 24 D2 85 B3 D0 2E 43 7F A3 32 D9 F1 D4 83
 48 2C 2E EC EF D0 D2 23 F3 9F AC 3B D6 95 C2 F8
 DC A4 DD 17 E2 91 DB 8D 08 F9 1A 6E 74 99 85 04
 73 F4 BE 18 76 40 2F 0B 14 B7 F9 7B A2 15 91 3B
 2F CA D5 EE 56 9B AE B5 96 50 F7 BE F7 2A 4D 93
 68 E3 91 66 3C 56 FF 43 BA E6 27 EA 84 80 F6 C5
 52 76 0E 67 75 DE 29 AD 94 D1 24 C5 36 BC D6 EF
 CC 7D B7 B8 DA DF 6F D1 37 B9 1A 7C 15 C6 2C A5
 3D 0C 07 9C 84 19 EA B2 D7 A8 E7 C8 B3 90 A5 FC
 29 5A 02 09 CC C3 1B D6 48 A2 DE C5 F2 91 75 00
 41 E5 EC AD B5 B9 E9 6B 21 BB FD 9A 73 E5 5E CA
 3A 5A 47 8B 51 40 68 6E C9 4A 82 43 C2 8A 20 91
 B8 A5 D3 4E 0A 71 7D D0 96 D9 3E CF 12 16 DE 24
 6A 75 81 1A A1 5D 46 39 AE 47 D8 F5 AC C6 17 46
 D4 8C 59 96 7F 5C 7A 9C C3 D6 53 1A B5 BD 85 93
 2F 23 9E 0D EF 1F 6A 54 65 D1 1F F7 64 68 8B 21
 8B 40 FA B3 75 1E FB 5D 17 BF B1 79 C7 61 34 D3
 C5 B8 71 41 56 9A E3 82 11 B6 BD E1 A4 F2 3B F0
 1B 12 B1 A4 83 DA 46 B3 8C 9D 49 38 57 6B 97 64
 8C 56 46 FA 7D C2 19 B6 4A FD D6 6A E3 D0 71 F2
 AA 3B 3C CA F7 F9 77 BC 56 23 C0 77 A1 BD F7 12
 92 DF C8 09 86 5D A0 37 4B E1 E2 BF BD 9C 25 18
 19 CA 0A E7 BA 4B 24 BF 0E F0 BD 9A 0B A7 72 B5
 C8 B1 7E 40 F1 22 EB DF B8 B2 86 37 02 C4 74 54
 10 21 94 66 B7 67 BB B9 89 FE 8A ED D5 55 DD 0B
 6F 37 17 D5 E4 BB 46 E0 02 AB 6F 5E F9 EA E5 B8
 C5 AA 5E FA 51 5A 8D D7 BD 74 F4 9C E8 4F A3 5E
 C9 C7 C7 AA 62 6A 10 7B 2B B1 08 00 02 3F B1 3E
 8F 9F D1 71 03 F5 B8 A5 5D 23 63 B6 E7 2A 85 D3
 6C 10 5E DB 55 FD BA 73 2F 2B D2 5D 18 B1 19 51
 20 A4 F6 B7 99 EE 07 F3 9E 26 F6 C0 45 72 08 C1
 2B D5 A3 B6 D5 F6 7D A7 CD 41 B3 CB 33 1D 75 05
 AC 57 06 32 A5 54 E4 27 E1 C7 C5 A9 F8 AA EA 54
 6A C7 1B 77 BA 7B 01 CF 68 88 DE E8 A2 50 82 DD
 96 A4 4B AF DA D0 2B 1C AB A1 F1 5D FE A6 8D 58
 84 53 00 BF C0 6C 94 A0 B5 C6 92 18 3D 7D AA 25
 E8 69 11 FA 55 93 7E 23 62 F8 21 C8 30 2B AB 4C
 3B 13 FC F0 9D 84 AA D1 B9 71 3D 67 1E EC 65 E1
 2E 2F DA 7E 86 CB E0 04 A0 83 C0 E3 77 C6 FA 7F
 34 70 B3 89 B5 62 5A 1E E6 30 9C 3A 9E 5E C3 D2
 21 D6 76 09 A1 F5 F5 8C 36 D8 D6 60 88 ED 3A 46
 08 56 39 A6 A0 18 9E 0F E8 A9 28 FA 69 12 A9 66
 97 2A 39 FA 60 72 19 6A 1E 19 1E B9 CE 12 5B 4A
 FB 12 EE 5E EA F6 70 05 8C 46 BD 2F F6 DB C4 0A
 81 26 50 AB 8A AE A1 7F 37 DC C7 41 84 52 25 22
 DE 57 2B 6E FA 13 22 74 E1 8D 99 B3 97 0C 6A 6C
 34 91 7C 0F D4 75 29 1F A2 94 9D 73 33 47 14 D2
 4F 85 28 A5 F7 61 B4 C7 7C 23 A5 70 39 47 C2 94
 5D 0C 0B 94 4D C9 6E 80 92 49 CB 5A A7 0F 1F 8C
 6F A1 D0 8B 95 7C 68 05 EF FF E8 84 EA BB D7 B3
 54 4D 7F 75 83 A8 C3 B0 78 1C A6 8B 74 B4 E3 BF
 47 3C 6F E8 0A FB C4 C4 2D 58 3A A2 CD 57 FF D6
 EE A2 38 60 7C 5B DD 72 6D 77 0C 85 DA 54 64 76
 E8 94 41 62 36 FF 3A 0D E2 5A 06 B2 86 66 17 6E
 5D 64 62 8E E5 40 22 44 02 AA DB E3 90 F6 C1 CA
 34 09 97 E1 1D 01 10 E0 09 5E 06 4A 3A 82 D9 99
 E1 D8 E2 CB A7 8C 9A 5E 47 CA 52 15 1F 3D 00 E8
 26 31 71 38 4B 76 4B F7 A2 8E F8 98 53 99 47 75
 3E 07 29 16 E4 43 49 4F C9 DA 73 9A 6D DB ED 14
 DB 7D 83 F3 DD BF 3C 99 A9 34 23 51 9A DF D9 BC
 3E 21 37 29 CB EF 5A 82 B1 D9 29 5B 3C 18 AD 76
 AE 33 1F BD 0F BC B8 0F 59 A9 09 84 70 65 FA 2B
 04 E0 41 70 07 91 81 52 76 C8 8F 3E 34 75 19 1B
 12 9D FC 12 4E AC F4 85 58 A4 C6 1D 2C B3 A4 B6
 49 E0 67 47 77 F5 98 78 0A 35 6B F6 12 5B 6A 67
 97 95 E2 55 3E 36 5E C2 74 70 30 4B 92 0D 1A FB
 03 98 DF 24 B8 36 D6 1B 35 C1 04 97 34 BE EE 42
 BB BD 29 B3 8F 34 D0 4C 3B F1 34 4D 6A 82 C1 02
 A3 61 D7 F5 F7 B3 D3 0B B0 57 00 11 24 54 5E 8A
 CB E6 16 01 26 47 8A B7 99 9B DE 5B 47 B3 55 D3
 3A EF 6B CE FC 73 16 65 30 0D FA D3 99 65 C2 E8
 8C 56 F2 C2 AF 6B F6 05 53 B4 E7 CF DC D7 E5 44
 C8 79 D5 5B 20 F6 22 43 5E D3 98 4F 21 E7 10 01
 D7 55 B0 02 1D 68 F9 0A 4D FC 7A 31 F9 15 BA C4
 F2 E2 B9 C6 5F 80 66 8E A6 7F 22 7B BC 1A 7B 5F
 F5 BF DD 58 FC AF A9 5C 3C B4 45 AC 4C 2D F3 A5
 F3 B0 63 FE F0 D9 A5 25 DD 39 A7 D5 A5 E7 97 23
 76 E3 49 D4 6B 3B 6C 0E CE 87 D5 4A CC C5 E1 C9
 A9 91 B4 F1 39 E6 94 65 12 DF C2 00 B5 B1 38 59
 A6 5A CB 4D 15 B9 B1 39 B5 EA FF D1 CF B7 87 56
 B0 39 D2 1C B6 17 0D C6 4F 49 7A 79 C5 9D C0 68
 71 32 9B 79 57 E8 5C CD 3B B4 F4 D6 35 4C 55 37
 B9 2A C7 96 06 27 30 51 55 B1 FA 3D DA 8B 3D BB
 4D BD F1 66 F8 7A 32 9D 65 C2 58 2E 57 84 50 0F
 6A 3A CA FC E5 EB 02 A2 DC 60 79 EF FE 56 36 4A
 7E 68 0D 94 BD 6A 2A C6 39 85 AA 75 0D 34 43 8F
 9A AB 01 C5 7D 7A DD 88 B0 2E 7E 4C 35 BC 90 02
 3A 45 DE AB 59 FA 26 32 E2 8B 75 28 09 0C C9 F6
 72 8C 06 34 DC 45 1C FE 01 02 D8 BB C6 B2 C0 2D
 F8 83 5E 73 BF D2 26 EF FF FB 4A EB DE 7B 26 4F
 02 91 0B 24 83 C3 17 8A A6 39 1B 0A 49 D1 FE 93
 A8 D2 86 AD E7 B9 B6 5A CC D1 52 14 61 23 7E 72
 DE 33 40 C5 49 06 84 F5 78 0A 6C 12 13 CB 2A B3
 97 B9 6E 7D F6 89 CD 83 E4 FF 43 4A C1 86 6F 00
 00 03 19 B7 D6 37 89 9C B9 D1 94 D7 DF 5F AA 50
 A6 FE 2C B8 5D 4A 26 03 D1 75 F6 8C 89 52 87 30
 B8 BF CB 67 6F 37 F5 57 B6 B7 0C 78 76 06 81 E8
 F1 1C EB A0 A5 5C 75 FC 8E 0F 89 F2 FD 61 A4 EF
 25 81 24 43 C8 FA F6 81 64 D3 0D 8B FE A1 1D 75
 BA CD 82 28 33 60 10 1C 4A B4 13 CF DD EC D5 8B
 B2 7A EF E6 1D B0 81 35 8F 2B CF BE 64 A9 A8 6C
 D3 7B AB 9E E7 EE 84 A9 79 AE 3D 1B 8D 8F 50 E7
 B3 85 73 9A 13 A9 7D DE 35 FD 8C ED 4B 6C 48 E6
 F9 0D EA 5E A2 7C CF AF DA C9 A2 69 70 A8 2D DA
 4B BE 66 80 77 1F EE AC 2D 6E 1A 62 DC 90 63 F6
 F5 D6 B2 3F 38 B0 90 DD 22 EF 58 6F 73 66 AB D8
 A2 14 66 AD 85 17 B8 D7 2C B3 FF 96 14 00 CB E1
 00 CE 81 A5 D9 1E 3E 6B 3B 9D C0 42 17 91 DE 02
 BE 15 79 B4 65 40 06 34 8C DC F9 83 D0 BA 29 73
 15 20 B3 3E 79 CC E4 B0 4A 5A 95 FB 7F 33 6F D5
 4B 39 6B 13 1A CF 96 A1 EF 9A 8B BC 4A 06 AC 7D
 71 B7 86 6C E1 FE 71 68 6B BE 46 87 C1 20 DE 88
 B4 CA D8 14 21 D4 FF D6 4E 78 EF DA 6B 09 30 C9
 50 33 CF E8 E9 4A 87 DA 90 B1 C3 B1 B9 1C D7 A4
 83 C9 12 47 63 43 39 F9 03 93 D4 EE 8D D6 D6 FE
 22 C5 1A AB AB 6A DE 85 D9 45 F2 E2 48 0A DC CB
 D4 2E 65 A8 48 A7 D8 91 68 C3 47 2F 40 FF 86 B1
 4A 38 08 14 7C 96 C5 B2 20 57 70 39 59 0E 49 6C
 84 62 33 DE 2D D3 5C EA B4 B7 C9 E6 ED 8C 9A 1E
 61 E3 8A DE 30 FE 00 32 F0 44 9F 38 AD 1F 58 59
 FC E6 43 3B AB 74 5C B0 9B A9 64 8D E5 6C 30 DC
 2E 0F 4A 3F FB C8 E3 54 7A 35 F8 C2 58 92 D7 83
 EE 1F FB F7 DE 90 74 57 A9 4D DD AC A2 BE 0D A9
 73 F1 50 3B 72 10 68 9D 83 49 2A DC 6A 7D DF 25
 70 34 4C D4 4E F0 73 D2 E3 BA CB FA 56 8E 54 4B
 14 6C 12 AA 4B 9E D0 D5 44 EA A6 7B 26 72 0E EC
 FA B2 58 DC E6 A0 D7 63 6D 90 2F B6 37 EF E8 A1
 CC 30 BF 77 48 CC 38 9F 4A 7C 72 99 07 EE 29 27
 4E 8B 3C CB 75 7B 6E 2F 72 FA 72 1F F5 75 07 7E
 79 C8 A4 97 EF 8D 33 5A 31 CA E5 67 F9 CC 03 38
 E3 65 3E C0 26 50 D6 21 CE 0C 3C B4 E5 CC A9 29
 E6 18 7B 6C 7A C9 EE 07 E0 24 4B 4E 4F 92 D4 A1
 24 D9 BC 29 43 A3 80 FD 6A 6D F3 0E 0A 69 B9 1E
 69 3B 76 2B 53 64 4D 0C A6 AA 35 8B EE 68 BD F4
 1A 93 5D E5 FD 8F 36 8A 2B 8E 04 12 89 8B 1B 64
 AF 6D 13 B2 13 DF CE 4D 42 B4 5F 7D FC 6C 35 A8
 0D 40 ED A1 E9 48 B8 66 EC 32 15 75 00 21 63 53
 A3 6D 35 45 59 DB 13 F9 B1 A2 5B 58 7B 0D 33 0E
 3A 65 67 4E 16 04 AE 06 34 2E 0D F2 72 24 92 3C
 94 C7 57 07 F6 FB D0 70 CB FB F8 D2 C7 F3 7A C7
 D1 90 1D 44 48 15 49 D6 25 05 81 A7 FF 43 CC 15
 1C E8 B6 57 D2 FA E0 BA BB E7 2C 45 18 33 7E 22
 83 7A FD 9E 27 A2 11 63 48 FA 92 90 02 1B 93 E9
 60 05 E5 A1 43 66 17 80 30 4B EE C3 70 74 8B 04
 BD CE BF DF 41 E7 CC 68 47 F2 55 84 E0 D7 E8 72
 36 41 CA DC 89 24 CE 38 C6 8E 0A 09 4A C2 32 14
 9C AE FC 2F 1C AF 41 19 31 99 08 88 F7 3B 6C 31
 B1 07 D4 32 5D 2E 7E AF 51 C7 37 EF 22 4E 28 9C
 57 DB 7D F3 FD 2C 01 E3 0E 56 78 ED 85 09 7F 01
 6A 5B 79 D3 94 1E 99 E2 A9 B2 87 2F B4 AA 08 3A
 2D 79 93 90 1B 4C 3C 29 1A F4 F0 92 E6 66 7B 8C
 F9 75 85 E3 57 82 A8 05 16 27 28 5A 13 E2 73 4C
 A0 B7 7D EC 05 CC F4 04 17 28 84 4D 40 92 E4 D4
 B0 79 34 EA 6C 7D 4F 19 79 54 40 C3 90 F2 20 53
 0F 6F CF F2 B8 9B 73 B6 0A A2 C5 7F 01 50 07 8B
 1F 97 B7 FA B5 76 39 BC F0 04 E5 3E A2 FB ED B2
 69 DF D7 DF B2 DE 9C 9A 4F 96 B4 F9 68 76 28 C4
 4D F8 0B B8 89 DD CA 7F A7 DF 9C 6A D1 2B 50 44
 C5 0C CA 76 59 DF 0D ED 89 FB E9 18 D0 56 6F 17
 0B 10 03 E3 66 7A A8 D2 84 79 25 1B 1E 6F 3F 81
 F4 5F 0F D4 99 26 B4 13 42 E3 7A CC 46 C7 D1 AF
 E4 08 87 AD 04 45 DB 42 63 F7 D8 94 3C 42 B0 B8
 91 A6 53 53 FF C3 31 C7 D3 FE 66 72 4B 26 F0 DF
 30 00 50 B0 81 2D F6 84 06 2C BA 77 2A E0 E3 FF
 5B F8 51 78 71 B4 18 00 06 C7 C8 8F 33 86 4C E2
 32 AE 94 B3 1F 50 6E 71 B6 B1 58 AC 48 F4 FB 4C
 2F 01 4F B0 AD 17 EA 59 16 24 94 9F 02 74 C9 AE
 8E 75 DB CA D2 6B B5 34 10 1A DD 33 1D 83 00 58
 5C A1 E4 6A BB A6 7C 2E A2 59 2A 83 12 5A 4A 4D
 DD EF 4A 12 54 57 D8 45 2E 8C B9 FF 65 BD 74 7D
 D4 92 F2 C3 72 9C DA A2 FF E1 D1 41 CE 5A 85 10
 80 C6 74 93 F5 30 F8 EC 8D 5C 78 68 D3 3A B1 50
 41 86 FC 44 25 26 20 A3 F5 61 49 A0 DB FB 92 BA
 92 2E AC 27 2B B4 7F E8 31 1D D0 53 08 18 C4 20
 40 58 A5 64 3A D7 0F C4 86 AF BF EC 49 AE B3 B5
 2F 5D A9 9E 27 8C 10 6E F4 8B 89 A7 62 00 ED BE
 85 12 D2 3E 12 4C 94 BD 05 03 CF FA 50 A5 C3 D0
 61 08 1A 0C 1F C4 70 62 DF DB F5 F0 64 8D D6 5B
 66 A5 C8 F1 BF 57 F9 52 17 78 FC EB 08 D6 58 FA
 84 6C 3F DC C5 CD 5D 45 BB C6 BB E7 6F B7 84 02
 B5 CF 6D 02 0B 08 20 EE 81 11 4B B6 41 3A AE B5
 2D 33 60 4D 81 D1 E0 AF 68 7F 10 20 D9 BC 82 41
 EF A7 43 FD 7C 32 AB 35 FD 69 7A 70 2A AF E6 B7
 A8 45 63 2F FD A1 83 17 F9 C4 E2 28 D8 45 0F 97
 47 0F 84 0C C1 CA 44 34 C6 2C 52 91 D8 8A 77 D1
 E1 B3 D2 5A 0F B8 B5 A0 F4 91 6A FF 45 BC D6 6C
 2B 81 4B FF FE EE BD CB D8 90 AF D3 8E 28 B9 D3
 2A 2E 5A 70 9E 54 FD 07 86 B4 C6 93 A4 DF ED FB
 D9 43 46 9F 59 CE ED 4F 87 60 15 B2 A5 CB 4C 63
 AF E1 B6 E1 99 59 5F A3 A2 90 54 4D EF 38 F2 07
 21 F4 B3 3B 5D 65 3E 72 CF 58 12 7F 88 AC BF 30
 33 22 32 C0 3F 20 F7 03 07 EC 65 FC 68 10 BE 92
 26 21 E0 FD BE 02 86 B0 3E E0 D2 02 2E 6C C9 93
 94 AA 46 31 F2 4F F0 93 48 CD 55 A3 9C 8D 45 BF
 37 0E C6 04 BF AB EA 67 44 F3 15 70 DE 18 12 B4
 BF DD 2F C5 9A 82 9D 3A 9C FA D8 8A 35 CB F5 17
 00 22 BE 67 C7 36 DF B2 33 27 C3 F9 31 F6 B8 9A
 CB 6D BE 74 19 DC CE D9 46 B6 26 EF 3A DC 28 9F
 53 26 50 A5 82 37 2E A9 6E D1 EE FE BD 10 F1 AB
 A8 15 64 CD F5 38 CA 3A 86 78 0B 91 A3 6F BE 6C
 A0 FE 6B CA 74 68 B0 D0 F0 93 B5 BF DA BE C4 94
 85 45 5B DE BA BE 78 04 1A EC C3 79 75 56 9C BA
 D9 09 63 D3 F2 4B BA 1D 62 E6 B9 60 88 E7 68 17
 C7 78 CD 46 1D 9A AD 52 86 54 8C DF 86 89 0C 1A
 7B 2A 3A 30 CA 6C 3F 91 4F 01 76 A6 A4 01 44 6F
 FA A3 EF 70 CD A0 51 76 7E 19 70 1A FF B7 F0 D2
 8D E2 11 31 2D CD 05 5E 42 FE 97 F8 3D 01 D7 C1
 A9 2B AD 2C 3B 25 1C 79 F4 E2 5B 81 E8 A7 24 A5
 C8 29 88 5F 82 56 8B 63 5B CA F5 E8 9B 17 A6 E1
 9F 84 AF 3D 90 79 1B 25 47 ED CC 00 EA D9 1E B5
 1B 33 F4 21 5E 25 FC 77 C7 F5 EC 4E 1E 2B 6C 51
 29 80 99 27 05 17 B0 49 98 CE B8 59 D9 5E 4E 25
 CC A8 6C 5F B9 E8 28 83 C7 84 C4 7E 0F 4C 85 36
 DD 58 FF 22 EB 46 EB 54 60 D4 5C 6D 2A D8 BD 7A
 0A 2E 4F 86 2D E1 EB AF EB EB 4F E9 5E FD 19 B2
 77 FD 81 4F 25 EA C1 8A 26 A8 29 C3 5E 8F 83 E6
 D5 E7 3F 97 AF 81 7C 46 51 78 75 12 17 7D 02 9A
 35 22 54 E2 E5 99 7C EE 48 B4 C6 00 8A 45 D5 63
 EB 93 5E 62 58 E5 A7 8D 0C 3C A0 7E DC BF CB B5
 0B D3 78 FA 4A A8 A8 2D A3 A7 E7 58 C0 C5 40 4F
 26 CB 5D 2C 85 13 EC FF 8D 8E D5 50 5C F1 5E 07
 8C 10 FC 6C 6B 83 DC 66 EE 12 7F 76 89 B4 73 98
 07 05 52 A7 0E 38 FC 4F E4 54 77 4E 8A 52 5E 0F
 8F E5 76 C5 D8 9F 34 5C 73 20 EE DE E6 00 A9 76
 34 C5 68 69 3F 62 6C DF A8 17 EF 73 D2 D7 37 E4
 E0 50 D2 1D 41 65 B9 25 82 DC 8D D7 1F 2D 51 C8
 86 B6 8D 35 B3 4E 4E FF 72 AE 89 24 2C 43 77 39
 FC 08 57 8A 1C 74 51 33 40 DB 85 6C 02 C2 F0 D7
 2F D6 97 8E BB 4A 1B 4E 96 4F 3A 2D 78 E1 F6 AB
 8C 4F E0 24 E3 6F 0B 5C A0 38 2F CD 75 EC 9C A8
 6D D4 4F 00 FF DF 41 E3 E8 3D 45 BB F0 D8 3C 4A
 FD 4C 7B 73 40 17 75 51 1F 71 AB 27 B3 19 92 75
 49 8C 1B A4 28 7C FF A0 9B 49 3D E3 3F 15 52 0A
 6A B4 1F 0E FF 7E F9 5B 40 2E 90 AE FA E6 CF 83
 18 14 BC 19 53 50 57 FA 75 48 B5 11 E0 18 A7 93
 CF 7D 45 A3 23 87 AB E4 93 9B 44 CC 45 F3 F0 1A
 1C 81 A7 9A 8D 42 94 99 AB FA 52 85 91 BC B8 9C
 EA 95 1F 8D 10 55 28 E4 60 67 D7 D4 50 70 01 D2
 AB 83 B3 93 71 60 5B 95 51 1F 4E C3 5C E1 89 D0
 5D 50 E1 C2 35 58 C2 B7 B3 6C 43 CD CF 9C 7F E5
 2C 53 79 E4 9A 72 F1 36 58 22 9E E0 AE 37 98 8C
 B1 FA F1 58 E4 D9 E5 AA 38 7F E2 DC 8A 6A 37 59
 00 FF A6 25 A4 19 C9 74 51 95 E2 06 05 AA BB F5
 50 92 DB B2 8C 41 2C 13 AA A4 AE 70 0A 76 C9 A2
 F5 D3 DF AC E8 DB 04 1F 4D 6D 18 7B 26 97 39 15
 62 C7 81 55 68 ED DF 22 1C 48 A7 0A E8 CF 16 84
 9C 26 3A 4F 70 74 D4 8C 64 A8 09 0C 4A 90 0F EE
 A4 A6 E4 62 9A E8 4A 58 B8 6F F7 1D 27 0C D4 50
 F1 60 3B EE 4B 3A 6F 80 ED 1F 8C 5A F0 9A 52 2A
 60 60 80 B1 63 BC 07 B7 EE DD CC 44 E0 0B 14 D2
 76 AE 1A 82 75 01 E6 74 B1 43 10 34 D4 61 B5 0C
 8F 34 78 76 6B AD 85 F7 43 D9 C7 59 E0 7C DE 91
 CC B5 5F B8 A7 14 F4 70 6C AD 03 C3 F8 55 66 9E
 90 35 DC 86 CC 95 AD FF 6B 39 32 DF 80 14 B6 DD
 11 E0 38 8A D3 61 0F 09 2F DD 2B BA EF 75 3D 25
 46 9B 6A AB D2 E1 12 AC 9B 83 08 9E F8 16 E3 CC
 AC E8 BB DA 94 3C 92 97 0D 4D 8B 1C 50 35 09 C4
 A3 30 25 0E C4 5D 69 B3 5C CD D7 8E 3C 37 EF A0
 1B 0B 90 DA FB 00 17 FD 4F 56 D2 7D 2E 75 94 18
 D2 D5 C7 59 2E 0E 5B 85 5C 87 87 98 4A 34 42 A9
 12 B4 75 6D 9E 3C 0D BD 0B FE E7 28 67 48 68 8B
 F6 A6 D2 6B 86 B6 4E 4B 57 30 26 6B D8 73 84 D5
 AC A4 8C F4 2B 5F BE D9 8C 72 68 7E E4 FB 8E 58
 13 E0 13 10 C5 1F 08 23 19 D8 85 B0 7E 9A A0 41
 86 E5 B2 06 C1 BE FC 19 34 96 CF 16 4D D5 7A F5
 95 59 AD 5C 6B 42 35 63 D3 45 FC 57 76 20 C1 71
 1B A7 B8 2C 21 69 7C 24 B0 99 03 7A 1E 82 0A E1
 EC C3 F2 3A 68 C9 67 A4 3E 92 11 1B E1 58 2D C7
 25 AF D0 79 A2 D0 50 2D 7F 75 DD D3 1E 6D DE E8
 EB BB 27 FC 18 EC 45 4A E1 FE A1 21 DA 44 F6 7D
 76 EF 6B AB 90 3E DE A0 B8 67 B0 F4 1C 35 33 70
 D3 2B 8B 91 B3 94 63 68 60 B9 D8 CD 01 32 48 05
 45 F9 62 5A B0 AD DA E3 D5 0F 45 E8 3A B0 EB D6
 5C 04 0E D6 0C 36 24 EB 33 BB D9 4B 8E AA A8 63
 E1 4C 07 39 8C 0F E8 8F 12 9D 1D D9 B5 9B 85 2B
 DE A8 34 E7 54 65 48 CB C2 75 0E 55 C7 07 52 0F
 81 62 51 B1 73 76 F9 3F 9C 90 CA 41 22 6E CC 54
 54 6F 48 90 0B 7D DB 48 69 F3 F7 8C 55 EF EA 77
 0F 08 38 B2 CB 3F 57 17 54 2E 2B 0A 7C 0C 30 71
 B4 A0 BF 59 A3 0A 50 C6 15 99 A0 C8 57 43 2A 9C
 33 FC 47 34 D2 43 FB 74 D1 F2 51 4F 46 13 F4 C9
 C4 0B A0 0B 51 7C 47 8B 7C F9 A5 32 60 6B 20 1E
 CD 8F 02 8F 97 9B E6 10 FC A1 65 64 8E F9 94 0F
 7B 46 25 88 89 70 13 6B 1D 54 BC DA 6D CE B8 39
 08 E3 83 1E B6 72 E5 C7 03 51 D6 8F 8B E2 27 27
 30 70 21 DF B6 A4 0A 0C 25 84 7F FB A4 5B 43 52
 BB 9B B5 FC 20 AB 23 33 9B CD 14 D2 C8 A2 91 A5
 FB ED C0 71 4C 98 AD 70 9D 55 58 7D DB 1C A4 13
 EA 27 8B 37 18 B5 FE 7B DF EF BB 38 8B B6 AF B5
 CB E4 BB E6 08 D6 69 67 9A 36 A7 1C 23 7D A7 E7
 A9 12 24 08 12 EA EC D7 77 1C AA 66 27 D3 29 B3
 C4 DF D0 E7 6F CF 05 CA F4 22 6E C1 6B 7F AA AE
 8D 16 5D 27 21 E2 8F E4 FA 70 A4 69 0A 0C DD 35
 2B 22 F1 09 0D 4A 73 0F C0 E7 CA 61 89 B7 84 F4
 B9 44 14 92 C2 7E 8C B6 DB 5E 43 C2 40 4F F6 C9
 01 FE 6F 94 AF 3D C2 BE 62 E8 E0 61 B6 AB 79 61
 FC 7C 88 7F C0 50 C0 18 6E F9 F2 5E 12 CC E4 94
 6D D1 78 EB A0 5E 8E FF 8A A7 61 D5 1C 99 BA 58
 64 4C 98 D4 82 A0 40 EB 7B 64 6F 83 4B 1C 76 2B
 5E C4 74 C9 F6 51 50 76 41 3D 82 FC 03 33 15 0D
 07 D9 6B 2D 0C DF 3B 48 DC F0 D8 33 0D D7 E7 8E
 A3 2E 29 98 03 02 54 D9 6F 76 6F B0 7B 5D 50 C8
 75 6D 26 69 5F F6 18 65 5E 0E 33 45 C0 1D DD 31
 D0 C9 66 47 6A A4 4F CA 75 13 71 AD 87 26 6A 33
 6C 4C 06 08 57 D3 3C 98 6C D1 4E FC 70 25 71 22
 8C BE E5 0A F0 BC 3C 77 4D 26 15 52 70 4B 56 BC
 CB 43 15 B1 45 9B BD 4C 9E 29 E6 1B 5B C0 39 4A
 49 87 9E F1 A8 1E B4 56 6E D3 50 E1 22 67 8D 32
 C3 58 88 AA 19 27 D5 E1 82 A4 C4 77 94 33 B6 D8
 8D 35 55 EC 73 DE 77 DF 27 46 3B 6C 99 B8 93 FF
 63 CB 34 7B FF 19 FF 9C 57 FB 65 F6 BC E0 10 E0
 F2 60 39 1B 10 C6 B7 D1 B0 70 AE 40 79 9B 5C B5
 05 D6 45 12 03 87 F4 0A 2F 0F DF 03 36 13 CC 6D
 2A 58 D3 72 BB E4 7A F3 AD D4 A7 D9 C7 9E FC AE
 7D E6 4E E6 9B 13 4F F2 5B B7 79 60 56 73 C2 62
 BD 6B 56 B0 74 3B FB 99 7A F9 0B 89 34 DE 9A FB
 3F E3 EC AF 9C 2B 4E 0E EC A8 A4 F7 D5 05 C2 D8
 5E 2A 91 5A 36 25 35 4E 54 84 F5 60 B8 91 E3 DB
 99 47 F9 3F 72 27 C8 21 01 D1 91 BF 94 77 7A 4D
 AB DC 6A 60 94 E9 B2 6A C1 E5 BB 6C 81 BC B9 EB
 5F C3 B6 65 94 56 16 10 DA AD 67 D2 96 45 32 DD
 50 82 5E 82 E8 84 71 A1 3D 18 BD F0 85 36 36 82
 97 A2 5D 24 0E 6D D3 54 AD 68 F7 51 E4 1A C4 93
 B3 5F 38 A5 CD 4E 08 54 3A AB 34 1D 07 4B DC F6
 97 5E 9A F2 A1 3C EF 87 43 E0 63 2F 12 66 FA 35
 FB 47 C6 D8 EF 38 F4 0A 7A 88 69 04 DC 64 AD 42
 4F DB 5C 58 54 F1 B3 1D 7C 5F DC 8D 18 FA 2F 89
 AA 84 C1 C9 84 85 90 51 A7 FA 71 25 BB FE 06 73
 02 F7 10 BB 6D 6F DD D9 2F CE 29 72 0B 95 D1 FA
 1C B2 5A 17 0B 80 37 D5 11 E4 E3 05 74 CD E2 06
 7C F3 C9 3A 58 E8 BA D0 94 A8 6E 15 3C A0 E3 13
 3C 56 73 60 E4 39 7B 3C AD 69 DA B2 12 ED DD C8
 B6 81 C4 50 67 4D ED 3E 58 27 CC EF 25 7D F5 E5
 EA F7 CD AB 72 2F 1F 8F 48 D3 69 68 4B 1C 43 D9
 16 B8 00 DC C9 9B 5B 0A 55 58 DE 49 C0 53 7F 21
 78 18 EC 74 AC 52 2C C7 41 20 CD 4F 25 D4 A3 7F
 DE CF 70 EA B1 1D E7 D4 31 11 51 BB 37 C8 23 96
 A4 72 5F 6E 2D 45 74 1F 87 6B 35 EF 45 49 17 E8
 C2 16 4A E9 E3 5E 2A 22 6A 7F 66 0F B2 E6 A4 BA
 C9 21 1C 7F E3 4B 83 A0 0A E5 BF DC 51 25 52 12
 9A B4 E7 77 DE ED E4 A2 32 02 16 60 F5 15 0C 0C
 B6 8F 79 1F 52 4A 8E D0 A9 A2 6B 9F 24 7E 1D E2
 F4 D6 83 85 7D D7 95 DE F0 65 77 11 60 33 2D AC
 F6 D3 3E 58 4D 85 95 C2 A0 06 DF 31 59 AC 10 A2
 92 6E 9C A8 5E BF EE DB 7E D1 29 80 48 2B 77 F1
 51 2F 32 E4 47 58 03 F2 5E 49 86 8D 85 17 C3 D1
 AA 73 66 98 9A 42 D7 39 3E 45 5F 3C 1F 1C 21 85
 20 B3 43 C8 3F 28 55 7C 2D B3 A4 58 37 43 A6 FE
 EA F6 47 1C D0 2E 58 5C 14 C6 CD 98 BF 26 7E 63
 9E A6 D6 46 3C 97 E0 1C 81 12 C5 81 E0 58 2E B4
 BC 59 67 00 3D 6C 84 F3 57 D7 62 B9 AB 94 65 25
 C7 88 3F A4 11 61 BD 45 6A 2F 36 34 61 65 4C 1B
 3D 15 36 08 98 7B E7 E5 13 89 4D 70 0F 39 4C A2
 71 28 BC 46 A3 BA D1 41 2E 5D 14 F6 E4 8D 5C D1
 B0 A6 BF 1F 75 EB F1 B7 49 4B 43 50 4D 4E FB 26
 9C 51 27 74 E8 CB 89 B3 97 FD D3 9C E5 A7 B9 F0
 10 23 01 6A 9E B7 8C 74 C2 9A EB DD 09 9C 21 E1
 76 AB EE 1E 8D 84 99 9A C4 58 97 5B CC 84 6D 67
 11 AF 56 63 6B 64 53 A9 0D B9 87 64 91 40 9C 85
 AB D1 10 57 A3 64 BD A6 A6 F0 45 3D D2 31 47 7F
 13 81 C3 C6 C3 C4 C7 DF DD 67 49 D1 6A FE 96 F3
 59 87 A5 96 27 AE AC 7F 39 C3 A2 67 36 1E 56 86
 AB 2F 12 10 42 8E 61 6F 5C 53 05 E1 C9 5B B7 B7
 18 F2 61 15 3E 53 A2 6A 7B AC 82 D8 49 C2 14 AB
 E8 DB FD 42 53 95 06 3B 73 08 60 9F AD D1 8A C2
 B3 C6 F2 64 09 7C 05 6A CF B1 A7 CE B8 F0 AB 74
 E2 81 14 AE F1 1C 5C EA 5A 80 0E A2 3A 39 AD 2E
 46 9D 36 C3 EF 7B 10 EF FC E9 65 43 AC D5 FE 8C
 66 6E CA 13 90 DE 9B 22 21 DA 96 0F 64 28 D6 39
 37 1D A2 EA AF 79 FB 90 96 74 0D B3 C1 FC 7B 0A
 B2 A8 F2 6F 93 98 2B 13 F0 DC E8 78 CB 2C D9 3B
 08 B5 B5 62 20 E5 AF 79 B2 B8 FD 40 66 0A 45 B6
 6A F6 3F 27 A6 CA 92 36 B1 9F ED 28 E3 33 A5 C9
 77 C4 C8 14 CB 2F DE 8D 87 FD 3E 8E 5B 36 79 5A
 2A 82 F2 AD 80 9D F8 47 8D 15 90 9A 40 6B 18 B8
 7B 20 A6 79 D2 52 B3 E9 9B 7B A7 3E 48 52 A5 0C
 82 09 10 0B 13 1C A2 AC 3F 04 7E E6 9D 14 BC A5
 0A 0C 36 AA 82 34 A1 58 43 C0 21 9C C8 E2 B6 43
 85 FB 88 A8 3B 26 BE D0 80 57 D6 CC 86 49 A8 DB
 32 2E A7 74 6B E3 D3 04 B1 F7 77 F2 27 F6 CE BE
 DB E8 D3 FA FC FB E3 23 99 3C 1E 75 57 DB 0A 09
 F0 2F CE 9D BE 91 0A 0B 48 5A 6B AF 3C E1 F1 7B
 7F 65 AF BC 16 B5 53 38 A3 9C 72 26 49 BC C8 6A
 67 1B 89 EC DD 2C 79 FE C8 1F EB 35 83 71 93 B7
 6D 35 F3 FB 52 F8 50 95 35 E1 B0 97 D5 1C 63 FE
 46 CF BE 0A 2D 8D FB 6A D9 A9 16 7E B1 F1 26 05
 6A F2 A5 D9 AB D4 0F 08 14 62 74 F2 17 9F 6B 4E
 2D 9C AC 04 16 4C 80 F3 98 D2 76 B0 E0 8B A8 F8
 FC 25 AA 64 B6 C2 8B 78 2A E0 80 4C 4B E3 E0 7A
 AC 49 11 59 D3 77 BF 60 5D 62 4B 3F D5 79 3B A7
 E2 9F 26 CC 71 48 28 93 6D D8 7F E0 90 A8 66 83
 E9 3C 46 36 7D 75 EE 5B BD 0A 81 61 2A 0D 2D 58
 0C 4A BD 50 BC 31 D9 C2 0F B2 AD F1 24 01 48 5A
 2D 3D 02 C4 71 E2 9E 73 4B 3E E7 E7 9E 1D 76 AA
 42 89 A7 50 25 9C BE B0 42 69 80 7C 0D 33 7C C1
 77 E8 DA D9 31 7F C2 88 32 17 0F 1F B5 F3 5B 34
 6F C8 9B 1A 82 A9 53 2B 72 76 35 7F 3C 34 57 45
 7B 00 D4 8F 45 8C A1 7D 6B 68 9C A6 70 B3 4C 4F
 24 32 68 1E 60 53 7E B3 8E 4C 84 CA 85 40 9A 07
 3E 10 BA C6 84 D8 FA EF 5B D5 6D D7 29 73 4B DC
 FB 95 00 BE 44 A1 12 86 93 AB 28 9C 4D 6A 9E C1
 79 35 73 E3 D8 22 A7 A0 92 99 D3 74 30 31 1F 9B
 88 2E B3 12 27 B4 B4 26 58 23 A0 43 22 89 75 85
 A2 3D 92 25 6F 22 E5 A5 CF 90 FA 75 97 8A 4F EE
 A8 D2 53 41 6F BD 4C C4 7E 24 49 B3 60 98 E2 30
 EA DA 2F F2 D9 DD 48 0C 44 23 D1 FD 88 88 D3 33
 DA FF ED 39 FF 92 BC FB 1A 46 1F 74 8B 9A D4 2E
 B6 70 AE FB 99 CE 30 10 DC 17 B9 32 F7 0E D6 3C
 6A 0B E4 FA E6 39 33 D1 14 B4 90 36 83 9E C4 23
 FD 6D 24 3D 70 01 B6 19 49 25 C4 63 72 AC 07 12
 CE 23 B7 91 18 15 AA A0 3D 23 20 08 0B B2 5A 06
 AD 2F 99 88 5C 7D 36 22 5C 67 18 62 03 02 4F FD
 30 67 12 63 CC 26 4D D4 5E E7 D5 52 72 5C 76 D5
 F1 42 0D 16 50 B6 E7 C8 5E F6 96 A7 95 1D 6A B3
 18 45 66 8D 09 D1 DF 97 58 DA 04 35 82 79 4E EA
 F0 E8 AF DE D9 66 D3 EB 61 D7 2B 05 CB 9B 08 CE
 73 53 A9 45 C1 CB BA D4 B6 83 B4 A3 4C 29 27 A3
 95 06 58 B8 5B 53 AF E1 70 63 60 30 19 ED 4E 97
 92 47 AF 18 0F AA 7A B4 BE B9 C0 6A 37 50 5F F5
 CF 45 3D 41 2A 7E 76 F2 92 15 9E 93 45 1B 81 C6
 51 6E 6A 24 E9 43 20 C2 99 64 19 94 8D 6F 9C 93
 24 45 30 B0 1A 0C 33 7A 02 8A 9F 87 40 9E 52 C7
 14 72 27 9F AA 12 5A 3A 38 88 DF F9 7B 4F EA 43
 60 1E CA BE 75 3C FC 75 92 A5 42 6F A8 AE CF BF
 B5 8D C6 9D DF 0B 91 CF 48 88 80 3D 01 1C 29 D6
 24 04 E9 BE 77 CF 65 39 9F 5D E6 3E 43 88 7C CE
 CA 54 FF 5B 58 64 C3 77 1F 41 82 80 0C D7 88 82
 07 94 A9 91 ED D6 51 8D 38 B5 BA 2E 2E A8 E2 99
 70 02 03 75 AF 27 E1 AC EF 79 7D 32 47 11 4C 23
 F3 47 89 64 FF 29 2E 8A CC 66 07 6C 27 05 55 95
 9F 97 0A DF 29 5C 73 68 FD 06 4E BD F4 BF 40 C6
 74 35 FD 5F 90 A2 97 1D D2 EC 98 77 05 CD E2 C1
 9F C5 17 88 05 2F DD 1A A5 E2 D7 D6 28 A7 88 93
 42 70 FF 70 01 A8 7A 51 17 37 BC 18 E6 AF 80 84
 43 EF 07 FB 2C 7E E6 E1 E1 D7 F2 13 13 46 75 0F
 D0 3F 16 86 2B 88 B9 91 55 B3 82 77 CA D0 9A 82
 AA 99 90 63 3C 2F BB B4 4F 6A 24 50 33 44 8D 00
 6D 17 1B E1 29 36 B1 63 D0 9F 48 80 50 77 68 82
 D3 7E 51 4C 7E 78 86 A2 5B 77 4F 85 11 92 21 A6
 F6 91 39 CC 54 2C 43 D8 DE B0 A5 88 08 21 88 F0
 20 21 9C 81 3E 86 04 A3 BC 34 06 89 92 24 A2 2E
 B0 3A E5 1C 7D C6 88 24 D4 F2 27 26 58 90 1C DC
 DE 1F 4C E8 B4 96 9C 1D 71 31 99 E4 44 40 1A 24
 27 23 65 40 A2 C4 8A 6F B1 4E C1 DE BE 90 4A EF
 CD DE 67 47 F3 43 6D 76 74 39 5B 66 D6 7A 23 9F
 6D DC C7 38 A0 3C D1 A5 0A 4F B1 F1 2D 0F 7A 29
 F1 48 58 6B 38 38 26 9D 9B 53 E7 CB E1 67 C1 4A
 E4 B9 9A 90 3B 58 EC 4D A9 50 28 24 90 53 A8 88
 94 D8 F8 37 4B A5 46 17 69 24 95 5C 5F 68 E9 32
 1D C1 C0 67 95 E5 06 76 F7 8F 2F 43 EA 8C 76 15
 3B 34 8F BC 46 64 B4 9F 1D 13 DF 40 E8 EF 9C FE
 E4 2E D1 BB 94 49 45 51 7A BC C3 47 F6 14 5F 04
 81 E4 B4 F8 55 39 E5 BE EE 5F F8 58 09 46 D1 90
 79 07 AF D0 15 B6 58 E0 7C 7D 29 6D D7 F0 47 B0
 C2 30 D5 E5 50 13 B1 23 4C 89 D0 F4 1C F5 9A 01
 B3 4F A5 9D A1 0F CA 28 8D 78 BF EE E9 D1 28 42
 B0 48 DF BD 3C 2E 70 F9 20 56 75 3D 20 D2 BB 7D
 1C FD 8F 73 B8 BF E7 3F B7 F4 A7 DC D9 96 65 8A
 92 22 B5 51 D4 4B 94 74 55 95 5C 87 6E FD 9E 9F
 11 DD 38 2F D0 31 C8 68 1F C4 96 30 F2 B0 C7 61
 E7 54 F9 9A 76 EB 2A C9 B0 54 AE 52 B8 61 83 D1
 A7 EE 2B 1C 7C 57 89 EF 1E 66 B1 E1 FB C7 43 30
 FA CF 55 8E AE C7 2E F9 C7 28 CC 7C 9E F8 7D BA
 45 8F B5 64 90 AD B4 1B 02 54 29 88 8F 34 97 81
 87 4C 76 7B B9 73 9A F0 6C 87 65 97 CC D2 D4 F7
 EE 86 01 22 AF F5 B0 05 81 21 0E FD BE 30 77 BA
 D6 2D FC 83 6A 49 13 B8 00 89 A3 4C A3 7B 3A E3
 D0 9E F9 DD C3 94 E5 81 85 61 39 FF 96 0E D5 4A
 D3 C5 D6 D5 FD 35 41 25 A0 87 C9 0D 54 55 E8 06
 44 6C 71 4E CA 83 14 43 73 7B C3 BD E6 FB 95 3A
 36 F1 73 BD DD 67 B3 25 52 2C DB F8 D0 DD 40 DF
 39 72 C4 7E E1 96 CC 23 15 37 13 85 A8 09 2D 65
 A4 85 8E 54 8B 6E 9F 58 63 66 ED 44 A5 43 6C 9E
 AA 83 C7 E4 58 FD 44 0D 88 FA 04 08 B5 EE F4 5F
 DB D4 3B A0 F7 3D C1 07 07 ED 7A F9 9A E1 D0 CB
 F3 2D 82 45 9A 3C A5 E1 66 14 2E 55 F7 17 59 9B
 09 53 CB 6C AC E9 45 13 5A 26 BB 2B 40 9E DE 26
 93 EA 4E 77 62 C6 32 59 4F AD 38 84 9E C8 97 88
 D2 1A 3D A8 C9 8C FC 8F 93 3B 2D 7D 1D 0B A9 33
 B3 EF 08 7D 39 89 0F 48 A5 18 FE EF D9 0B AD F9
 2C E3 89 0C 4E 9E 10 66 3B 36 33 A4 D6 E2 E9 EB
 86 31 59 53 C6 CA 72 B2 04 37 95 AD BE 59 D1 37
 E6 58 D0 BC 0F 1F 5B 65 7F DC 9B 86 FB B2 D8 8D
 01 60 1C FF C6 35 BE 07 2F 5A 41 FC 53 CC 12 50
 F7 F7 78 27 7C 67 62 79 9A 8E 6B B8 E3 79 87 54
 1A FE 62 E9 BB 40 C4 53 92 C2 61 EB 6C F5 DC 76
 50 54 3E CF 50 2A 9F 3F F2 67 58 77 68 3B DD 76
 F9 63 36 52 9C 95 FF FF E3 5C 44 82 B6 D2 85 AE
 81 3F 66 39 FA 23 26 97 C2 BD 3D 46 53 6D 8A B8
 65 2B 26 AD DD A3 9F 55 33 D3 3F 74 16 11 07 DD
 3E 55 54 D1 E9 CF F1 FD 3B 52 1E 0C 49 30 BB A9
 35 F9 47 FE A5 3B 11 B7 95 C2 77 9A 04 C0 9E A3
 89 FD 17 30 35 71 7E 5F 29 09 11 02 98 55 9A 7D
 D0 88 4F 41 EA 51 57 90 BD 09 65 83 21 E5 17 05
 42 09 BF D0 FF C9 DA 6B 2F F2 7A 26 48 E8 6D 03
 54 2F D6 24 60 DC 1D 16 E8 1B 70 23 76 95 CC 6D
 2B 7D 08 6E 7A FC 97 89 A5 72 75 31 4C 5B 07 03
 41 83 5E FC F5 4C AF C9 18 BC 25 C5 09 95 99 18
 62 D9 DF 6F 89 86 F7 9B BD 93 7B E3 80 61 FF B2
 BA 38 EB E1 C3 42 94 E9 65 C0 75 84 7A AE BD E0
 7E 28 22 58 43 44 16 03 AF 48 E1 C3 7C 9F FD 32
 F1 99 E0 0A 37 A8 EA 0E F8 DA 3A 22 DA 72 14 3D
 E7 F5 F1 A4 3E 84 2D 7A A3 01 C4 F8 45 F6 FA AF
 2D 33 B8 01 8A 16 DB 39 E8 BF 22 0F 30 BA 2B 9D
 50 A1 33 35 F3 23 87 2F 56 02 79 A2 8F 4F 74 2A
 6D 81 31 DC 27 46 24 BB D9 A1 B2 91 DC 49 A1 0A
 06 F5 D0 A2 2C 39 83 BE 68 8C F6 02 EA 09 65 6E
 53 A7 23 D6 4B BD 00 FA 33 0B D2 F9 8F 77 32 80
 83 A8 0A 76 6C A1 AC E8 A0 81 6A AB DA DD 49 86
 F2 24 93 14 D3 B7 1D F0 0C 5E CB 8A B6 F1 96 0E
 06 1F DE 58 5D C5 88 6D A6 E3 86 19 CC A4 1B 10
 3C 1A 31 12 A1 28 23 F2 FC 9F 6F B6 A4 48 0C 05
 A7 BF 02 B8 49 44 9F 6A CE 9A 99 23 2A 74 C1 E4
 2E AF 79 45 23 16 E1 5A 3E 35 1F 41 E2 E6 3D 9D
 48 1E BB 05 28 17 FF 44 BA 05 A1 41 82 8D AD 42
 91 C6 3E B9 C1 FD 3E 65 C8 B4 91 D0 B7 CC 02 0E
 30 7A 46 86 9E 05 5D 63 EC 4E C9 E4 40 9D B6 D2
 C6 61 F4 35 FC 14 FB BB BB D8 2F C7 BE FD 76 84
 E3 98 49 15 96 BB 21 08 0A 44 21 CC E6 25 18 E8
 22 2E D7 19 1A E9 3F 0B 23 A9 1C 8A 1A 3E 36 BB
 3D B5 95 86 5B 48 C1 A2 C2 A9 E9 F8 51 DF E6 2F
 BE 1C 1B 25 14 9B 05 C5 26 3F F5 4B 32 9E 5B 9B
 6C 23 2E F9 EA 23 FC 91 1A 19 4F 28 0D 6C E2 2C
 14 70 BB 23 3B 86 D7 F9 9C 9F 0B 39 0A FB 04 D1
 1E EC 04 C3 A1 13 76 25 BB 57 75 D8 2E 8B 5C D5
 60 34 EE F1 43 32 F0 98 8F 9B A0 02 D7 C2 1A 67
 90 E6 AB C2 57 8B 56 F4 D8 C1 0D 52 5B 3D 05 FD
 21 A2 4F 5A 63 E1 C1 AA F0 73 F1 28 69 0B A1 B8
 FA 92 4C A5 92 83 1D 78 7A 76 8C 7A 43 FC 97 67
 CC AC D3 62 FB D0 1C 86 4D 4A 9C 6F 6D 40 DF 48
 5B 37 B6 33 F4 42 92 AD CA 26 C1 2B DE 6F 81 4E
 3E EC C3 0A 8E 4F 43 BE FE 7A B2 61 11 F8 54 09
 26 00 93 2D C0 A2 76 3B AF 2D 0B 2F 41 5B 93 C7
 89 12 F2 CF 32 46 81 E1 EF 47 48 9D 1F 1E 35 C1
 F1 6C 22 59 81 FA 72 E0 1E 64 BD 0F 77 E6 A4 EB
 9E 47 79 0E FE 5D 7B FB 51 A6 CE E2 9B E6 76 D8
 61 0E AB 73 98 BA 5E 6B C6 24 FD B7 2C 35 41 A9
 B5 03 52 B3 5E 77 CA 2B 40 EF 4A 7E 6A A7 C3 20
 C1 D5 60 49 DB 9B 19 69 A9 54 AE CE 13 F7 F2 38
 32 66 04 2B A5 A4 05 A6 8E B8 96 67 12 B0 64 43
 73 29 22 B7 C5 F7 A2 50 0C 9D E6 B5 03 FC A1 68
 8B 1F C4 A9 2E DE A3 6C 20 FA D3 95 5F 46 0F 60
 0F 1A E0 29 E7 09 00 FB 63 CE D0 61 76 89 35 CC
 E7 46 87 69 D4 6E 67 B3 7A 00 00 28 75 70 C4 CC
 BE 22 E8 D9 72 3A 46 CE FB 4A 72 C4 74 D1 1F 40
 5E 28 92 7D 06 09 D8 AA EE 94 E3 BF CC 61 12 13
 FB 2C E0 33 9A 56 29 43 25 30 BE E6 57 62 4B 04
 88 D3 FF 56 FC 3A 1D 25 08 24 98 85 FB 19 1E 7E
 C8 7E 8D 75 E2 9F 8E 8D 92 36 D3 5F F1 DE A8 63
 38 FC D8 98 2F A7 12 CF 01 66 66 A3 5E 0B 7D 7B
 83 2D AF CA 0A 3D 8D A6 DB C1 30 0E 3A 04 73 92
 84 C7 4F CA E5 CA 21 9B 86 B4 1C 27 13 B6 70 69
 4F 24 7A 0A 7A 1F DD 4A 4E C8 A9 84 6C 88 CF DF
 15 FB 3C B3 22 62 4A 6D 44 14 85 F5 D0 AD 4B F0
 09 CD E5 F7 F0 0C 3B DC 65 69 01 5F 15 5B 67 24
 DD CA C0 B8 54 E0 55 21 A7 9E 3B 7A 6F 47 91 30
 C5 EA 0C 97 5A B7 E2 2F 9E C1 73 40 98 76 CD 3C
 B8 6E F6 EC 40 91 53 0B 12 F6 1C 44 D7 A7 40 1F
 FD 54 89 9F 98 9E 4D 7A 1B C0 C0 EF 00 2B FB 64
 B0 0B 45 76 41 FD B6 BF A6 51 D2 A9 15 EC AA 92
 F3 A8 9B 2B 42 AC AD 80 45 22 69 AC 5D 0C 3D A2
 45 29 F9 77 61 01 33 09 CE A5 84 4B E6 49 28 76
 5D DB 73 38 0C B8 2F C6 4B AA D8 4A D6 1D E4 CA
 25 CE 4C 00 57 D6 42 A1 78 5C 8C 7D E2 94 DA 9B
 D5 7B AB D3 72 FF C1 32 5A EF 29 66 96 39 39 08
 A5 26 DF 7E 80 A5 99 4B 5C 6F 63 6C 4C 6B BE FA
 FE 37 75 0C 0D D6 88 7D 5D 76 99 DD 0A C5 54 64
 E9 24 17 C0 49 22 75 91 9B A0 17 85 28 75 91 32
 84 B3 6D 1F 37 39 81 2B 51 A1 68 8C CF F0 80 09
 98 B5 B9 80 D8 B6 68 4D 17 79 C6 75 09 7B 75 58
 27 AE 32 8F C4 D3 3B 26 38 D9 C8 A2 77 70 50 2A
 DF 41 15 3E FF 1F 4A 7F 37 DD F7 5F 95 3A 5E 87
 20 F6 B2 E1 CD D1 A7 F3 98 3A 97 AE 6C 30 FA 18
 0C FA BB CD 0C AE 13 74 C3 91 40 84 C2 9F B4 03
 66 57 05 08 96 5B 4D 3F 56 AE 12 7E CA 1E 2A 53
 06 D4 5D E9 4B 1A C6 30 51 B4 B1 18 CB B9 E6 DF
 82 55 FC 8B 8F 01 44 8F 42 FA D8 97 CC A2 77 3F
 F7 0C C9 05 E4 DD 7A 80 08 D8 B0 0A EA C0 C4 D8
 5E 2D FE 9C D9 46 AD 53 65 4E F9 58 1E 26 B0 4A
 D3 72 CF 2F 77 63 A5 8F 06 D9 0F DA 2E 82 36 8E
 64 86 62 3A 9D A4 80 F3 A4 2D EF 14 6C A4 9E F5
 41 B4 6A CC 56 8D C2 3D E2 91 5F 78 75 59 62 C8
 25 7B 79 19 A3 34 D5 0F CF AC B2 32 28 F9 EE C8
 8D 0E 5B 4E 9A B3 D9 D1 C3 AE 4D 7E ED F5 D8 A3
 A3 88 B4 80 69 A6 54 70 26 93 97 EF 38 03 67 34
 A3 6B BB 8B D1 D1 AF F2 09 9E C8 06 CD DD 43 D1
 C0 99 0C 07 5D 83 40 86 07 31 7B C2 FC 88 18 C4
 A4 78 68 71 7D 62 1B DD 04 D5 A4 E5 8E 4D 44 A6
 3E 97 0F 4C 71 02 3A 98 EF C1 7B 4E 2A C2 AD 69
 39 42 45 03 12 2E E2 F3 02 FE 65 2E A2 89 8A C7
 E9 A8 46 82 9E 93 EB 4C 5E AD D8 38 1E C4 0C 01
 6E 2C F6 B6 69 EF 1D FA E3 0B B4 4D 90 55 0C BC
 C0 1F 3D B2 54 DA 96 E1 BD FE 5F B9 10 EA E1 90
 5B 54 7B 66 61 52 2A 54 67 F8 DB 88 73 D9 E7 BF
 29 E9 F9 6D 36 69 70 A4 CC 62 5D FA 8B 34 F9 FC
 6E 30 96 8C 67 54 7C 54 FB 7F FD A6 7B 99 8A 18
 82 E0 FB 79 73 EF 21 7C 59 DB 5C 3E 2A 35 0E DC
 F7 7A 80 4C D8 75 D2 AB 93 F5 A6 29 D7 DA 77 94
 72 28 37 42 05 5A 77 6A 77 64 60 E3 C0 0E 24 94
 D9 6D 4C 31 97 90 63 1D B2 91 45 AF 25 3D AC 2F
 04 75 47 BD DE BA 6B 3E 6C E7 6D 3F 6D C0 4C 3B
 3D 86 A2 CF 6C 74 C3 C9 1F 8E C6 2B 45 A3 C9 F0
 1A E4 AF 08 1F D4 06 92 BC 1A B3 B5 C4 73 18 C9
 F4 B3 70 C5 06 C6 07 0B EF 4A 8A 43 E4 C5 53 AA
 01 BF CE 9F F9 0E FE 90 E5 4F B3 AB BF C9 AB EE
 E5 F0 94 60 DA EC C0 E5 54 2E EF 89 E5 EF 36 DB
 0F 79 BF 3D F7 0D 37 1E 5A 36 82 16 35 18 3C 6E
 C8 F1 0E 02 95 C4 9B C1 9F 13 EC 40 D9 67 6B A6
 C1 6D FA 38 00 63 F5 46 79 A1 79 A9 B1 14 45 EF
 B3 55 17 28 4E 2F 41 4C 25 B3 D9 34 65 D8 66 29
 67 9F D9 ED FE EF 17 E3 78 F5 D9 8A 56 0E 59 4F
 38 83 1C 4D 35 09 08 1B AC 71 4E 91 45 D7 C9 87
 48 76 C7 64 93 06 88 78 B1 12 6D D3 4B 59 82 C9
 26 0E 73 D4 30 C7 A0 99 9E 3D CA D1 AF CF BB C1
 05 92 E7 15 87 C7 EC 0F 3F 1B 5C C0 B3 17 D0 CF
 D4 D1 8B 0B 9B A9 AF D6 99 F5 A2 90 64 BF BA 75
 30 40 22 9C D0 2B 7C 10 DA AC B9 79 8A 2B CD 61
 84 6E 59 A0 46 7C AD 39 0A 5C 23 96 F7 86 9B AB
 42 D4 A2 C1 7F CC 9E F8 4A 01 48 F4 9B 0A 5F A9
 DA 53 FD CF 4A 4A 08 C8 23 6C 42 0E BD 6C 32 BB
 52 1F 61 FB 8B 34 E4 EA 4D BD A7 8D 04 F8 F6 65
 41 1E 74 CE 51 C5 67 5D B7 1A FA 3D 6E 51 66 F7
 1B A5 31 B0 6E 19 1E 0C 92 4B EC 06 11 BD 20 2C
 56 0B F4 76 6E 57 B1 CF 35 B0 F8 29 20 74 87 4B
 15 B5 64 90 ED C2 B9 13 3D 7E F7 C9 51 22 96 B4
 EB 3C 80 D0 BD 29 A9 E6 4D B2 7D DA E8 F9 5B 97
 F8 26 89 20 17 EF DC 16 4B CD E1 8C 92 E2 1D EC
 40 42 C0 6F 4A 5B 60 09 39 23 2B BA 9B 9D CD 44
 78 57 E3 C6 B4 F9 6A 46 AC D2 0A 43 FE 57 7C 47
 25 15 E2 26 FF 17 93 05 2B F9 40 F5 05 07 D2 FB
 9B 75 CC 0D E8 E6 45 7E 91 3A 2F CD B7 AE C5 7D
 C4 B7 E2 93 3E D8 B6 32 0C E0 D1 3A A0 96 3E E2
 E8 BC 4B DC AC FC DB 8B 28 2B 8E FB 66 14 7C E2
 3D 29 0F 69 9F C2 28 31 41 68 42 50 38 46 9E AD
 92 59 C3 E1 26 92 B5 90 8C 54 00 78 28 79 C0 B4
 09 8D 4C BA D0 4F E6 B4 19 C4 C8 21 3A 81 27 E0
 42 D7 95 DB CD F7 45 F6 1C 57 21 03 64 6D 2E 7D
 21 3B F1 E0 61 2E 8A 18 E4 11 78 B8 FA E5 52 32
 C8 BE 96 BA B4 EF 21 A9 14 43 54 EA 2D 8A 73 95
 C8 75 06 8B 04 51 DB F6 10 20 0F 0A 77 B9 A1 60
 92 7E C3 6F 9B 96 78 8A 49 BF 91 31 11 5E 03 04
 01 DC 90 BD 5A 50 1B 3D 9C 09 34 4E 84 86 F2 BF
 94 63 8B 45 C3 E8 2C 51 76 11 AA 73 AA BC 40 F6
 35 4E 53 B0 4C 1F 24 86 52 C0 CB E8 9C D9 15 B0
 4A 3B 56 F8 35 53 89 9E 89 21 BB 1A C6 F2 D9 05
 E2 F2 F8 6F 11 EF 10 5D B1 6C 6E 45 18 80 39 41
 24 0D 26 3D B2 30 CA 1D 3F C8 17 F7 DD 87 55 69
 F5 C3 C0 DE 30 BD C2 CD EE F9 D4 F3 DE 9A D6 0C
 F5 09 B8 29 A0 19 E7 4A 75 EF 66 D9 85 64 E2 6D
 AE 80 F2 E2 3B DD E3 30 26 CD 00 DF 7A 33 22 7A
 83 49 21 83 8F DA 39 F2 94 DF 9F AE 2B 9F DD 4C
 55 5A 0B CF E9 0E 99 F6 0E F2 99 9A 3D 74 70 56
 89 E5 9B 67 4C 3B 8C 89 6F A1 95 77 5B 34 D9 A8
 62 28 09 91 9B 3D 67 0F E6 F9 2D 10 5E 3F F3 99
 34 BE 26 C8 DD 10 7B 20 3A B6 F4 10 99 74 08 7E
 5B 2B D7 2B 24 E2 14 CC 19 DC 7C FF 18 C5 97 2E
 E5 A2 3F AC B0 71 33 D1 BE 23 C3 23 58 55 87 32
 90 59 FB BD 23 12 AF 33 0B 02 53 86 6F F8 27 B0
 33 78 0C 8C 11 4A C3 90 D8 EC F1 C5 78 E5 EC 53
 2B 7D D7 DF E4 7B B2 DF 6D 7A 4A 66 C0 D3 4F 47
 E0 53 C0 7F FD 8D 2D F5 3E 30 90 DA CD C4 F5 68
 FF 1B 6A 20 BB 5D 59 F3 8D 91 FC 6F 4E 31 41 97
 2A 79 B5 C3 50 8B 1F BE 08 68 73 1C F2 77 81 04
 B0 32 0E 93 A6 2D 18 D1 EE 65 E5 CE 9D 80 A4 B4
 1B 6C 3A 00 2D 95 54 46 FE D3 71 2A 38 28 06 88
 BE 42 00 91 D6 46 27 56 08 29 79 6D 64 B4 34 92
 D6 BC 7D 27 1B A8 DA 73 A6 79 98 DA EA AA 8B 74
 EF 0B F9 0B DF 18 DE 70 5E 52 1D 3A 0D BC F0 D1
 1D B8 1D 39 84 23 23 66 86 B3 85 93 96 96 71 81
 E1 F4 37 E5 7D 87 A9 BB 2A 31 19 E5 CE C3 C2 05
 DD F7 48 D1 78 B3 37 94 66 3C EF F2 2F CA 40 C7
 94 42 A2 1B C9 A0 B0 51 4B C7 28 C4 B7 A9 02 B1
 AE 91 4D 1D C9 80 55 38 AA 2B 3A 22 9E C2 D4 7D
 12 24 D6 DA 5D 0E 5E 8C 3B D9 AA DE 98 83 AA 46
 BD 91 B3 86 11 F3 92 7D 53 37 2D 5B FC 20 94 2A
 37 53 1F CE FD 1B F3 34 E1 A5 26 A9 63 7F A4 2E
 5C D6 36 93 6D 54 AD 73 E5 15 A2 B9 5F 92 FE 7A
 E4 9A 82 BA 90 80 E8 66 B3 1E 0D E1 6A DF D4 61
 B5 39 F3 08 91 30 46 E4 DE CE 4D 34 52 51 2D E8
 53 5C B7 4F 93 7D 7C 9C 09 AB 3E 71 F9 AB E7 A7
 5C 74 46 4D B9 ED 25 81 78 DB 4D EC 65 35 35 9B
 31 16 58 73 73 BC 9A 55 6B 18 5A 34 AD C6 BE 2D
 1C E0 33 30 D9 C1 9A 96 6A 3D 8A E2 AB D8 AC 0C
 48 10 28 82 8C C5 D4 A3 FC FD 1D 12 BB 3E 39 AA
 5E 96 ED 5A C5 99 0A D3 00 AB B1 F4 65 27 6A 08
 12 33 6D 2C C9 6F 66 B6 F4 F9 7A 90 14 40 B4 71
 C6 B7 CE 57 FB 8C EF D5 45 27 C8 FD B6 CC 1A 76
 3C E3 2C F4 5C B4 4A 67 33 CD C6 C8 4E BC 92 E7
 45 6F 91 2D 95 6D 8D ED E5 4A 90 58 EB 76 A7 9B
 44 49 B1 D1 FC 25 97 2C 94 C4 ED EF BD B4 4D E3
 B1 FA B3 99 2B BC 83 6B 4D 97 09 9C 4E 99 D6 83
 69 13 A8 F1 D0 DA A3 FD 10 5F 90 0D 3E 1B E0 9D
 71 C8 51 4B 99 BE 3F 67 58 B8 82 9B DA 05 E8 F5
 35 1D 64 62 C3 69 11 76 AA B4 77 2B B6 5C 9E 37
 8D D2 2F 5C 3B 1D F7 14 09 87 E8 58 F0 D1 A5 19
 61 35 0E 70 2B CA C3 20 FD 14 88 7A 1E D0 BB 18
 EE B2 EE A8 29 8C C1 A9 32 DF EC DE 84 FC 46 5B
 E1 FA 5B 02 A2 A0 CF D5 09 98 1F 09 84 24 BC AC
 27 59 AD 65 04 81 41 45 25 69 BC CE 47 5D 11 D9
 DB 6C 18 46 D3 4D C4 89 22 59 96 2F 3C 5E 81 7D
 75 64 99 5A 9B 4A E8 DA 8D 54 02 DD 64 7D D7 B2
 E9 5F D7 93 FE 77 B5 93 7D 18 82 93 79 8E 6E D8
 B8 82 C0 33 4D AC 16 E5 FA D2 48 4A 22 AA 7A EF
 C1 AA 37 D1 A2 91 76 22 69 F9 22 51 E3 71 90 95
 7A AA D0 9E AD 5C 18 A7 85 ED 25 B5 9B 8F 9A F1
 00 A1 34 90 72 DB C9 27 F5 BA AD 1D CC CA A1 15
 6E 7D 01 E4 E1 3D C3 82 D7 02 7F 5B 50 44 42 4C
 6F 8A 05 3A 48 F1 D7 66 2B 68 0D 88 F9 95 DF 23
 DE CE 1F 88 2B 00 37 54 6F A1 02 C1 C0 BD 09 1C
 48 0A 9D 3A 76 72 13 5E 7A 5A C4 ED 8F BF D8 62
 A2 99 82 97 A6 8A C6 A1 64 68 A5 36 98 41 7E 7D
 98 E2 56 4A C3 A9 71 66 64 1A 5B 4A 2B F8 EE A3
 05 63 E8 09 6C 8B 8C 60 DC 9C 9B AA 02 8C 4C 8D
 7D 95 B2 E5 E7 D3 C1 A9 75 30 13 09 CF 64 5E 93
 4A F7 6D 6C C4 21 AF C4 B2 86 45 D9 AD 4A 16 B4
 B1 05 AF 59 74 11 07 6B C5 9D BA DD E2 27 06 30
 21 14 97 BE 8E B9 CC 96 12 46 25 8B 90 DB 21 B5
 89 CD 14 24 A7 4C 17 43 1B 26 E7 FC F3 21 33 9E
 4C 7B 28 76 D6 9E 09 E2 56 C9 2A B9 98 EE 3A BE
 1F A0 C6 60 DE 73 B9 AB 45 8E 44 AD 5B 17 FF 4D
 E5 B7 7D 59 19 22 9F E8 D3 C1 E5 0F EB 70 BE 64
 EC CA CA 42 1D 48 43 A4 4F F4 42 D1 6B F0 8E 26
 EC B5 78 CD 66 CF 76 E3 00 DC 0B 14 9C 9D 7E 91
 A0 9D A7 F1 DF F1 78 63 FB 0E 2D 8D D4 7D 5E 2D
 0A E7 67 FD FB 05 7B B9 4B F1 3F 8E 17 C5 70 AB
 7A 4B 7A A7 00 93 C9 67 C9 DA A4 E5 40 1A E0 4E
 E5 5C 1B 40 F4 C2 F3 12 87 DF 1C CD 4F A1 37 F7
 06 2B D0 3A 72 62 A8 1B DF 7E 96 CF EE 29 EF 71
 13 E7 32 70 DB A6 BB D5 CC 19 AF 90 FE 9A E6 D1
 68 A0 F5 6D 6C 6B A7 1F 5F C1 B6 CA BB D2 61 2C
 F7 18 50 0C E9 76 41 52 61 7B C8 82 37 F0 FF 96
 34 FB 58 D8 C4 2C 93 5F E1 05 11 37 65 AD B2 B6
 FC A3 8B 94 28 B2 01 54 5C 35 2A A5 FB F4 AB C5
 5B CE 38 6A 61 0B DC 41 71 E3 12 E1 A6 DA 16 2E
 21 CA 2C B0 C2 96 27 F9 3C 46 42 D1 6B EA D8 02
 81 49 2F 0A A6 18 8E 78 46 A9 37 F6 E5 02 FD 6B
 C7 3D 9B FF 44 FB EF 27 24 63 6E BA A2 70 14 3E
 92 1C 9F 62 4E 8F 95 BB 48 DC D5 DA E4 86 85 04
 88 A5 2F 3B 2E 6B 24 3B 62 69 EC B4 E4 ED 17 16
 FE 8B 55 92 10 9E E7 A1 6A AD 88 16 74 34 3C 36
 A9 DB E8 88 C7 20 7D 53 37 DC 53 B6 A7 2C F2 2A
 64 48 35 56 BD 6E 0C 31 A4 D1 EF D5 5D 15 B1 C4
 17 3A 62 2D 08 47 BF 4B DC 6C 2A C8 79 DE 69 EC
 E3 03 34 6A DC FA 2A C9 17 C0 F8 29 AC 76 9F BF
 3D 99 77 AC 01 37 C6 C6 D9 A4 D4 D3 70 8E 9F 7B
 4A 4C E2 0E 35 80 C6 7F 9B A8 A0 30 67 AC 18 48
 B9 00 3B CC 61 6E C3 99 3E 75 68 75 86 1F 8A D4
 0F FA 4A A4 36 53 A1 6C 8D 76 DF 9E 53 0F 00 83
 3B 46 1F 75 22 51 34 58 63 FF 15 79 E6 E6 09 DE
 C9 52 AD DB 18 FF 15 7F 2D 49 B4 B0 43 A8 B8 E1
 5A 4C 9D 63 CE 34 BA 09 43 A9 17 2A 00 5E 39 0E
 3F C7 55 C7 7D E5 F5 36 B6 35 82 40 68 F9 4D DE
 7E 8F 41 38 1F 22 55 0C 47 81 73 04 78 ED F5 46
 2B E1 7B 80 1E 96 15 ED B3 C2 A0 A9 D8 F2 85 E9
 D6 46 08 31 BD C8 55 C8 AC 6B CF 7F 10 02 A1 37
 88 60 34 43 1C FC 5C 32 A4 8B F2 F8 A8 52 A6 FF
 83 37 09 48 E6 30 8B 8E 03 FD 57 67 13 AC C5 2F
 9D F6 7D F7 46 31 93 FE 0C C8 69 2F C6 AC 35 81
 1D 7A A1 76 BD 6B A5 43 02 A0 BD 04 06 2B 76 9A
 1B C8 EF 97 35 0A 18 06 84 3D 56 F1 BA E5 67 5F
 A8 F3 41 56 8D 8F BD 17 D8 82 06 1C 4C CA 73 3A
 B8 F9 E0 19 4F A8 D9 B0 0E 2D 0B 59 CF 7A AA D4
 B2 96 16 46 4E 07 4E 29 D4 47 66 F3 F1 74 01 51
 7C 5C 2C 62 6C F1 F8 BB 55 DA F7 42 EC B4 C2 6F
 4A 41 49 85 94 CD 47 B3 78 24 2A 12 BA 40 F2 C0
 C0 F6 0C FB 14 5A 1A 90 79 21 A7 50 12 19 2E 5D
 5E DD 11 B6 9C 82 ED FE 65 B8 22 D9 47 58 77 52
 47 2E F4 CD 25 F0 DC 54 95 D9 A1 47 BA F4 CC 1F
 FC A5 2C 2D 33 24 A8 ED F4 A1 9A 9B 15 E4 77 82
 AD CB 95 A7 C4 F6 F4 60 0C AA B2 DF EB 41 3D 3C
 BF DD 0A DF 2C 23 1B 32 1F 9C C1 37 6B 20 08 66
 34 C7 50 0A E2 CB DA 1A F6 9A 10 DB D4 DC E5 39
 10 16 6B 65 E5 B4 7F D4 11 7C 74 19 E8 3B 61 B8
 03 CC 0F C2 2E 91 57 99 5B 99 20 BB C8 27 19 D6
 FB F7 9A 09 8A 0E 2B 1C 83 4D 0D 0D 43 0A 55 72
 72 E5 B6 1B 66 40 56 78 13 68 27 D1 5C 81 19 1A
 C1 4B C7 94 E2 A7 80 84 A0 C4 DB A7 48 D4 A5 57
 74 FF B7 6F BB B7 4B DE 18 82 A1 05 01 AA 9F 93
 BD 49 35 33 81 66 0B 87 D7 F0 52 AB 1C AA 3E 23
 B7 A7 14 90 5B 73 4D 93 DE C9 93 DE E1 85 5E 0D
 CE 59 3A 59 17 14 9C 85 51 08 07 30 15 7E F5 71
 F1 BF 1C 98 10 9D 40 BF A8 86 EC 62 4F 88 95 41
 04 03 23 DA 04 E7 3F D4 7A D6 CC 9D A8 E0 0D 6B
 82 59 63 AF C6 DD BC 22 EA E7 71 EA 80 EE 54 76
 16 73 10 5C B1 01 36 9E 31 67 4E 2E E0 1E 9F 0D
 58 F3 EC 21 BD 9B 19 F0 43 94 EB 86 E3 0F 9A 92
 AF 16 A9 59 D2 5A 3B 92 DE B2 A8 DC F5 1E 23 2D
 BE E7 38 E1 F1 46 8F B4 DE 1A FE A1 76 05 CD 36
 32 18 A2 0B 69 AC F5 A0 4B D3 6A 5F DB 9F 00 50
 19 3F 93 A8 C1 07 BF 3E 84 6A AF F0 4F 38 94 47
 E7 0C 62 B4 73 81 17 D5 74 E9 7A A6 AC 4D 00 CB
 9D DD 37 02 C5 40 72 9F BA CC A2 DD 1E 67 99 16
 60 29 55 2D 0B FF DC 03 9E AC 6A 96 46 6B 1E 80
 FB 9A 3E 67 9B FC 2D 3E 0E C4 3C D0 62 E1 3C 7A
 46 4E 40 2C F4 FA 90 7E EC 15 1C 9B A7 CC 6D D2
 B7 2F 4B 4E F9 80 53 FA 4C 8F E8 C4 34 7B 7C 7F
 BB 7F 5C CE 7F 0A 12 50 BD 58 B4 47 E9 25 07 D4
 10 59 74 A4 DF A8 5E B5 DB 20 2F 45 88 DA F3 2F
 CD A9 77 D9 8E 93 90 40 E2 08 CA 8A 94 AC 93 71
 AE 47 4C AF CB 04 B4 7B 58 09 14 AD EE C5 CC 24
 C4 46 91 6E 05 A8 68 B8 F1 75 DC 21 F9 EA A2 E1
 9D 87 2C FA 1D 8B B1 13 B8 68 30 98 77 AF 1D E9
 A0 FD 41 5D 13 69 76 63 AE C2 49 17 FA ED 31 C2
 0A 69 60 B3 98 72 67 F1 C4 98 B7 E4 FF B8 48 8F
 98 04 48 2B F4 2C AB 8D 8A 54 ED D6 8B 6C B2 11
 34 C4 E9 61 47 D4 CE 17 BB D1 88 41 72 16 E3 D7
 59 73 8C 6F 4A 33 36 17 61 31 8B 8D 46 7A 7C FE
 9B 94 41 1F C3 CA 7E BA 28 1F CA A4 E9 71 6B B7
 AD 07 68 B6 6F 03 69 A9 94 BC 7F 64 49 12 6D 59
 A0 B2 DF 77 E1 F0 BE 28 08 CD FF 77 88 AC F1 5C
 CA 3B 52 E2 66 EF D3 85 D7 F2 3F 1A 0E 5C 20 DF
 4B C2 B8 34 66 DE D8 9C 73 22 50 05 C8 40 4E EB
 06 10 99 F1 2E 30 C9 F5 6C 62 10 7A FB 3B 9B 0F
 9E CF 52 D3 CB 2D 25 E6 BD E6 9B 6D E1 DE C2 A8
 2F 86 04 14 0F F7 6C F5 54 AC EE 13 7B F9 DA 11
 46 0D FA E1 C6 55 31 E7 60 C8 24 A2 45 A4 FF 9B
 49 91 B9 98 32 52 98 D8 5D 95 16 AE D8 D8 94 40
 7B E1 9F DF EC F5 C3 42 58 21 3C 86 25 A2 E1 BE
 20 57 00 C4 E3 51 7E 87 60 03 B6 0E 8D 73 E9 07
 45 4D 68 2D 4E E2 DA AB B5 11 BE B9 FA 51 6F B5
 F4 31 07 F0 C3 E2 E7 7C D2 E3 71 BF F0 39 EA F5
 EC AF 5C 89 F7 D7 96 6C 0B F5 4C 4A 09 A3 66 12
 7C 46 72 1E 4C 2B 4C 0A 04 B4 17 68 5A DB 5E 0D
 F3 C2 67 C5 80 9A 9B DA E0 97 49 C7 10 54 80 3B
 7C EA 3C 8D DE 82 ED 5E 52 54 C0 FB 58 B6 27 38
 6E E8 C7 54 A4 44 6E 82 77 39 3D 00 4F 64 D3 D5
 BA 78 D6 EE 21 80 03 84 B5 23 17 D5 71 17 E3 50
 72 78 EE 6F 0C 66 D4 3C 9E A4 FF 5A 5F A2 20 C6
 03 21 3E 96 17 39 08 2A 4A 87 A1 B9 FB 40 FE AF
 8E 2C BA 06 E0 6D C3 37 AF 00 FB 66 6D EF 6F 14
 CE 8D FE 91 97 07 F9 3B 85 3C 1C 25 95 D0 0D 2D
 14 17 A8 45 62 C1 34 F5 37 D4 BC F1 EB 97 54 3F
 7E 31 4A 8A 98 1C 4F C3 A8 D5 65 C8 D9 C7 53 F0
 4E EB 31 17 D3 36 EE BE 6F 7F D6 2A 97 DE 21 C3
 0F 87 B2 74 7A 42 64 EA E6 45 73 EA B5 2A F9 A8
 E3 97 4C 75 8D AC 48 5A 0E 3E 05 1C CD 78 C3 3D
 70 14 73 AA 08 D8 42 F0 52 FB DC 30 57 A8 79 57
 10 CC 92 8D 0B 45 7F C3 6F 65 89 1B B3 25 62 9E
 0F 02 C8 B8 7A 99 DF 6A EE E8 5C 98 76 83 2F 60
 6C 70 5D AA BA D7 95 DC 21 C1 A3 F9 BF D4 77 2B
 D7 D5 A5 FD D2 11 33 18 7E EF 0A C2 5C 86 2F 4D
 4A BC 4F 87 84 3F 2F D2 56 4D 2C 10 51 42 76 BD
 FA B3 57 18 64 4B E2 53 4E A2 0B 89 74 00 2C A6
 E1 13 95 02 D2 B4 55 65 91 FD 20 FC 01 98 89 DE
 4E FC 8E 34 E5 7D 4D 83 80 66 AA 4E 3C 83 E8 70
 D0 A1 0C FC B1 72 5A 38 DF 91 2A 0F 14 C0 42 D0
 35 2F 01 F8 D1 92 E5 BE 76 52 9F AB DE 49 70 58
 83 36 44 1B BC 49 41 BF 10 58 B2 F8 B2 8C 4C 8F
 32 D9 54 E1 F8 D9 F0 75 8C D0 4A 28 03 E4 5C 27
 DC 5D 30 66 B6 BF CC D1 EF 40 EB A0 C5 D8 3A 38
 B6 C2 C1 DB 35 09 7E ED 2C BF EC C7 A6 83 60 76
 ED FB F2 9D 8A D2 23 4F 72 09 96 2A 6D EF 81 28
 16 5B 3D 38 17 EA 3A 38 33 96 15 C3 37 CA 0E 8D
 C6 9A 63 96 FC 2F 3C 39 5A C9 B6 02 FC EB FC D9
 61 11 24 1B F6 37 FA EF 57 C9 C7 AC 74 11 B2 EE
 A1 B5 13 88 53 8A 7B 61 E4 05 89 2B D3 56 24 B1
 6B 53 6A 57 E5 F2 E1 73 C2 91 42 50 4C EB 00 C3
 35 8E 09 5E 6A 33 65 6E 39 52 E2 7E 6A B9 9D E0
 85 D6 B4 0D 11 62 49 51 AE 43 D4 EA CD AE 16 07
 2F E8 FE 2E CA 03 0A 10 5E 39 7E 8A D8 52 52 D0
 67 87 45 84 10 63 5D B8 7A A3 90 F7 2A 9C F7 5F
 F5 68 E5 BD 39 8C C2 A0 3C D5 4E B0 3E 3B 46 97
 B7 E9 FD A5 17 89 87 D8 5E 07 71 74 53 F0 7D 3C
 B2 08 01 C7 8D CB C6 C0 E3 B6 6F C0 DA DF 6A AC
 55 74 46 CE 45 D0 9C D6 21 D6 06 F3 A6 46 C0 7F
 B4 02 25 B2 BD B9 FA BE 08 E0 CE BC 19 BC 11 7E
 C4 EC E1 A4 15 8A FA 34 2E A7 34 30 D0 24 02 82
 9B 0B 62 21 FE FE 8D 35 02 2A C4 62 9A DE C1 93
 1B 00 B8 B3 C4 97 50 6E AC E9 60 18 C7 21 56 81
 ED 51 B7 CA 6E 54 82 79 3A 31 BC 90 23 AA 9E 31
 C5 0B 7B 8C 6E AD 22 74 22 88 55 52 F9 40 15 76
 E1 4D 46 82 F4 52 15 CA 4B FE CA 7A 01 28 98 18
 AC DB EB 57 C0 D9 B7 EB F8 C4 5C A5 9F 7F 3F D2
 8A 82 29 D4 41 78 35 FF 98 26 EA 8B 3D 3B 08 D8
 4F FF 35 59 1E 42 63 00 71 A2 14 5C EA EB A0 CE
 F6 C5 7E 98 29 82 C9 A1 25 F6 C2 B9 F2 5E 96 7F
 A5 BE C0 86 78 62 8C C2 70 E6 E6 06 3D 6D 0B DB
 97 25 33 79 BE 51 9F 3C 9D 9B A4 05 60 C6 2A 0F
 42 4A F3 02 7A 48 12 68 98 F4 40 97 24 F9 CC 78
 E5 08 DF F2 A9 8F 47 D4 11 17 7A F0 FB 58 30 97
 73 0F 2F E1 B9 04 CE 17 8B 71 DE 71 EC 82 8C C2
 31 DF 0A 50 DB 5B 59 31 93 45 83 99 F5 4A 27 50
 C4 B8 4A BB 65 55 9B E3 FC 60 C7 02 75 DB BF D3
 9A 28 29 56 1B C9 62 A0 1A 12 8B 02 B9 52 A8 93
 C3 A7 E1 0F 2A EF 57 BC 7E 8B 77 94 2D C8 E6 3C
 09 F3 07 76 E9 4D 05 E7 A2 F8 65 6B BA 4A E8 BE
 A8 3C B5 E5 4A 9C C9 4B 97 68 1B E0 8A 19 00 C7
 E1 DF F1 DD 4D 3D 0E E7 35 DD C1 DB D9 3E C1 99
 F4 46 D8 B5 73 45 ED CD 29 FA C2 A2 C2 9B AB 43
 70 07 71 DB 98 C1 26 9A 34 A7 41 48 5D 06 15 77
 2C DB 0F AC 95 A4 61 BB A8 F4 5E A1 37 1F D5 CA
 07 48 F6 A9 AD 59 13 91 E3 8D CA 27 4D F7 35 5E
 1A 31 17 16 8B 6D 25 89 BC 3E 87 83 92 7D 32 4F
 AA 70 CB 9F 46 72 91 DF CF F7 38 39 53 62 32 5A
 5D E9 07 49 8E 47 CD A4 20 81 BB 23 88 39 B8 AE
 55 73 46 AA 21 0C A1 F3 26 E8 DC 17 EF B8 86 15
 3B EB 20 A4 0E F7 83 86 38 0A D3 F3 23 37 7B EC
 AB 0A 0A AF 0F 86 29 FB 97 B6 FA 21 A6 FF 74 8A
 97 4B 57 34 35 A2 C0 FD A0 23 D3 BB 83 2C 93 DA
 A1 F4 16 2F 80 DD 0C D7 85 AE A6 8F D2 86 8C 79
 9D 7F 09 B9 87 8B 83 5E E8 18 2C 2E 1D 16 AD E2
 32 60 68 76 35 CD CF 35 30 76 B2 C4 38 09 58 21
 78 89 94 5B E1 0F 3D 20 B8 2A 7E 54 8A 20 E1 34
 F8 D0 ED E6 05 A0 C9 2A 8E 39 33 1F CB 52 A2 76
 99 E9 00 59 3F E1 06 48 06 7F 52 4A 47 45 CF 80
 5D B5 09 5A FF AA AD 97 5F 93 1C 02 A6 8D C4 CB
 F2 01 51 B7 7C 18 83 F5 14 0C 2F 10 3C 87 71 77
 10 2F 48 CC 90 94 6C B1 71 B3 64 31 06 7A 56 23
 8E 82 CB 51 CC 93 2C E4 AB 37 B6 97 7E F1 90 94
 41 2D 20 FE 6F 2E 2A 8D 01 8A C7 9A 33 86 7C 47
 6E D8 0B 53 D7 05 81 2B 11 D6 F2 EC 01 6E D1 88
 00 99 74 D1 3F 97 EF B4 75 95 00 AD 77 15 DC D4
 B6 D5 54 30 85 0B EF 33 3D 94 BD 4D 1D F4 AC 6F
 C1 E9 22 C7 3F 52 E8 6C 85 AC 37 32 C9 58 DB E3
 8E 99 BF 43 23 D9 03 D0 41 AB E5 75 02 CF 9F 27
 EE 26 45 95 04 29 1B A6 1E EC 60 7A 51 92 11 73
 A2 B9 D0 A5 5C B2 5C 0C CF DF F8 37 26 8E 5A B2
 D6 19 4E EF A8 86 94 B4 FF D0 74 32 8F 24 10 F3
 89 83 4C E2 C5 4E 54 37 DA 50 9C 57 7F 73 21 C5
 08 73 AA EE D6 56 69 4C 34 EF 46 3A AD 07 47 1A
 56 55 64 C1 74 B1 EB 31 E8 24 D9 2D 4D 72 98 96
 B4 45 1C 82 B5 7D F8 E3 10 D8 65 B1 90 50 75 DD
 FF AE E0 EF FF B7 2E 89 E9 26 98 9E B4 6F 8A 32
 E2 50 91 6E 4C 2E E4 97 FB 02 C1 EC 80 9F F4 E4
 79 60 80 05 E3 2E AE 85 E6 D0 62 07 FC 42 37 75
 EC C8 7A CE 0E 7B EF 83 9C 0A 91 20 DF B8 21 82
 04 BA 94 CE 8E 41 75 05 22 F9 C1 0B F8 15 BF F2
 E0 FB 82 10 6C 49 3B 77 52 DD F9 E6 45 5A ED 97
 16 51 28 33 E6 00 8C 7C 37 E8 B8 6C 8A DC F4 B7
 15 05 77 DC AD E1 3E C9 CE 26 8C 54 DD D5 1C A5
 C4 0E 31 22 3C 08 05 44 E7 FB 94 C1 2B 26 58 87
 D4 49 F0 DF 5A 4C 19 C6 2B 4F 54 B9 36 B9 21 06
 B9 E6 67 15 C6 C6 EE B1 5A 46 2B 83 D0 DE 38 3C
 EA DC 08 25 3C 4A 0B 4D C5 25 7D B8 63 C9 92 16
 9A 89 E7 50 92 89 FD 7A 31 47 27 E4 E3 18 11 57
 D5 51 CE 5C E8 8C 24 E4 1C B5 BB 6A DA 58 2C D4
 61 28 3E FA 4E 6C C7 62 29 C5 5F 56 97 D8 5E 3D
 BE 0E 48 E1 7F 60 44 2E E8 8B 4E E5 CE 86 7E 31
 0D E9 ED 14 63 94 16 85 94 FB A0 0C B9 30 11 E5
 CB 38 34 D7 B4 26 BC FA 97 7C 20 A6 15 15 7D 3F
 BD 24 E9 84 CB 83 EC 33 75 A9 66 E2 76 A5 8E A6
 E5 6A 02 28 13 C7 53 D8 67 15 90 99 AC 6D AE A5
 00 45 B9 40 E0 11 03 07 71 02 A2 3F 92 5F 28 6E
 20 2E 31 51 47 E4 E7 37 76 F7 04 BC CD 1F 76 87
 88 63 18 0E EF 24 A9 61 0B 13 A5 04 D5 DE 15 6C
 D5 E1 84 7A B8 32 7B E2 30 8E 8C 86 D8 27 6B 1E
 FC 82 C0 37 D2 91 AC C1 D0 30 1A E2 D8 3F 05 77
 B1 45 6B 6A 9A 82 EC 9F 5A 63 DA 94 AD F1 30 FC
 DB EB B7 3B D9 C2 3F 51 1A 4C 75 DA 95 FD BF A8
 09 BA 59 95 C2 71 4A BD 29 73 98 6D 0C 7A DC 46
 74 6B 1F 9B BA 72 3C DF D1 C1 78 27 F4 2B 45 15
 CB 0D 7D A6 9F 59 DD 99 1B 15 D0 22 6D AD B8 BB
 87 31 BA CC EA 39 05 6C CE CA 65 43 F3 2B D9 6D
 8A C0 AB E8 31 37 15 4B B1 30 FF 7F B8 CF 0B 45
 C5 29 92 AC 78 3A 22 CB 3E C8 80 7C C8 1E 55 CE
 0A A9 46 86 6B BB 24 A4 CA AB 8D CE 12 32 1D 88
 A5 78 AC BF D5 B4 14 94 0C 5A E1 26 51 B2 04 22
 3C 8D 0D F2 9C 34 DE F7 B7 4A 40 C9 60 1B 10 6F
 A6 4D F3 D2 3A B4 B1 46 74 6E B8 3D 31 38 52 CB
 94 83 1F D8 A0 83 7F 46 13 B7 AB B3 8F 40 ED 49
 ED FC 4F 64 67 F9 C3 C8 1C 5A 26 69 EA B2 12 90
 5B 26 AA 30 51 71 2C F1 FB DD F8 DD 7B 73 34 8F
 71 4D 3F EB DD BF 64 0A 84 59 98 1D EC C1 21 B4
 1C 53 E0 D7 EF 4B 85 36 1A 6D 31 EC 3D 0D 14 C5
 4B 96 24 BE 64 45 00 67 0C 42 38 E4 90 66 EC A6
 8D 06 F7 7E D3 92 21 9B AF A9 02 D3 50 80 31 97
 12 A7 0E 8E DA EA E2 CE 04 D7 4F A8 20 13 D6 39
 68 64 B5 7D A1 5F 16 F1 95 E9 05 63 03 B8 C7 1B
 E6 A8 91 55 9C 7D 0F 4B 0B 4C F1 BB E2 FF 2B 7F
 79 47 4C D3 CA D1 D5 10 9F 66 B3 CC FC D6 6C 54
 88 EA 20 C0 D4 BE 9C E8 A8 F9 A4 5C 1B A6 6E DD
 C8 61 36 C2 2B 08 26 73 5E 3B F6 AA 7F 06 07 7F
 BF 58 06 19 C6 85 81 D5 0D C0 AA 77 5B 5A CD 04
 61 11 32 EF 52 31 A9 3E E0 CE CA AE DA FA 25 C0
 D8 BB 38 DA 94 89 87 BA 27 51 6E A6 6A 3B 59 46
 79 9A E8 D9 29 BD 71 4F 19 DA 50 FA 57 FD 1D A7
 F5 7E 0F 16 E6 C1 43 9F 6F B8 06 F1 EE 6D E9 FA
 01 D0 E8 22 11 5A 94 74 F2 62 76 69 CC 4B ED 26
 E3 91 C1 E7 72 B5 2A EC 0D 3D 7A A6 A8 FC 90 3A
 00 02 03 5D 00 1D 67 D6 2A E2 DB AD 94 93 A0 3D
 AA 4A 18 29 6A 2C AC 0C 77 8F 4A 21 04 8D 43 FD
 EA 79 59 F9 10 2D C3 51 71 8A B1 80 05 47 9D 04
 42 0C 08 CE AD 67 E3 94 03 E0 27 12 69 97 FD AF
 93 62 B2 B2 7F 2B 63 63 DA 31 B5 28 07 DC A4 12
 16 70 47 1B 34 80 2F C2 53 41 54 43 FA 78 01 7A
 3E 4A 91 22 55 4D 44 DD 84 BB F4 6C 45 92 F5 F6
 20 17 96 F6 8A C7 FE D5 6B C6 61 3C B5 CC F2 5D
 C0 46 A5 EB C4 36 D0 E5 97 08 D7 EE BC EE 8D 9D
 36 77 3C 2F 89 B2 99 E7 32 98 25 30 97 38 1B 26
 77 71 D2 7A AD D5 15 B3 96 57 00 95 0A 7A 82 5B
 EA DA C8 65 72 2D 77 48 51 F8 E6 C2 8C BD 5C F6
 AC FE 36 1D 16 9A 39 4D D7 30 EC D2 D8 ED 07 99
 4E C1 55 B9 3D F4 AF 78 A8 1E 41 C3 83 A5 41 EC
 5F F8 19 7C 01 0E B9 BB 9E 8A 48 A8 AE F4 A2 B1
 34 2F 82 F1 E2 E7 00 74 10 62 D0 41 0E 89 53 7D
 2A 7F B8 C8 61 CA F1 22 80 2A C2 E5 58 7E B1 F3
 73 8E B4 19 F7 B8 6E BB 6D D3 0D 69 55 59 2A C9
 6F FE B4 25 D5 FF C3 AB 7E BD EB AF 97 96 E0 62
 47 E1 1A 49 15 1A C5 3D 77 5D 51 99 71 DB 14 FA
 AD E0 38 B4 B4 24 BF 93 16 45 A3 16 E6 96 F1 C0
 B6 86 C6 0D EE 90 95 B7 D0 29 3E 16 3F 82 48 06
 CB 39 90 9E 4C 9D 7C 62 D3 CB 6E 8E FC 92 A6 5F
 F5 9B 12 99 A5 1D B6 08 9F 07 BB 5D AF 4A D3 F0
 3D 9A 8B F9 C8 17 60 A3 27 E8 32 84 48 AC 8D 90
 8C A2 F6 3C C8 71 DF 03 0D C5 CC 25 65 4C B8 BC
 F4 94 E1 63 30 88 D5 36 71 08 E1 F7 B1 B4 69 3A
 8C 74 90 D5 4F 0D 16 12 ED B1 7C F7 B7 70 25 54
 41 5D A5 14 32 7D 2D 8C 33 7D 43 05 92 0B 92 B6
 4B 94 EE 2F D5 8F 00 48 5C 00 E2 BE 66 DB 26 15
 D3 76 53 92 A3 F9 73 E8 E9 B4 9B 14 C7 7E 76 F5
 C6 42 D8 55 AD A6 BF 85 6A FA EA 28 E1 17 CE 06
 DD CD EE B0 DB 40 F0 23 A3 84 07 06 56 2F 4E 72
 7F F5 99 07 8D C5 E2 F5 DF C2 BD 4A 7D 76 4B DD
 8E 21 FE C6 2E 41 7E 30 73 39 0A C0 98 F3 A5 8A
 FE 4B 27 1C 83 0F A6 88 09 51 B7 68 63 FD EF 7B
 D1 61 2B 9B 24 2B 68 30 B1 DE B6 A1 69 DB 39 F6
 EB F4 42 11 0A FA 12 0C EF B5 78 D2 6B 14 7E 08
 52 CA 76 E2 D6 C5 AA B4 02 1E C8 95 34 F8 DF C3
 3B 06 70 28 93 7B 5D A8 8B 36 4D 65 D2 75 86 CB
 E4 64 EB 3C A8 D0 A9 E3 CA AB 71 2C 97 6F 64 E8
 FC E5 05 A0 10 E6 FE 5B CB 9E 51 1B 91 22 68 F0
 EA 7B B0 CB AD DF 3C C9 21 4F A1 88 07 A0 7B AF
 AB 3B 8C E9 ED E2 C3 DB 61 43 FA 47 1B 9F D5 0E
 22 6D 43 AE F3 B1 02 F3 73 BA BF 13 06 72 88 1C
 DF 37 18 B6 89 F2 77 60 EC 9C D5 C1 CB 0A 0A 7D
 EE E9 4A 2E D3 7A 09 59 7A 8C E8 10 43 F8 C1 18
 31 78 5F F6 AC 47 C6 6B 3F 81 86 60 AB A7 EA AB
 BC B2 16 6A 3E DB 2A A6 88 00 C8 A6 A1 57 78 41
 07 5E 37 E9 28 FF 4F 0F 33 41 D4 CA 0B D2 8B 1A
 89 38 02 A8 04 19 19 9C 1C B4 71 60 24 43 B1 24
 4E AD 55 C0 7B B1 CA CE 75 64 B0 D6 7F 05 35 CB
 A0 67 91 38 19 C3 C4 3E A1 D3 E8 E8 E4 6C E3 22
 6B 3F B9 DA CD 7C 4A E6 E1 45 40 A7 A2 A3 0B 91
 E5 D7 C0 81 E1 50 5D AC B2 DB 77 D4 83 D4 E1 80
 19 99 16 60 C6 47 4E 2A 06 7C E6 95 BF CD E0 21
 23 27 8C 45 9E ED 6B 59 F8 9A EB CE 10 05 4B 90
 EF 6A 13 D5 F0 53 53 52 48 6A E8 34 4C 2F 79 77
 F0 D9 A3 C4 F7 17 1D 27 A3 04 38 36 4F 2B E5 42
 EB 9F 47 55 02 24 CA 01 B6 41 FE 59 71 0E D9 58
 EA 6D 4C E0 57 D5 5C DD BF 8C 18 C6 CC B9 D2 CD
 04 96 C6 C2 62 CD F6 CE 8B B7 1A 18 91 15 CE 10
 1C AA 1C C1 0E 0A 46 22 1F 02 10 6A F3 83 F9 2C
 AF DE EB 6C 6D 2B 90 35 AD CB 76 AD E9 9E 81 FA
 A6 31 06 46 A8 B1 B5 0F 6F C3 09 32 F4 9D 4E 6F
 B5 E2 42 54 AC A5 40 F7 99 FB 9F E6 8F 03 D9 21
 D0 77 AD 6D AA 40 DC 2E 38 BA 43 25 D5 13 83 FC
 08 9D 2E F4 8D 4A 6E 29 AA 30 EF 80 A3 4A 89 7E
 80 75 E6 D7 EE 2A 0C 41 F3 ED 67 22 3E 54 93 54
 E7 75 0D 10 7E AB 6B A8 11 AB 4B 7E 63 69 0B 32
 10 44 DF 16 2C E3 00 0A AE B5 4D 02 61 6B BF AF
 0F 3F 4F 1F C9 AD 3C 84 F6 2F B2 79 55 56 89 55
 7F 06 F8 C6 E7 13 B8 FA 40 78 60 67 C5 DB CC 9D
 19 26 EA 75 57 17 7F A7 AB F0 C8 B3 AC 92 98 02
 4C DC 95 DE 74 F4 27 8E E7 4C EC 10 B9 56 73 EC
 4E 7B 44 63 46 CD A9 73 5A C3 29 E9 D8 C4 F2 A5
 18 8D 3D 3C 18 BC D6 F3 C3 73 9F 06 49 D0 95 20
 BE 3D 34 33 9F 7B 46 0F 41 CC E7 B2 38 66 0B 78
 0A 19 39 29 04 A9 D1 65 1F F8 40 51 77 BE 78 1C
 9F B6 3D 8D C4 62 A1 B0 DE 69 AA FF 99 CE 3E A2
 CF 58 03 1A 28 30 C5 A2 F3 06 6D E3 A6 50 A2 4E
 8A 7C 20 66 C6 5D A0 1A 48 B8 66 B0 0F DD F7 C0
 DE 18 36 F6 A5 27 9B D3 BD E9 7B 39 2C 58 C9 E2
 37 87 42 70 97 CB A7 04 79 C9 DD C5 C0 0D 88 A8
 9B 03 C7 56 1B 85 7F B2 A4 04 CE 3D A6 36 A1 D6
 A3 33 D4 82 DA D5 F2 20 BF EA 04 97 9B 81 D2 A6
 E7 6E AB 20 50 74 93 EA AE DC 60 36 A6 F7 69 16
 FB 5B 88 2A D6 DF 83 57 11 C3 C0 92 78 60 8E 97
 CD 15 77 CC 10 06 C9 4B D0 9F 21 E1 C6 F0 3E 4C
 08 49 1E BB E4 5F 40 24 46 E6 79 61 A9 0B 56 AA
 C3 B0 5F EB 94 87 65 34 81 CC 4A E8 9D F0 69 BB
 29 75 1D 72 66 38 21 9B 88 19 19 3C 42 FD A6 C5
 3F 51 83 2E 3F D7 5C E2 51 19 AB E2 10 EF 97 8A
 2A D0 58 DF 7B 88 20 B8 57 79 D5 21 8D 23 3C C0
 62 1D 5D F5 C7 39 D9 19 DA 6E 44 B7 51 23 7D 3F
 62 72 12 CC B5 A8 D0 DC 36 CD B6 89 E4 13 32 36
 AD 8A 47 4C 80 52 E3 AE A4 7B E2 66 27 E6 CB AA
 CC DD EB B0 E0 69 5A 78 06 1B 82 2D D3 82 04 E5
 FB C9 C1 35 C6 54 DC F6 FD 31 24 20 2C 2C ED B4
 CA A4 97 58 32 E2 7F AD 90 77 39 F4 21 C2 A8 86
 BE 56 F5 9A 60 71 3B 04 B9 85 85 D8 A9 79 76 4B
 7D 7E B8 D6 EA 95 1E DC F4 03 F9 C3 08 61 2B D0
 E1 2F 2E 8A 8D 68 64 E5 D8 46 3B 47 5E 9A FE D6
 76 F6 81 4A 3B 2E 88 DA 2A F5 19 29 36 EB 40 8D
 1E 3E 92 46 C1 69 73 A4 E1 5C 45 71 68 3A F0 12
 52 9C 03 7D A3 D9 01 FF FB F9 73 B2 91 F7 54 D0
 E0 94 93 B3 73 EC D2 99 3D 8A 7E A9 89 C2 44 FA
 32 D7 EC 7C B5 CC E0 E1 4F 8C 4F B5 61 5D AF B5
 1B 2C 75 9D 3B EE 47 9E 2A 86 92 A1 EE DF EB 43
 C9 BF 12 4D 16 62 47 AB F0 17 17 71 01 EF 38 42
 34 55 EB B4 46 AB 05 8E F1 7F 81 BB 32 19 0E D3
 9C 56 72 EB F2 5C 1E B4 5E 0B 63 B1 1B DE 4A AE
 5A 39 E3 52 B3 91 EA 2A 99 B0 07 C1 8B 21 1C 2D
 33 CE 73 6B 44 52 E6 29 EB 8A B3 46 CC 6C 5A 3A
 B0 5C 10 FC ED 4D 43 BB D1 33 33 58 E5 1E DB 4E
 D0 12 7F 67 EB E8 31 A5 58 C6 F4 AA F5 36 75 79
 58 51 3A 8F 18 1A DA A4 63 3E A1 EB E3 68 D5 64
 C8 29 62 4C FA F1 0A D9 08 1D 60 77 22 3F 63 A4
 CA E2 46 C8 1F EB 50 50 66 82 B8 A2 FB D7 27 BA
 D3 49 68 D9 4B 72 85 42 79 E4 39 EA 24 63 BD 16
 D7 89 19 B0 FA A3 3E 5F 13 64 A1 18 DA 31 FD 60
 4E A8 54 8A 94 25 62 4A 39 50 73 A3 D3 7E A3 54
 FA 2E 9C B4 C8 96 F7 D0 F5 05 2B 23 3D 11 F4 25
 5E F1 27 AF A7 EB 22 AC 1D 3D DD B7 71 F9 2B 16
 8C AF E8 AA F8 14 28 13 FD B3 B9 48 FD 0B 9E CD
 92 B9 E9 70 C4 9D A0 17 E8 7B 05 65 A0 D3 21 F8
 11 B8 F6 E6 28 01 98 26 E4 A9 C8 31 51 55 98 2A
 25 44 C9 C0 90 C9 4D 08 62 82 A6 4F B5 37 AA C8
 F2 9F 31 E2 87 A7 B0 CC 4C 71 1D F0 8A DD 4C DD
 69 5C 63 F2 4D E5 1A 33 33 BF 96 63 4C D5 57 7E
 5A EB D5 20 E0 81 51 56 4C 43 62 52 82 5A 62 A9
 CB 93 30 B5 A1 BC 28 19 E9 8F 69 C8 43 A3 44 39
 C8 0A BE E2 E3 7F A8 C5 D2 70 0D 60 80 58 0F 09
 24 7D 80 84 98 44 AB B9 EF 39 47 9D 30 A7 D8 6E
 DE 16 AC 53 69 23 4D 76 85 F4 A4 AD 01 AF 94 B4
 16 06 C2 B9 86 33 E4 FD 0D B9 0D C7 81 39 A9 4D
 A6 61 1B 1A 02 5A 50 69 59 50 99 9B 43 F6 C2 BC
 27 0B CF 3C 78 F2 6E 33 46 DA 8B DE 0D 7E 3F 5B
 16 3F DE 4C C2 8F 2E 5F D0 B0 31 B1 C2 F7 CE 29
 65 87 77 3C BE 41 C5 7B A6 6F 06 83 9C 8E 14 24
 7B 27 E6 C9 2D 19 48 7D 1C A2 AC FA AD EF F8 E1
 DD 94 A7 E9 FD 26 16 94 9E E2 2E E8 EC A1 9C 53
 F6 9F D3 D5 A7 9F 78 7F E3 B9 9B F9 08 01 BC 08
 3E 0D 78 07 A0 31 04 5E 15 C6 A7 B9 02 F2 6B 70
 56 89 B2 EA 8D 58 3C 23 B2 34 E1 0F 88 BD F2 97
 5E 90 46 0F 82 94 4A D9 37 6C 35 B7 FD D5 A4 BF
 95 E6 8E 2C E1 76 E3 9F 69 1E 64 17 0F 1C D2 00
 0F A5 39 2F E2 D9 A1 2C 05 66 AD 40 AD B8 11 A0
 A7 9A 34 48 AC B0 20 CD 12 FD 5F C9 FD 1E F2 76
 F2 C6 E4 CF E0 23 70 D5 E8 99 C6 63 50 BE A1 AB
 41 A7 7F 5E F5 47 F0 89 68 D2 47 C1 13 DA 40 53
 AD 98 DD 67 20 2D 9B 89 6F DE 71 EE CB 70 85 73
 29 15 23 C8 82 BD C7 6B A3 0D 3A 0D 78 57 78 99
 F1 38 7E C6 38 9F CB 63 47 19 B9 63 B5 30 10 F0
 E9 EF 9A 2F 5F 00 8D E7 4F E3 2E 09 02 F7 BE 4D
 87 94 68 72 23 FE C0 B7 A3 16 A1 76 FB DD 89 02
 2A A0 B5 C6 BD 6C 8C 6A 38 44 94 E5 60 83 48 CF
 2C 8C 16 B2 EA 8B 2E 31 5C 08 AD 59 32 E3 F8 0E
 41 38 21 F8 1A 29 96 5B FA 79 80 32 CB 55 4F 22
 15 41 86 F2 F3 8E FF 49 7D 3B 01 97 7B 7B A9 A3
 25 BD B7 D1 B1 3B B4 E9 AB 33 B6 AD DD E5 E0 7C
 A6 FF 97 63 B8 78 9E D4 91 07 02 D2 C1 B3 47 B3
 72 4E A2 62 C7 77 17 93 33 04 F6 6D 81 FB C4 12
 B3 3E 30 91 D2 DF 1D D0 7E B1 FB 46 51 87 D6 B1
 CA D5 7B A8 F6 DE E7 E6 C4 7E AB EF 40 10 EA 2A
 64 85 68 33 F7 36 C1 39 BC 23 3F 77 4A 68 58 1E
 08 BB 7A 26 8E 81 E3 CE D1 33 6B A3 CC FF CB 83
 B5 52 E8 7D F8 99 56 85 22 68 0B CD 40 E4 CD B2
 81 F2 47 76 94 CB D8 F3 DE 44 DF B4 66 6A 47 C0
 B2 5B CE EC D8 FA 15 64 26 9E A4 22 FE 16 74 1B
 4E 4B 25 B9 E9 3D 5F E6 33 1C 5D AB 76 61 B4 30
 CA A5 3B 78 15 6A F7 5D E2 E2 E0 56 67 1B 1D FC
 F2 64 F6 AB 08 FE 4D CE 86 FB 31 8E B0 D4 9D 30
 82 4D 75 1B 9F EA A8 D4 84 A0 A4 0E D9 44 45 9E
 15 91 13 BF CE 62 C9 B6 37 57 D2 E4 00 BD 18 FC
 95 1F CF 0B 34 30 87 FB C5 9A B8 67 79 FD B5 62
 E0 C4 E6 B4 C6 9A 6A E7 6B 8D 2B ED D3 6E 63 73
 5B CA 9A 2D CA 34 7C 1E AA 1C 5A A2 49 77 AE C1
 DB FE 29 79 3E CB C0 26 7B 29 55 09 DD 76 7F 54
 5D 09 17 ED 1B 81 C0 FC 24 DD 91 12 D0 D1 C6 77
 93 9B 60 A6 B0 BD 93 8A AF 09 EC 1B D9 8F F0 57
 BB 58 97 C9 D1 CD 52 96 65 A6 38 80 A5 4B 3D F6
 69 64 E5 C4 CA E8 CB EA 1A 83 62 87 BA D1 48 30
 58 6C 8E 89 99 D2 A6 CB 88 2E DF DF AB 91 8B 92
 80 9B F7 4F 2C 95 29 75 4E 49 1B 5D AE B0 BE 1F
 3C 11 DA 77 32 1A CE 84 0B BC CF 70 98 43 57 4D
 FD EB 72 79 F5 D7 04 4D F0 2D CE FE EA E0 D7 80
 54 76 2E 0A 52 A4 A0 C0 0F AC DA 9E C3 A3 5E 19
 10 42 9C 32 13 74 91 3E 85 D0 E1 AB 56 16 0F 94
 37 5D 69 B5 03 40 A1 02 44 74 A7 72 48 89 10 52
 32 2F 70 77 60 B7 78 45 B0 8B B8 2C A5 6C 01 7C
 65 2D A0 4A 60 4A 9A 57 DA 7B F5 0F 91 2B FA FA
 F6 B1 08 9A A8 71 29 B8 A3 08 60 F2 46 24 12 58
 D7 38 78 01 E0 16 77 90 11 3A 7D EA E0 6A BF 44
 06 D7 A6 D1 A4 D5 F6 A2 96 1A 63 DB AD EB BB 08
 52 CD E0 64 FF 10 A2 FC 1D 50 23 BD 28 27 1E 98
 50 D5 27 14 47 E6 5E EE AF 1A 66 64 0F 90 CE 2C
 64 C4 8D 87 48 81 C1 87 A1 6D 65 55 A1 79 6C 27
 83 B7 AF 6A 26 D2 E8 E5 E6 8B 23 E3 C0 6E 8A 14
 92 6E 18 59 AA B9 8C 43 90 AF 2E 04 72 2A 26 E9
 C5 E9 83 4B 03 16 18 60 6D 9E CE 76 4D 10 7E C9
 98 7F A7 54 37 C4 60 7F 22 9A F4 4D 2E 21 A7 DE
 29 F2 D8 66 4E 5D 02 12 9B 80 2E 0F 4F 37 8B 09
 C4 FF 4A 06 FA BD 42 EC 3B 7C 57 BE 11 7F A1 F0
 08 23 96 05 36 49 E6 03 67 F5 BE 25 8C D1 59 88
 52 24 4E F7 87 A6 30 3A F1 20 AA DC C8 96 11 36
 77 2C 0D 97 68 9D E5 AA A9 B5 FE A4 73 7B 27 7A
 31 2C 49 C0 87 CE B6 8A 02 89 FE 95 7E 72 D8 BB
 B1 D9 51 D0 EA 1C 6C 26 81 61 AE 87 E8 5D E6 E6
 2A B0 C3 CE 4A B9 14 C5 58 7A 84 72 DC 80 ED 35
 22 37 B3 58 2F 6A CA 8E 2B 71 92 69 12 E3 23 05
 D8 D7 2D 82 99 C5 3E 7A B5 7D 29 26 50 C1 DE 4F
 2F 47 E0 16 38 EF 20 B1 73 6F F8 8D 45 34 35 45
 98 14 D1 6A 6F F1 28 95 1B 67 2E 2A 2A AD 76 91
 7B 78 31 F7 49 3D C5 20 0A C8 AB BA 6E 6B FC C1
 7A F6 78 AF A8 DF EB AF D3 B2 13 83 38 90 4A 88
 3F FF 34 B8 0E A9 DD 94 88 64 B1 37 10 E4 C2 85
 D3 06 3D 96 26 3E E0 12 B4 56 06 38 34 CB 6B A5
 1A 9E B5 92 54 5D 89 0F 69 49 D0 F3 31 FF 87 1C
 49 0E 7C FE C2 19 1B A1 FB 65 9B CA 78 0E B5 87
 DF 08 2F 79 63 06 E1 A9 36 EA E7 64 88 BD 1F BF
 32 DC F5 00 2E FA 0F 0F C2 19 90 53 EC D3 C6 BC
 DD 1A 8E 38 9A 9E DD 42 D5 00 4C C6 80 53 E8 A4
 8C 59 57 40 50 E4 2A 58 86 C1 F7 B0 97 64 42 E5
 C5 C3 A8 A0 E5 7E 98 5F 82 8B E0 AC F0 6D 65 94
 0E 5F A7 47 BC 6F AF 99 86 70 57 F0 D5 8C FF 42
 9F 2C 16 90 DA 0C 76 1D DE 46 E5 BA 4A 80 61 AD
 7D 2C A4 BA D1 20 66 8F 13 0C 9D 40 D8 0E 52 BC
 82 86 C5 CF 6A DD 31 57 59 6D 71 58 C5 F9 90 9A
 6B 0F 93 EF 44 82 2A 91 7A 1A 34 48 20 01 FF C9
 72 52 1D 90 78 BF 63 F8 48 67 B5 D3 7B 05 2B B9
 A7 D1 62 E6 80 BA 64 B5 28 DE B5 D2 42 D6 28 BD
 38 0D 87 1A 86 40 DA 0B 03 46 0B A9 70 53 CF 5E
 11 8F AF 9F 69 B0 8E 00 9E 53 12 57 7F D8 C3 60
 27 BE 96 D0 8A C3 CE 96 C4 4A A1 A4 50 39 D3 5C
 69 A6 AA 91 CB 11 CB 39 6E 41 5B 0F 3D 14 A4 5C
 77 48 E9 04 8B 08 2C 74 A0 68 50 11 92 8C D3 83
 2D 97 E1 66 24 33 AF F0 98 E3 AC 79 95 96 E5 15
 F7 FA 4A 92 71 CF 9B CD 39 98 C2 86 B7 8E 7C 8A
 F5 B8 12 B2 E3 71 86 0B 7B BC 55 20 F2 6F 7E 95
 E1 74 54 48 F1 B4 A4 91 9D 21 26 34 CD 8C 57 AA
 44 F0 8E 2F D5 B5 0C 4B C0 5F 64 C2 D7 35 F0 5B
 F3 2D E0 DB 86 17 3C 00 76 6E E9 92 F3 FE 54 38
 4B 41 2E D2 35 7E 38 92 EC 2A FE D0 D8 AF 5F A7
 8E 0F B6 86 20 8A C2 F5 D8 0D 96 E5 EC 9E 73 D5
 D1 CA D9 9E 40 90 8C 1E 74 72 67 18 B9 63 9D 4B
 BE 34 11 73 39 25 BE 76 56 61 AA C5 DD C0 A1 2F
 B7 C8 D9 54 C7 4D D0 6F CE 78 32 51 F0 A0 6F FA
 D3 78 FA B7 2E 4C CC BF 7C 31 C5 5E 08 6C FB 60
 7F 33 EA 39 ED 1A D2 BF 4A 0E D5 F4 4F 59 EB EB
 00 30 77 ED C3 E4 17 FD 95 85 5D 52 D2 97 E3 EE
 B0 12 78 AB C5 C1 AA B9 06 9A 86 67 40 B4 26 3B
 36 2D 1C B2 62 A4 05 3C 63 1F 01 F2 30 33 1B 51
 AB 9C 67 31 17 4A 83 0B C6 46 92 8C 14 8C 14 33
 F8 E0 49 4A 70 03 0E 20 33 4E 95 62 F4 D7 7E DE
 45 40 D7 05 9F BB A4 2E D7 76 4C E3 F4 38 33 C7
 12 F9 3A 91 D0 63 A7 D4 FD 8B 4B DE 6F B4 40 1F
 F6 BD CF 74 BA 9E F3 C9 DB D3 8A 74 67 66 95 6D
 D1 0B F8 B2 1D 95 C9 8B 35 7F CD A3 0B AF 87 35
 8B AC 78 FE 6C F5 DB 0E 7B 21 80 E3 41 C6 7F E3
 02 80 D8 8D DA BA 72 0E 16 7A 33 44 CC D5 ED 6B
 69 36 EB 6A 5B 9E 29 F9 6B 99 68 61 D9 FF A2 B3
 21 B9 F9 1A EF 5B 9E 66 D7 24 8D BC 43 09 79 2F
 0E D5 61 4A 52 42 C9 60 81 73 94 97 AB 9F 79 51
 E5 EB AB 50 D3 9F 6C A2 42 14 FE 14 6C 75 6D 89
 66 10 3F E1 53 0D 21 0F 6C 0B CA 21 D9 BE 4D 25
 01 06 ED 3B 38 0C 78 37 00 D9 84 55 69 BA 37 6F
 D8 8E 37 57 65 5B C6 17 86 A5 DE 36 5F A2 8B 47
 62 5B CE 62 01 AC 6C 2D 6B 8D CC 26 DB D2 49 9B
 0D 8D 0E F6 E7 CA A3 09 1F 74 2D 5C CF 5F 7C 5A
 14 61 60 AF CC 87 A6 73 E2 60 59 34 CC 9D 89 F1
 15 1C 39 93 99 0C E4 2A 7C DD C9 7E EC B3 BA AE
 55 C7 A1 FF 86 BC DE 41 92 6C DB 89 E3 A2 02 A2
 32 20 46 B7 AA 45 C0 7A 15 50 AC 96 54 C8 0F AA
 01 1B 4F DC 58 B8 2A 56 38 D9 92 B7 E0 F8 69 B1
 9C 1D 66 28 F0 70 87 2A FD 54 1A C1 A8 BA 6F 78
 CF 8A EB 9D 77 1B 47 30 2D 51 AC 66 64 B4 43 67
 A2 2F 65 0D 23 B0 1F CE 89 AE BA F7 72 BD DA 59
 18 FB 94 0B 89 41 86 19 87 DA E8 C5 25 92 A2 0D
 3F D2 E3 70 07 AA 26 4A AA 77 C9 A3 CE 58 45 A9
 89 96 4F BF D0 A6 3C 9F FB AD AD 1F EF 6C 26 DF
 25 34 00 53 9D 2B 71 6D 5C 1E 73 45 D0 1C 17 BD
 05 AC 93 AE A7 26 38 45 FC 69 09 83 B5 9B 1E 24
 05 2F 0B E1 0B 41 74 DF 6E CB 94 0F B2 A7 20 0D
 0E CE B7 86 F6 FF 3F 76 92 E9 1D 75 1E AF D4 9C
 7D 5E 24 2F FE 29 AC C7 42 0A 30 C4 BB E2 C8 9A
 3A A0 C6 F8 61 99 23 41 AB D2 14 84 B8 B8 9A 1A
 21 FE 49 B9 B8 0E 16 2A 85 B9 E2 D9 E8 8E 2E B9
 1B BC E3 F3 80 A6 32 AD A0 4D 39 DE 75 93 D9 A2
 3A FA ED 38 47 09 3C 9D 73 A2 24 32 4B 07 9A 7C
 8F FF D1 3E C2 F8 EB 94 66 2D 9E 3C 4E 95 7B 22
 70 56 C3 C3 E9 F8 C8 43 1C 29 8D 5D D5 C3 CB DC
 2D DB D3 A2 FE 1E C5 1C C0 60 BE 96 45 A7 71 86
 9E 49 EB 2D 1E 0D 0F BC 23 CC A5 E9 87 33 99 9C
 59 95 59 C1 54 27 9A D7 2B 15 82 E5 0C 8A 7F B4
 F0 B0 00 37 1E 05 EA 12 FC 55 A5 02 4B 2F 27 F2
 99 93 49 97 E6 6C 54 70 A3 17 28 94 12 4D A7 6E
 A1 49 7D 70 7B 52 9B 61 17 74 C1 79 32 6F E6 DA
 22 48 D4 87 68 8C AC 7D C0 3B 53 E4 F6 63 D0 66
 11 28 11 19 14 A6 6D 0B 3D 68 18 61 9B 4B 00 D7
 40 2F 0F EA 6A 07 C9 8E C1 92 BA 13 D5 86 6F CD
 64 60 29 4D AA 8D FF 09 73 4B A9 A7 24 9C 46 47
 FE FC 06 67 2E F1 41 13 05 B8 9D 27 3D 73 E1 79
 94 FA A8 27 27 59 07 0C 64 9E A5 F0 3E 4A 7C D6
 4D EA F5 4F EC 1C 5C F2 57 5E E0 1D 3F 76 78 FE
 B7 34 40 34 66 08 DC 30 24 C8 2F F5 22 A8 1C 64
 AD F6 92 26 EC AA 5E 9E A9 8D 1E 4A 1F FE 62 5C
 76 49 80 20 31 8C 29 28 4F CC 6C F1 C4 B8 B3 04
 1E 59 07 33 F0 4B 1C 7B 57 95 C4 DD C5 56 6F E6
 D1 77 69 2F A0 89 6C 56 13 0E 12 C2 37 D2 E6 8B
 0D 7D 00 52 0B 45 E8 35 B6 F0 D5 5C FC 90 2E 1A
 4D 82 C8 85 3A 8E 47 CB 5B 89 45 A6 2F 7E A0 14
 FC AA D2 B0 9E 3B 1E 37 7E 8D BC DF 18 E5 BE AB
 E6 3A 6B CB F5 D4 6A AA C6 CF 8E BB 15 07 D8 0E
 C3 09 4D 86 63 00 46 6D 8B AF 48 45 B2 8A 0B 9C
 4B 30 77 B9 C0 92 5A 98 64 EE 0E 2D 7A C4 49 5D
 D3 92 15 C3 7B 5F 21 FC EB 79 49 D1 1B 32 B7 9D
 97 CD 24 EE 18 E5 7B 08 91 AE 92 8F 8C E2 C0 93
 ED 69 9F B2 41 FB 8E 63 2F F9 AD BD 63 0C 48 D5
 CF EE 76 30 8C BE 24 0F A4 51 4C 94 F3 09 BA 8F
 2E 54 8A 1B 54 D7 E2 78 B4 F8 3F 9D 99 1E 88 A9
 CA E7 76 D3 93 E0 6B A5 FD EE 3E 5F AA 69 F3 3F
 91 51 D1 43 28 7C 1D 7B 56 FD 4D 57 B3 BC 8A 4E
 54 96 90 CF A1 5F 7F 39 1A 7E 6E A7 27 9D F5 29
 51 B8 B6 A9 4B F6 E7 35 AE 96 05 F3 AC 31 14 E2
 F5 44 91 B7 19 78 97 A9 53 65 FF 88 FD A8 21 4D
 4A C0 53 8D F6 A1 B4 98 78 84 6E CC 7E C8 DD C7
 03 B3 75 E6 63 D8 F2 4C D1 E7 55 79 16 3E E8 1E
 13 99 CF F3 E7 CF 31 BB 27 B7 30 C4 A0 24 A1 C8
 1C 83 3B 63 65 1C 9D 54 7D 91 7F 82 05 5F 64 B9
 69 B3 57 50 4B 91 54 C0 37 6D BB 9C 93 07 C0 B6
 94 3D 28 F4 0A 6E 9A 93 CC 3F F2 A0 4C B0 F7 2E
 87 A8 F3 6C EF CE 3A F3 51 92 EB E8 1E A4 D1 D6
 26 D2 8A 8B 16 CB 42 F3 C5 F4 1F 88 8E 64 3D E7
 6B 2C DD 2B A2 C9 7C EE 15 D8 02 D1 B8 1B 2A 54
 69 EB 65 A4 FB D5 6C CF F1 D9 2C B5 EB 11 A4 51
 82 E4 C8 F6 50 02 E6 2E A8 9F 47 79 69 6B CF EB
 1F DB 3F 08 3B 09 53 0C 73 A0 F1 10 BC 58 2E F4
 BB 5F 39 C5 49 C2 3E 84 CA 36 6C AF 8D 71 67 57
 BA DC 94 91 F6 56 FE EA B9 9D 50 34 97 C6 28 6C
 CF 09 98 2C 09 0F 6E 26 A1 C2 AF 0E 7B D9 7C DB
 0C D8 24 82 F5 5A 86 3B 5B 94 F4 50 C4 BA 3B C3
 D4 80 AC A1 CE 29 6D 5F 60 CC FD B6 18 E7 18 49
 31 31 25 AD 2E 75 50 FC 00 59 66 F9 80 AB C9 21
 85 D9 52 4E 8E 17 3A CA 02 96 B1 55 48 EB 00 5B
 4F BD 26 E0 66 F6 88 44 19 0F 0D B1 0E 4D 42 AA
 2D F0 DC FA 7C CC 0D 9B 41 54 8B 02 7F D8 37 03
 45 9C 9D 83 9B C0 0F 7B F5 39 E4 E9 C2 2F 58 8B
 EF 05 16 6F 15 08 77 B5 4D 54 5E C0 4E 1F 0B 79
 9F A0 25 BB 65 34 63 BA 4B 16 52 E3 61 AB BE B7
 48 5C 6B 6B 36 13 1A E7 C2 54 61 CF AE C9 2D 9D
 F4 C3 D4 47 02 43 CB B1 B7 BD 9F FF CB 35 A4 AF
 B0 1A 0F 50 CA D5 40 C5 B5 DA 44 FB 99 0D BA 60
 8D 47 31 3A 38 C1 2E C8 26 05 1B C3 BD BA E9 82
 BA ED E0 5D 48 BB B0 68 FF D1 C7 EE 7A DE EB 0F
 D1 FA E0 A8 2D 19 52 12 3B 8E 88 5C CE 1C 2E DB
 C3 8E 98 3E 70 46 66 10 80 CC 23 67 C5 0F 8E 5F
 E7 84 5F F3 E7 ED FA 8A B2 3F 9A 3B F1 34 09 B0
 91 7A AA A2 65 32 76 6F FB 05 19 C2 9A FF F7 58
 76 27 29 DC C3 18 49 F6 92 3B 68 EF 68 30 0A 82
 E0 A8 40 E6 EC 09 0C 8A 07 87 9A 98 6C FF 80 9C
 0B 66 84 04 B4 2B DF 44 A5 BA 02 E9 39 35 27 DF
 05 C5 40 3C C9 49 A5 AB 99 86 1D E8 50 8F 2D FA
 CA 16 BC 2C 93 F4 61 2B 99 92 CE A9 EE C2 97 E6
 73 24 81 AD F0 43 EF 8B 49 13 35 AF 77 B7 95 29
 D6 9E 54 7C 93 C3 9E FB C9 20 B8 65 61 D7 3F B2
 F5 C0 FB A5 DB 87 E7 D6 3F 1C 76 C1 2F 79 2F 73
 AA CE EA E7 3F F9 F8 CC 48 D7 A0 FF C6 5F 00 70
 43 DA D9 39 A8 17 CD B1 59 76 8E 4E 58 41 CA E4
 DC 09 39 88 21 C6 8F E3 4C F6 0B CF C7 6D 8D 06
 85 6B 4D 6B 1C 32 85 BE B1 7E C8 58 C4 84 BC 6D
 08 8D 8C 0B DA 40 E9 D8 D8 D1 51 E6 9D 7D 8E 6E
 F8 E5 D5 E6 7C 58 75 6B 6C 9B 27 72 9E 01 92 65
 24 00 2B 20 F8 3E 2A 86 D3 87 1D D2 3A 1B 2D 8F
 3F C1 03 3C EE 2D 45 8D D0 DB A1 41 D7 55 23 9E
 66 4D 49 CB 2B F9 28 54 34 94 D6 15 6A 37 E3 00
 06 CE 8F F0 B0 B2 3A D0 3B 0B 10 6E 68 46 8B C3
 98 0D BF A6 AB 97 41 53 EA 6C C8 64 B3 20 EC 9F
 A5 EE 9C 48 C9 7E 91 EF 80 82 23 7A AB 02 37 E8
 FC 15 2F E5 14 A2 0E 57 2A 20 18 1A 4D FE 3F 49
 0F 2A 6E F1 CF 8E 85 23 78 D4 CF 78 EC FF C8 8B
 07 66 CC F4 DD 9B FA 51 34 4F 6E F7 DB B4 B5 62
 8F E6 08 E1 20 97 01 59 74 A9 12 F6 EB 8C 8B 40
 8E E0 57 45 B8 9F 80 5B 59 71 03 BF 76 D0 CA 9C
 5D 0F 61 77 F5 93 1D 26 57 31 77 86 19 CF 19 41
 AC 8F D5 CA EF 8D 48 2E 62 12 34 0A BF A8 8B 2C
 42 A6 1C 69 3D 7E 94 77 2E 17 75 10 59 F4 2D 54
 36 54 15 89 E0 FE FC 81 3E CF B5 8A 6A 3D 60 F7
 B8 5A 67 8E 68 49 7C A8 D1 AC 00 85 92 C3 6F E9
 0E C0 39 1E A9 9A AD 89 2A 34 3F 2D 36 FB 95 50
 6C 3C 40 62 E3 29 AA 66 03 1E 0F 0E 1E 16 AC 61
 0A E4 A3 4C 2B AE 3B 40 E3 57 C0 0F 3C 8B B4 85
 5A 6E D0 0F 61 80 82 71 D7 E2 9D 34 87 CF F8 67
 7C 3A 1F 2B EC E4 36 5A D9 D0 86 E3 B5 42 25 99
 1A 57 32 E8 E4 8B CF CC F6 EF CE 13 F3 7D A9 51
 E8 BB 79 FE F5 5A 70 F2 C7 5F 47 CE 3F D0 BD 2D
 42 42 D3 52 8A E9 DD 75 CE 8A 7C 09 F1 68 DB 5E
 75 40 9D 9C 5B 9B A5 BB 7C 12 B0 16 31 43 40 EB
 77 06 E1 75 D6 D2 CB 16 37 89 E5 95 02 E8 62 01
 97 34 4F 2E 47 3B 12 1B D4 A1 47 94 A1 6C 52 E0
 39 B4 8A 54 76 AE 00 10 DD 3A F0 AC 28 9D B7 25
 BB C1 8E 7C C8 9F 58 AD 55 DE 45 94 42 40 59 56
 70 E7 0C 0A 36 D8 2A F5 0E 2C 25 47 87 6D DB AA
 AA 94 27 D3 9A B0 19 58 55 73 1D 67 9D 58 64 16
 B9 91 9D A9 5B EB 37 DF F3 F2 AA E2 12 65 08 27
 FC C0 14 DD 7E 3A D5 77 D6 9A 23 4E B6 84 D8 9F
 A2 53 41 82 8D D1 E7 30 24 EB 6B 1F 38 46 53 21
 F4 BD C0 EC 6A 5A 28 A9 F5 D5 E5 B1 AE 10 99 C1
 9D C7 EE E0 60 9F 9F C4 C7 98 ED 9B FA 63 13 73
 F7 7C DC A3 35 87 FB 48 9A 54 CE 30 83 30 3A A7
 2E 77 2F 3E 89 0C F7 A5 C2 69 49 4B 09 DD 9D 3A
 3A 7F 98 60 85 03 88 87 33 18 F2 76 54 63 24 1C
 85 99 5F 8B C2 C5 B6 EC 92 56 3E 0E 0E 57 35 40
 DD B9 34 56 44 F6 DE 4E DB EE F6 4D AF 24 0F 51
 89 E2 75 03 38 CB E3 F5 B4 48 2F B4 F2 81 C4 17
 59 6D 6A BC D5 F8 C1 EB B1 D5 3D 47 93 9F E6 92
 CC E8 0F C4 4B 5D 4B CD 07 FD C1 76 17 82 6E 5F
 86 27 CB F7 52 38 36 F1 8F B0 59 41 1A 25 EB 2C
 0F 44 0F 75 B0 6A A0 5F A5 03 0E 88 A9 FC BE 47
 E1 27 DD 14 EA 3A 08 34 81 9D 25 B1 63 D7 D9 1C
 08 93 F5 77 D5 A3 0F 69 50 FA 81 EA 32 E8 5B 45
 85 C6 04 C2 0B C4 36 B8 EA 3D 63 DE F7 EE 53 83
 4A D2 B9 93 D0 0A E3 9A 5E 94 12 79 30 8D 7D B3
 4D 50 BB 64 70 08 28 0A 29 82 C8 03 36 7D 2F 0F
 9F 75 A3 F8 6C C4 9F 84 E1 D8 E7 0A A0 C9 83 D0
 1C 0F DE 84 30 EE 83 A0 B2 94 D8 0E 60 EB 32 B6
 F5 D4 4F 5B BD CC 1D 10 79 2C 84 4A 0E C0 B3 06
 CD 7A 4C 78 81 B7 BC F6 1F 11 FF 2A C0 B6 85 10
 3F 8D 14 5F CC C6 40 1A B4 A3 35 36 76 22 C2 8B
 65 17 08 9C D5 92 B6 F8 46 40 C5 A3 82 ED 1F CC
 52 44 A5 15 88 1B BC 62 5C 1E 2D A4 4A 3A EE BF
 89 2B C2 13 5E 17 B4 EF 83 7C D5 4A 7D 1B AB C8
 67 5F F3 5F 0A E9 C8 81 42 C2 7E 1E 5D 49 BE DB
 E8 74 2B 16 C3 A0 51 E1 CB 9A 7F 44 61 46 A2 9F
 8F 69 13 1C 06 8D DB 7E 59 83 F1 BB 73 81 62 1D
 96 A0 29 0F 86 3D 9E 01 53 EF 56 4B 99 9D 06 48
 44 A9 9E A9 58 EE EC F6 B1 82 DC 11 31 9C D1 1C
 8A 7F 07 90 8E CE 87 8F 2F FD 51 07 E1 41 F9 B6
 83 CD 36 2B 9D 72 2D E6 EB C7 B6 A8 0E 18 FA 66
 73 40 1F F7 2C 2E 48 CE B5 21 77 83 8D 31 87 AD
 03 7A 50 B7 00 8C 70 50 3D 31 8C B4 4B 7F 09 B2
 2E 35 14 A9 2B 69 69 86 AA 6D 4D 91 C8 BC BD C0
 A2 E7 0B A8 95 8A FC A3 E6 8E D5 D1 25 EB A7 0F
 55 F7 78 CF A6 34 63 92 24 26 DD 16 37 ED 5D 17
 7D 24 FB 55 87 43 81 7B 22 DA 5D EC 92 BD 0C 0F
 CF C6 01 DF FC F3 6B 4F 80 10 BF 7A BC 57 BC 57
 52 7E 92 4F E3 DF 24 C4 D5 29 51 7A AE 34 3A 6D
 D2 E9 60 72 F6 97 92 8A 4E 38 2B 39 CB 23 1D 94
 C5 7E ED DA 0A CE BE 82 0E 47 3B 9F 07 0A 7B 6D
 F2 B7 BA 74 F3 31 91 F8 FE D0 24 55 67 D9 D1 5D
 1E A6 43 A3 26 74 71 D3 FA 40 2E 7C 9F EA 97 34
 68 14 6C C2 0B C1 B9 C4 1B B1 5E 1C A4 A8 06 2C
 20 CB 8F 41 62 2E A9 4E F7 6E 12 AA C2 6B 25 23
 34 02 4A 8B 5B 17 0C B8 A5 B7 11 6C EF 10 DC B6
 A5 A0 E6 86 E2 A0 B7 99 ED 18 80 78 BF B9 9D 6E
 BC 5E 81 F8 55 FF 00 F3 03 A9 23 BF 0E E3 D9 CC
 53 71 20 CB F7 2D 21 54 E1 1F BF 93 27 E4 41 2F
 E1 AB 34 78 B7 F2 42 8B B9 F0 DC EE 71 BF 88 83
 A9 EF 43 32 1F 9C 2E 70 59 90 0F D7 8E 9A D6 5E
 E0 1C 31 61 FA 18 3B F6 CB 4F B5 F8 64 62 95 72
 81 B7 A7 12 DD B7 29 E1 7F 88 0D 55 6C C1 84 A5
 0C 17 57 40 6B 19 11 DD B1 19 04 3D E5 8F 11 80
 73 E7 85 00 88 99 48 23 AC 8A 1F F8 F0 07 54 C3
 1D A0 94 64 BB 47 3D 47 BD 77 31 B1 C6 89 CF BB
 0E F7 10 E2 D8 2B 45 F6 40 59 CE 8D 05 E0 D3 19
 37 56 7D 37 45 85 9D 4D 4B BF 06 E2 88 DD B1 A3
 1D D2 0D 48 C5 FC 8E 70 FA CC 41 DD AB C6 E3 BE
 3D E5 05 7A 23 1B 96 4A 17 E3 0A AE AD 95 93 B3
 3A 05 74 31 DE D7 51 0F EB E3 56 7B 08 E8 AD C3
 B1 87 6E C5 58 76 94 DF 44 0E 20 15 72 B9 C5 25
 80 04 84 CD FA E2 82 13 17 91 61 7E 63 0E 32 D5
 09 B1 AC 2A B8 11 95 90 DF E9 77 68 EC C1 8B E5
 E7 A2 3C FB 52 8F A1 DD F4 D1 F8 95 13 B2 FF 01
 74 5C F9 50 55 9F 37 B1 E4 EF 07 AA B2 5F 81 61
 AA ED 88 04 CA 20 2D BF 4F A7 B0 8D 50 35 FA 92
 D3 57 E9 19 2E C3 E2 D0 75 31 F3 03 59 E8 44 25
 E3 F2 E2 04 FE 85 A8 41 EB 00 E3 84 56 CF E1 D3
 A1 B4 D4 13 66 19 8B 46 E7 C8 BA B1 B8 3E 2A B9
 EC 2E 05 44 66 CF 8B 5C 3D 2B 79 B9 D8 E9 45 24
 67 20 55 21 D2 36 C6 C3 75 02 C8 E4 CC 80 61 B4
 3F 8A BF 01 DD 60 C1 44 8F 10 10 33 FE 6F 18 B6
 7B 60 4B 7A 98 EB 39 0D 9A 95 DC 13 31 69 C8 00
 6B 16 52 05 5F C6 77 B7 FA D6 E7 A6 8F A4 38 11
 74 23 99 96 11 D7 DA BD 03 50 16 D3 08 17 B8 CD
 98 6C B9 78 65 5F 3B 5A DA E5 92 DC AE 83 49 83
 19 DB 39 E1 D6 47 EB 24 71 CA A9 9F 10 0A 2D A9
 1F 45 59 96 65 D3 11 6A 28 E3 0E F6 26 90 18 EA
 02 47 88 87 78 6E EB 53 65 36 E2 E7 D4 21 AC BA
 D9 13 8E B9 78 00 8A E8 20 9D 6F 3B 9C DA EC F7
 AE 21 78 37 DF 91 9B BF 1C 4B 8F 9A 40 D5 E8 15
 49 83 EC 47 71 2A 74 23 A9 DE 2B 08 9C 91 CE 19
 81 E2 3E 56 7E 76 22 FC 62 A7 3D 00 09 94 21 4F
 68 CF B7 FE 1D 17 03 55 F6 E2 D3 D2 76 03 AD 4B
 9B 21 06 8F EE 91 7A 87 DD 4D 73 C8 D6 91 67 E2
 C1 75 C3 1D C8 9C A9 E5 B1 6B BD DB 9B 36 21 7F
 CB 6E 97 68 59 AC 76 C2 78 B5 53 7B ED 62 F9 A8
 53 49 4D EE 34 3F FE D3 6C 37 26 6E 9B BF C6 A1
 E6 D8 B8 C2 F8 99 90 43 6B AD DD F4 45 A0 7B DA
 9B 19 90 92 1E 58 54 25 D3 E6 4E 00 C3 FB 80 28
 B8 CE 73 46 A4 68 AD B2 B9 35 FE 16 90 1E 4E 0B
 E4 08 35 25 BE 6D B6 06 9A AE 61 94 69 AC 3A 9E
 25 DC A1 DD 69 C3 8E B3 48 37 65 F2 09 7E C5 83
 3D 8D C1 55 2B C7 53 A9 EB 7E 21 D0 FC F2 8A 29
 3A 0E AD D4 06 EF 8B 51 61 AC 50 10 CA 72 B0 C1
 57 38 D4 45 62 F3 EA 26 63 51 63 3E 80 8B 28 96
 91 BF 02 42 A8 0F 04 90 9D EF 05 BC F0 00 B3 6C
 80 48 3F 1A 70 B8 E3 D2 98 08 02 E8 40 62 F7 CC
 A0 F3 B2 E6 B6 3D 22 0D FB FD E6 64 E1 62 D1 D0
 F9 A3 94 F2 7E A2 CC 16 75 99 FD 42 C4 08 4D DC
 81 06 FF 5D DE 07 80 33 15 6C 99 A9 B1 9F 7E 34
 86 B2 AE 37 D6 3E 59 1E 76 3A 5B 42 65 41 AD 61
 E1 A8 1F 5B 74 9D A5 FE BE C9 53 98 F9 2E C1 93
 73 15 29 62 BE 72 A9 43 E1 03 80 CA 59 CC 70 13
 BB CC 9D E8 42 84 5F 8A C2 8E F1 A3 7E D9 3E 23
 D6 EC 4F 86 37 20 46 4D E4 5F 78 3A CC F5 8B 62
 FE 40 54 9F 22 64 3A 33 03 4A C4 E0 B2 04 EC 45
 57 CF 5F F8 CD EA A3 CB 23 7A E5 17 66 E1 44 0B
 98 AE D0 85 36 3D 4C 27 9F 17 4D 75 E8 0B 96 31
 98 5A F1 97 D1 4B 72 67 00 E4 FA EF 58 CA 7C 5A
 7A 41 EA 3E B2 42 10 50 CF 65 C8 15 DD E3 97 88
 4F 76 F6 71 B6 9C BB B9 74 00 B7 95 25 71 73 58
 13 23 7D B1 7E 0D 75 E3 A8 FC 0C 44 DC B7 75 80
 DD 95 F7 C8 5E 6A BC 23 BF 8F F3 A0 30 CC EE 87
 AA 78 AF 85 F4 72 64 DB 8A E9 27 1B FE 1F F0 17
 57 81 3A D5 8F 48 6D 25 72 E1 9D 9C 19 75 13 EA
 1A BC B8 ED 79 87 CC B1 55 CD 00 FA E5 05 43 CD
 20 6E C7 E0 04 40 9D 00 83 E3 32 42 D6 E5 D7 9F
 6C 5B 62 35 21 40 0B 51 1B CA ED 63 38 BE D9 5E
 97 85 11 56 76 9E 05 AC 21 16 37 61 E7 24 F3 D5
 BF 25 02 BE 11 1E 87 CC A1 04 22 8A DB 58 FE 6D
 DE 6C 84 25 20 8E 14 90 6E 03 96 3F 4E 49 A2 14
 5B 05 37 66 A7 D3 7F B0 D3 75 AF C9 07 98 48 85
 07 8D C5 3B 6F 3D D0 FC 40 7A 8C 38 E1 D9 79 7A
 2F 08 D9 46 A0 25 F7 B8 07 D9 78 A2 FB E7 E6 70
 EC C4 18 C4 29 92 58 25 86 2D 10 31 97 01 DB B4
 11 43 1E 77 57 C2 59 AB 85 70 9B B3 16 59 51 58
 05 A1 48 62 CA DB 83 F5 5E 2E AE FE 5F 03 4A 09
 D8 F5 DA C1 43 B2 A2 22 0A 89 55 33 D3 4B B9 15
 08 7D 0C 8C FF 65 96 0B 40 67 42 B4 3B 17 30 E2
 19 C6 3B 27 68 B7 AB 97 50 A1 2E FB D4 15 88 1A
 D0 84 B0 9D 11 01 5D 4C D1 89 F7 05 64 08 DE 5A
 B5 FD FB 1F 06 A5 BA AC F8 A5 CE 62 E0 83 BD 2A
 D4 64 A2 9B C0 35 4D 66 7A E2 E5 74 AE 2A C1 DC
 F0 67 16 F4 DE B8 01 70 12 E5 0A 4A 0C 67 28 4D
 9C 4F CA 5B AC 13 18 9D 90 51 C8 9B B3 A0 7D 14
 5C E2 42 F8 38 C0 A1 2F 28 40 3D 20 A1 80 2C 9D
 B5 25 7F 98 7A 1C CD 35 DA 47 6E 76 6F 98 7B 91
 4A 19 9C 3F EF 3D B6 80 F6 7D 3E 1D 1C 22 92 C3
 65 00 C6 EB F3 EE 8A 7D FE 6B 9C 85 53 49 69 A5
 67 EE E3 0C 39 59 A4 A7 D2 19 52 18 BD 1C 02 5B
 93 5F A5 5B 4F 0A DB 21 F5 4E C8 43 74 BD A8 DC
 96 13 81 4B FE 0B 21 2B 80 4B 6F F5 74 9C E4 D4
 A8 C5 79 F9 C2 A2 CD 3E 41 C8 B4 96 A4 2B 76 E3
 71 99 B5 F5 56 2D 24 15 1F F2 90 53 C7 EE 34 BD
 F2 B6 7B 8F 51 11 33 E9 33 C9 86 5C 51 86 0F 1B
 E1 CA E6 B0 A0 51 E9 20 FA 6B C7 4C C4 A4 83 42
 D4 A9 72 5B 35 53 32 55 F9 06 3F 84 27 F1 28 E3
 D7 F5 A6 5C 1B B1 25 50 0A 5B 3C 8E 1D F2 96 6A
 CF 18 DE E7 1E 89 C8 87 3C DC A9 C5 AA 80 AB 8F
 EB AC 99 D7 81 36 DA C9 7D DA FA 29 C1 A2 9A 6F
 CD CB 0D 08 8B 3E 9A 2E 4B 26 2F 78 D8 23 A2 53
 B4 A0 F6 21 CA 29 C0 68 E1 24 7B BD AB 7B 79 4C
 A4 E1 D8 09 7B 28 88 B4 3E A0 E5 0C 50 07 39 39
 90 1C EE 2F ED 71 A6 31 1D E5 10 6E A3 A8 90 52
 E9 0A 90 43 20 52 7F 3D 21 32 FA BB E1 67 17 FF
 33 15 0B 52 D4 D9 94 20 CB A1 F0 9B 71 18 04 2F
 B6 0A A3 FC 4F F4 42 C3 25 5C A6 A7 E7 FD A2 22
 8B 16 61 29 24 86 5B B5 CC CC 09 BF 25 3D A2 59
 B9 C2 05 CE C2 68 3F 00 2B 26 09 61 78 19 75 0B
 63 85 3B 44 87 77 91 A9 F4 6F 31 80 84 E4 E2 FC
 FD 8C 69 63 B9 4A 0D 20 F0 C4 15 0B 1B C1 F8 BB
 6C 3D 12 09 07 E2 04 9C 1F 3D A4 96 F7 F4 E1 FD
 EA C3 8E D0 A3 E7 77 6A 69 EA 0C 38 1F 89 0A 3D
 1A 9A 56 82 C9 8D 70 76 21 6B 4F 8F A7 45 C6 B2
 B2 F5 7E 80 2B FC A4 3C 53 BD FC 83 81 CE 94 5D
 E0 A7 9A D4 E0 49 67 EF C7 E2 2E 9E 51 65 6C 8A
 26 2A D8 38 6B 5B 81 0F AB C0 D9 ED D1 6F F9 86
 55 A3 FF 7B DC 72 07 CF E3 C3 69 83 58 B1 9D 56
 17 BF C9 C1 50 19 7B A5 B3 DD 28 00 DB 0F 7B 92
 84 68 34 13 49 C3 88 A0 EB E7 77 92 17 A9 AA 60
 B2 56 33 8A 35 ED C9 BF B6 BE C3 18 F1 AD 4A 2A
 E7 AC 3A 4F D1 33 71 40 B9 57 48 03 BE 78 A9 0D
 AB FB FC 6D FE 39 E4 91 B6 31 65 AD 48 71 02 92
 F8 8D 47 AC BA 99 CB A6 E9 C4 8B 54 56 8F F4 D9
 A5 FD A5 13 FE D3 DA 74 02 29 A9 0E C4 0C BE C7
 41 D3 CF DA 09 38 DF EB ED E2 58 41 2F AB 19 3E
 35 4D 9F 26 BF 60 79 25 C5 27 DE 6F CE 20 2B 38
 71 32 D6 09 9D 76 C1 58 28 0A D8 25 96 BC 39 D9
 26 10 50 6C 2A 49 E3 0A 8D ED E6 61 EE C3 5E 8E
 C9 1F 37 CA CB 0F A0 2D C2 80 E2 4D 99 C1 9C 9E
 13 A3 13 A0 48 02 23 5C 98 83 BB E5 9D 67 BD 71
 CC F4 03 98 B7 2E 6F CF 03 A5 37 71 FC 27 11 4A
 14 9B 3D 59 02 4E B0 30 9F 59 F9 75 67 E4 DA D5
 AD D9 12 69 CB 07 66 74 24 BE 18 1D 21 B6 B6 49
 35 DB 8C 76 33 E6 41 7B F7 AF 7F 74 45 C0 DA BA
 A4 83 70 D0 BB C7 2E F3 3E C1 1E D8 4E E1 8E 46
 BC 38 70 05 8E 69 C4 29 22 7C 75 FF 69 EE 86 A6
 DB D0 BB B6 E3 09 87 42 AA 64 68 20 68 E7 A6 BE
 17 62 B6 57 5B 7A 14 21 0B 59 AD 0E D7 76 58 28
 24 25 C9 C2 B1 25 B0 42 8A A9 1E 42 B4 63 65 EF
 59 30 F0 DB CF 8F C5 6D 33 E7 6A 8C 5A 4E 5D B6
 1E 63 B8 8A 99 72 5C FC 74 7B 2D C4 26 0F 0E D4
 E5 8B 7A C4 A8 FC 2B B5 40 82 D8 BF B4 D4 DE 27
 96 11 35 F1 06 A6 56 E8 72 45 0B 80 F4 26 08 5F
 96 ED 42 C8 EC 0D 9E 8C 9B C8 0D 66 0F C2 1B 36
 61 09 6C 86 EB C4 66 7F 27 4F C4 3D 28 9E 56 70
 12 03 4E BF 2B 39 8C 8D 64 3C 7A BE 42 67 B0 40
 A8 70 B3 A6 0B 9B 6E 05 C3 AC 47 2B C1 BC 29 44
 F0 8E 4D 7D 55 28 D9 81 5B 60 A9 5E 0B 02 E0 C8
 DC 61 E4 3C E2 FC C1 04 7F DC E5 6B 37 18 CD D0
 70 D4 2A 3E 31 7A BB D1 4D 70 C0 E5 1C B9 50 52
 E1 0D 46 14 E1 AA 02 6A B3 67 57 24 0F 41 0E BA
 BC B1 8B E3 6D F8 AA 1B BC FC 1C 37 57 E8 FD A0
 B8 91 86 0D 93 66 BD 97 E2 64 64 50 A8 2F 8B 98
 3A E1 94 D5 B8 78 D7 CF 37 66 E4 C2 B5 B4 95 98
 E4 B5 02 41 24 46 CB 82 25 09 28 B5 9E 8B 98 33
 B8 56 15 89 09 9F 85 70 4C DE A7 2E 59 5D 55 99
 4B BC EB 7B 01 96 53 A3 C3 2B 46 06 5E 59 78 89
 4C D2 D9 7E 6C 66 D5 62 2C 85 83 B8 93 03 9E 15
 1C E8 B1 C7 D4 FB 10 6A 43 48 5B 9A 2A D9 28 F1
 53 C8 1A 1F F3 AF A9 65 F4 1B 9B 7E 5A 2B A0 9D
 B1 50 59 A9 09 5A 88 48 36 A9 3A 8B EE 59 4C 1E
 8F AF 1F 43 4B E2 D8 82 89 84 64 54 B0 6B 21 FE
 5A C6 1D 03 92 B5 48 3B 72 03 E0 1D B4 4B 9D 9B
 70 05 4D AA 02 D9 1E 52 68 40 FC 2F FA 28 EB 1E
 79 B7 F4 B7 F6 CD 90 80 A8 E0 4C BF FD 4B 7D 64
 29 CF 07 80 5F 76 21 0E 6C B8 AE 11 18 3A 06 E1
 4D 89 BC 87 C5 8C 96 9F C7 D0 33 62 5A D2 82 03
 3C 35 2C 2E 5E 41 13 02 10 30 8D F8 76 3A 83 9E
 08 00 4C 6E C9 BD F6 DD E1 BC 3F 3E 3E 98 70 E5
 97 B7 13 5D F1 A8 12 F2 20 2B 63 CE A7 55 05 FE
 24 F6 25 48 D7 A5 0E B1 19 82 E0 BF 90 9F FF 51
 07 E4 C4 5C A5 00 9C 16 45 CB BF 72 3E BF 6A A1
 0A 90 18 4A 36 09 0E 47 F0 EA C2 AE 6E 60 25 3D
 B2 82 AB 4B 20 E5 4F 73 91 85 92 5A D6 B5 06 4C
 BA E4 4E 5C 30 EF 98 E2 8D 14 B0 2A C0 EE 2A 1D
 37 F5 50 B2 77 25 09 E2 A9 28 41 82 77 F2 B1 76
 47 BF 35 FC 7B A2 1F C2 23 76 31 45 03 A1 2F 7E
 2E 5E 68 6C 46 9A 47 15 1C 88 60 DD DD F1 4A 75
 20 2D 94 FA 69 FA 65 9F 23 93 8C 81 69 97 3B EF
 60 BA 5D EB 34 63 E1 C6 4F EA 8A 5C 4C BE 21 92
 DA A9 69 42 FF D3 42 32 FD 84 B6 53 E7 BD 1D 5E
 AC BB B3 13 8E 3B 26 D3 64 75 0E 4F 4C DB 33 E3
 DC DF BF D5 D8 87 46 0E AC CB FD F1 FD 1F 57 D0
 A5 04 85 79 D8 11 ED FD EF E2 74 1D A6 CC 3D 05
 AD 94 73 B1 6A 11 56 46 5F 07 9B D0 3E 34 4C B9
 1E AB 96 72 D9 84 B5 20 3F EF 2A B4 2C 80 25 A0
 F1 F9 04 A1 91 8B D1 A9 50 22 48 A4 12 ED 5C 1E
 76 CB 9C 77 46 87 BB 61 78 25 46 1F F8 27 6F 5C
 47 D8 F4 83 C4 72 98 AA 52 9C 61 12 F6 B7 16 2F
 F8 F0 5E 92 39 01 4A 11 36 4F C1 17 CB C5 A4 78
 9F DF B9 AF EE 7D AC BA 61 AC 71 1C 72 95 F5 93
 D1 D7 6A D8 6C A8 5C 42 49 3C 52 6E 4C 08 3A 7C
 44 B4 8B C1 FD 48 7D 2B 90 B0 79 7D BE 0B BE FE
 81 F1 35 D6 70 42 E4 FE 3E 97 7D 8E 54 7D 8A 4F
 B2 00 94 DA 00 AF 0A 05 19 53 6C 8D 3F 17 73 8C
 F9 62 24 B1 50 9F 5B 6F 42 D1 AF 06 47 F5 26 E4
 66 31 60 26 74 AC 7B F5 E6 84 DD F2 08 B8 61 17
 E3 01 91 46 54 84 0C 9D 66 0B 1D 13 7C E5 B9 56
 DB A7 26 29 F1 98 62 DF 1F AD 8E D0 1D BE 3F 92
 5D A4 25 00 0E 58 10 37 DC 63 3E B6 AD 9A D0 83
 03 BB 16 CF 5D B8 C4 3C 31 13 37 2F F8 12 05 41
 90 8E 53 34 52 11 D5 26 69 FD 5D 8D 63 40 0C CC
 B4 FD 56 54 2F BA 09 41 42 11 EC BE 44 A7 54 70
 D6 E6 29 4B 7F 2F D2 AB E7 B7 76 1A 43 3F 77 96
 CC 54 F6 5E 28 B3 49 B6 E0 92 68 1D EE BD 47 59
 05 17 35 E6 8F E5 2A A9 60 B0 F7 80 74 39 35 08
 48 02 5F C1 22 80 6E 78 91 F8 EA 21 74 35 CB 49
 8F 06 DC 2D 1F F1 1B 99 D7 D0 16 A9 F3 EA B6 96
 7A CA CE 66 00 38 53 4A D2 CF 2E 7E 6B 13 10 16
 0A 5D D1 E1 39 BE D5 BD A2 B6 9D 40 F0 99 D0 F5
 AB 56 28 85 75 7A 42 60 30 2D 3C 5F CE EB 1C 16
 0E 6A DA E5 F5 CD AE 34 B7 26 0F 76 82 91 32 56
 AA 61 10 B8 6E 5C 99 87 60 12 C3 88 DF 15 65 A2
 39 BD E5 B2 1F E8 89 A5 DC 97 19 E5 AC 82 0B C5
 74 8E 4C D1 BC 0B E4 2A FB ED 6A C1 A2 3E E6 BB
 8E 47 52 BC 92 DA 71 6A C6 C7 79 99 F2 AF E3 16
 CD D7 2A 08 D3 D3 77 19 A9 FE 8A FD FD BC 7C 53
 8C 05 94 CA 8A C6 E2 21 A9 9B 7E D2 F2 15 D7 E0
 F2 04 EE B8 DC C3 39 9C B7 EE 35 FB ED E5 E2 54
 4A F2 A6 7C 5E E9 48 50 34 12 7D 85 79 33 C5 5B
 6A D0 7C 24 F0 AF E8 EC E9 AA 53 89 40 E4 19 B8
 39 B7 91 21 53 B4 8B F9 77 A8 17 4B 25 21 FF C3
 D3 22 A4 67 F2 8A 92 73 2C 0D 9B 9D 72 18 1B 7D
 D3 E7 B2 3D 62 9F 59 28 C4 11 D3 EF 13 67 E6 F1
 56 85 FF 2F 24 DD E0 1C 23 74 7D D3 35 F9 58 38
 54 47 83 BE 96 10 FB 69 14 5C 89 2F 6A F7 38 C2
 B4 14 18 95 76 56 4F 1E DF 1E 47 30 87 0E B0 BF
 0C 17 D6 BB CB 4C 7A 3F AB FA 31 85 79 DB 52 38
 45 DA BD 55 F0 CA 4E FF 2E 67 AB 8E BE 4A E9 F6
 FE 36 A5 CD F3 4E BE 69 10 E7 55 55 B4 9E 3C 49
 4A 38 C0 B9 C0 CE 73 BA 61 4B 0A E8 6A E4 83 6F
 9F 19 B9 3B E5 1E 78 C9 9E 8A 0B 86 10 3D 15 0A
 AA 8D F0 7F 3A F7 AC CA 0E D8 E5 61 A1 65 F1 A2
 B1 C6 CE 7A 64 38 6E F9 F5 DC 2F 97 ED B8 39 7E
 4F 0C D8 AE 70 5B D5 F2 19 D9 CB 9C 7A EF F8 18
 C2 20 C2 24 4D 69 ED 6D 3F 81 3F 86 64 88 5B A7
 07 FB 80 2F 83 4A 40 0C C7 CD E9 61 E5 C3 65 B9
 C6 75 74 51 56 C5 F4 2E CB 1D 06 30 5A 1F 80 B5
 53 10 8B 1E F0 D4 C9 3B 3E E6 4B 08 46 7F BF 6A
 B2 01 9B D7 87 3B B1 A9 3D 05 B5 1C 70 29 92 22
 EF 6D EE F5 C6 CF 23 61 99 D7 D8 0A 76 B3 57 5C
 CA CC 41 96 92 BE 1B 8C 14 08 9B 3B 7D A4 62 3A
 48 D7 F4 3B 06 80 37 CF 34 E6 3F B1 C1 2E 78 5A
 57 DF F9 A1 53 71 42 5A 5F 6C DE A0 AE FA 3D 82
 25 80 39 3E 9E 12 CF E7 EE 2E BB 8F 19 11 6F 78
 7D 5D 96 6D 1A 76 C9 03 DF 18 F1 0A 5C 29 8D 0D
 60 81 BD 46 CE 5C 3A 3C FB 0F C1 FA 82 6E 8D 0C
 01 52 01 9A 58 11 94 CC 0A 85 83 29 56 98 AD 70
 64 32 5E C9 B5 40 27 00 22 85 E7 65 84 83 0B 4C
 EE 64 9A 4D BE 63 3E 88 50 18 89 02 C0 47 DA 35
 69 A5 7D FB 98 8C 10 42 1D 1A 42 F4 F6 4D 9E A5
 B9 34 EB 8D FC 7B 3B 6B 23 36 79 54 3A C8 A7 6B
 5C FA 41 39 E2 9B 70 EB 53 E7 E9 A2 B3 B8 B9 32
 F8 1E 75 F2 41 D2 3D 24 E1 C2 F8 E4 91 3C C6 D6
 34 99 3A AF AD D2 80 CA AB 65 EA 8C 21 02 35 24
 8E 53 F0 FB E2 16 93 84 CB 6F A8 A6 D2 85 11 D5
 7A 8E 11 DF 1D 2A FC AC 97 27 C0 1C 02 3A 6B 76
 78 41 24 7A 5D 97 7E 5E D1 14 1E 7A 36 D0 13 3E
 94 E8 35 0D B4 8E A2 6D D3 7D 4F 6F 87 79 3D 1C
 3E F4 00 BB E5 20 D9 6F CC CB 50 22 07 CA 25 C6
 AC 17 21 FC D7 A6 47 BC A1 8D EA 82 14 78 6F 51
 4C B3 EE BD CE 41 34 F5 53 D3 F6 96 B0 D0 91 C3
 D4 CB 0A 1A AC 6B EA 99 EC B6 F7 2A F9 9C 8C E4
 F5 23 B8 F1 8D 57 C0 43 41 31 DB 7C 17 AB 88 9F
 A1 0B B0 AB AE 6E 2B 97 36 C6 5D 2A BE 72 43 17
 4E 73 C5 EC 02 1E FA 2B EE B2 AE 15 EE 65 1B DE
 F0 8F 2D 4B 61 1E 72 F7 F3 98 1D FA 05 7B E3 77
 C7 12 DB 93 02 77 C5 A1 59 7A DB 88 27 96 4C A9
 1C 5B 81 73 A2 CB BE 97 D2 ED 55 E3 C2 6D 3D AA
 A8 EA 23 F9 06 C8 29 D6 48 E9 D2 4D 5F 96 5E D3
 EE 97 02 C0 1F 60 D2 85 5E 7D AC 2A 05 BD 01 A8
 CC B3 C4 1A 30 AD 75 CA D7 8C FA A7 78 25 15 6B
 BA CF A0 F5 39 B6 3F 2A E1 5F 9D FD 34 12 2B 6A
 E1 29 56 35 D8 20 C3 44 A2 56 C5 81 80 17 09 3C
 AF 26 01 56 DF 6A 58 6D 12 06 E6 39 9A 7D 88 3D
 64 FC 0B 53 F8 84 20 8B 74 E9 5C EB 53 EA A7 63
 CE D4 B9 23 98 5E B1 7C 58 44 10 C4 29 D3 95 1C
 A1 AE 76 75 93 B1 5E 2C 4C 2D EB 5C C9 08 74 6A
 67 BD 72 53 9A BC 99 16 37 27 48 EE 09 52 DA CF
 D5 2D A0 0E 14 4B 0C 24 B9 54 BB 3B EA 1F 22 37
 15 F3 F5 82 87 E4 F1 4B 64 18 AB B3 59 EE 03 78
 C7 0F DB 03 27 EC 03 12 7E 2D 3C 13 41 F0 44 B1
 BB B9 72 A8 EF 23 CE 1E ED 82 A6 92 0F 33 C6 17
 0F DB 33 C2 AD A1 BA 01 E6 A2 7A E7 58 3F 2C 51
 80 77 DD 62 BD FC 85 B6 13 BF B4 F8 14 9A E5 55
 44 91 3F 9F FF 1D 86 35 49 64 83 54 08 20 40 66
 6A B3 40 70 5E F6 C2 14 FB 78 5C 21 B0 AB AD AC
 00 B7 9B 25 99 F5 5E 3B FD D7 82 16 19 A4 37 8D
 80 91 F7 3E 47 A6 98 80 9F 41 79 24 94 03 9E 99
 CE AA 8C 48 20 8D 73 BB 0E B2 63 17 C2 6C 96 75
 42 66 75 A1 95 B4 AB 30 EE 75 FF 0B 75 4E 6D 9F
 A5 B5 3F 7E 91 D4 48 7B 7F 01 8D 32 20 4C 51 60
 1C 79 BA 55 7F FC B2 9C 9E AD 28 0A 8D 88 60 30
 E0 86 4A A5 A7 50 7F 3A 65 EC D0 C1 8E 78 E4 D2
 5F 65 1B CC DB 10 77 6C 2D 2A 8A 0B BC C9 EC FD
 F4 FF FA 62 1F 99 63 22 4D B6 30 8D 50 72 6E CC
 4C 0B CC 62 6D A0 5F C8 9C 92 61 4F 6A B1 9F E1
 39 A7 FF 77 0E 9D 65 19 39 85 3E DB 7F F0 96 47
 00 AF 85 B3 02 FD 98 CA 16 91 E7 D4 FA CD C0 A0
 B7 38 74 F2 8F 76 A0 60 7A B6 D9 56 12 D1 2F A6
 D3 AB 3D 87 79 88 4E A7 BB 12 6A 23 37 B0 DD 6F
 2D 0B E2 C2 0F 82 32 9F 0F 64 F1 C3 C7 1C C8 3F
 DA 57 18 C3 0B 4C 03 F2 25 B1 0C 13 92 2D 77 97
 10 27 3D 6E 90 25 AC 78 AE 98 68 C8 9C 88 07 2F
 6A F2 03 66 45 E0 D0 42 C3 BF 97 8C F7 45 68 BF
 B6 B2 36 7B E7 13 49 26 BF 78 C7 04 37 8E 3A 7D
 88 85 4A 1D 7E 27 54 12 21 9C D7 FB 6F F3 99 F8
 31 58 4A 10 75 E7 35 C6 F0 9A 78 5B FD 74 F8 BE
 97 E0 5C 16 C8 3F 1B 69 72 A7 03 44 FE 6A C1 52
 67 D7 B9 4F 90 96 AD D9 60 CA 55 0A E4 ED 58 E3
 70 DD 9F E4 3E 47 41 C2 E6 34 C3 5D 85 8C 41 16
 02 31 22 F5 9C 24 81 34 01 E3 89 34 45 FD 2D F1
 9C ED E3 3D EC 8D 02 FB AD B3 D4 0F 44 AC 2D 3B
 E3 C1 98 05 16 41 2F F3 1B 56 93 58 FF 4D 20 50
 F2 83 CE B2 B0 06 B1 8F 80 F4 BD A6 BD 5A E4 69
 CC 68 06 95 61 6B 21 16 3D 21 99 70 EA 8F 25 0D
 68 56 33 1D 7E 46 BC 12 05 23 73 3B D2 7B 38 DB
 3E 90 69 4A EA 2A FB 5C 2D A9 BE 3C DB D4 66 67
 98 87 EB 67 E0 A9 DE 3F E4 25 10 73 D2 AE BF BF
 16 D3 B9 7C 9F 9A AE F9 F1 6F D9 6D 33 9C 36 1C
 10 74 0B C7 9F 32 56 3C 12 C6 5A 3B 11 4E 5C 5D
 A1 BD AD B0 B5 22 75 18 E0 51 0E 80 C8 E0 46 E8
 9D 79 BF F1 4F 77 00 D3 87 89 84 01 58 BA 84 AD
 68 3F 54 D5 D4 9E 44 BE C9 33 96 45 12 E8 CD 97
 7F EE BD D8 73 26 B1 A4 7E 91 81 D8 2A A8 CB 37
 32 B3 9F 0A 58 24 6F 0D 5D 5C 53 5E 7D 52 6A 56
 35 33 ED 6C 4D B3 3A DC AC 6F 94 B7 FB 5F 9E 32
 31 C7 14 8F 90 63 47 E3 4A A5 22 27 29 1E F5 52
 C9 C3 37 E5 0F 30 E1 A3 58 DA 16 85 C4 45 5D B6
 D1 FE 79 1B D4 F0 0B 9F 55 69 32 00 08 0E 2B 38
 A5 E8 77 25 53 1C F0 C5 6A 1E EC 78 A6 D0 E7 D2
 BE 3F ED D0 D9 E9 AA F7 71 DB 24 3F FF A6 B8 E8
 D2 5A C1 0E 1C 61 C4 63 17 8E B7 FC 75 BF 8D C3
 1D 78 45 26 82 65 B0 DE 52 54 DD AC 1D A7 48 70
 84 E8 24 D1 C7 8E 8D 67 A1 9B 26 B4 2B 24 A5 02
 23 4A 1A 65 BF E3 1E EB 7A FC 43 E7 79 C4 20 BB
 73 8F B7 32 4F E0 FC 4C 27 14 BF B6 E1 79 A8 38
 0C 43 F9 A8 2F 11 7D EA A5 35 BD 5C 48 F8 64 BC
 A7 E8 D3 2C 55 29 20 1B 77 A5 91 C1 4D 1A BC 92
 34 61 FD 2A E6 96 81 81 53 DD 4E 00 E2 3F CD B8
 54 FC AD 09 95 ED C8 D4 07 A9 DC 69 07 2C 6C 38
 08 8A BE DB 75 E3 F5 8A A7 6A 02 CA 6B 9F 87 E0
 EB A5 9A CE 29 4D 36 35 DE EE A1 F0 46 56 79 09
 0E 86 F6 9C B5 A8 13 03 97 0A AF 79 E4 25 87 6C
 B9 C5 0F 1F 41 A3 E7 D1 1A AF 97 DA EF 12 13 FC
 7E E0 39 2D FF EF A8 79 94 AE FC 0C 46 72 13 6F
 09 4D F9 75 45 ED 78 BB 7A 24 76 89 E3 1D B8 D7
 74 C9 C0 ED 38 C9 C4 D0 62 AA D7 F1 AB 0B 73 63
 25 3C A0 7D 6E B4 5F 1B CD 07 63 6B D2 3C 03 A4
 D0 42 A3 48 5E B4 88 FA ED D9 67 11 2C 13 76 9F
 D6 B5 EE 6D CA 43 24 58 52 CB 93 65 9A 6F BD 04
 83 F9 DF F4 C4 80 C6 51 08 F6 02 3C 61 EF 33 23
 BF 7F 52 4D 1F BD 68 90 A5 F9 2F 0D 9F 56 AB 5F
 B7 EE D7 FD 61 98 F4 66 0A 99 3E 16 8F 47 E5 02
 34 11 29 7C DC 73 AD F6 EF 87 F2 23 F4 59 6F 6B
 BC 73 D2 C6 9F 7D 7F 24 23 CD 2A 0E 5F F1 A9 D7
 F4 56 BA 36 2D 7C E3 FC 02 62 E6 1A 01 3C 39 A3
 7D 57 1B 14 87 55 9A 64 8B 22 C4 19 29 7A A8 A2
 DF B1 81 06 33 67 2B D3 F2 37 B8 AD B5 B5 51 AF
 C4 69 B0 92 9F BF 8A A7 08 11 3E 88 75 3A EC E5
 5C 49 6B B9 AE 5D 27 24 67 CA 23 16 73 63 ED F2
 62 6A AB 67 0F B0 12 68 BD 8A D6 31 DE FF 6A D3
 44 8C 40 0F BF 74 86 24 A8 39 49 C5 2C 48 40 DC
 F2 78 F2 C6 BD 43 10 9F 20 A2 3D D5 8E 6D AF CE
 9E 93 5D 31 89 54 1A 78 88 80 7F DB D3 48 67 0F
 F5 1D 21 5A 34 40 00 03 B5 EF A0 A0 22 AC E6 15
 40 5A C5 B7 32 52 9F E7 78 99 8E 67 A7 90 CF 86
 BF AF 08 6D 5A 90 0D CA 5C 50 80 A3 C3 D2 E3 CA
 B9 82 F2 D5 16 97 ED EE EF E0 BC 2E 68 78 1D 92
 58 A0 F1 5F F6 31 2B 02 64 90 16 BA 43 88 4A A6
 5F 81 F2 C8 33 8F 41 EA 1B 49 5D CD 86 C2 05 2F
 8C 17 5B 38 15 BF 9F 30 82 D8 6C 00 78 01 A8 B5
 40 7C 81 A7 21 93 51 32 17 E1 64 30 DA F3 24 ED
 A2 3F 73 5B 91 7D DA 24 41 80 05 08 A8 59 6B 59
 9D 41 AD BA 5D F1 9B 0C 11 35 CF 52 E6 0D 34 78
 DE 52 A9 A4 C5 1F D6 04 E5 AF 02 B3 6F BD 29 EE
 E7 C2 7C FD 25 51 53 92 A7 1D 99 1A C9 49 6E F9
 CF 04 7A C6 00 38 39 7A 65 C3 87 70 D2 E6 0B B9
 5D 55 C0 F4 E3 01 0C 35 EE 8A CC F6 39 9D A4 9B
 B0 13 FA DD AA 30 08 56 C9 F9 4C 2A DB B5 2D 27
 F0 1D D9 7B A3 37 30 63 B6 04 A0 D8 E6 C0 A1 40
 26 41 55 BA 87 C2 F1 78 74 9E FC 46 E2 41 44 DB
 E3 49 81 96 A6 08 43 A7 83 B5 8B C6 86 87 CA 36
 01 EC 5C B0 7C F8 FF D6 2C 58 5C 10 F7 87 7D 1D
 5F 48 DE AE AD C4 04 39 83 E1 CA DA 6D 89 B5 E7
 8C 9F CD A1 44 5C A2 0F 7B EE DB 49 56 2B 20 EB
 85 3E 6B 81 DB 2A 07 DD AB 13 0B D8 97 27 B6 B1
 CD 64 D4 20 6B 87 6D 18 D3 BF D6 B6 41 AB 04 E1
 81 50 36 97 C7 D1 BF 45 65 83 44 2A 76 B3 0B A4
 02 92 22 73 76 10 41 E9 00 36 80 4D 50 CA 7B 73
 C6 C9 35 9D CC 78 38 A9 0B AC 8F 69 AF 97 CF B6
 39 3D 8A EB 39 C4 40 79 3C A1 72 7D 27 C5 15 73
 D8 4F 31 94 C6 24 C4 75 03 B0 E5 B5 B6 5B 0D B6
 7D AA 9C DE 2C 44 8A 96 5F 07 76 F5 8E C4 7E 80
 B0 74 AD C5 D8 B2 CC 97 B0 74 42 56 E4 1D 42 0D
 4B AF 26 BE 20 E1 01 6D A5 AF 5E AD 93 20 61 7B
 20 F9 7F 71 0B 5D 5E CC 0D BB 23 38 CE F7 62 D2
 2A E3 78 25 5A DC C5 87 90 9A E8 24 0A 5C 60 13
 45 2C 0A 43 92 6D 38 A5 67 FC 74 4C 8C B1 7D 56
 D0 72 73 F8 FC 9D 86 E7 8B 57 E7 2D CB 3C 9E 55
 E7 1F D8 13 79 65 92 FF 7F A7 84 B5 DE BF 08 4D
 50 7F AD 83 2F 17 2A B8 E4 4B 30 7A A5 EA 9E DD
 9A E9 8E 18 49 73 FD CB E3 7B 93 78 2A 0E 2F 25
 2C 3B 2E 57 F1 22 D5 45 45 D1 E8 42 A1 44 78 7F
 E9 E2 9A DE DF 74 52 EE 11 C9 B2 D3 7A 55 AA F4
 DD A6 17 49 C6 71 7E E9 36 36 78 C8 E1 F8 54 18
 B2 59 E0 85 3F E1 C1 45 08 BB AE 81 C1 4D C0 B3
 CD 12 11 AD 20 C2 AD FB 56 3E 53 35 99 A3 19 47
 C1 11 E3 38 04 32 A7 54 A5 0B CE DA BE 65 6B 60
 E9 D6 F7 2A CA 38 19 D1 DC 08 AC F2 E5 8C 65 50
 28 93 13 55 3E D5 02 59 1F B5 51 5D CD A3 32 A3
 E6 05 6A C5 C5 C3 F8 20 04 2B BB 5D 11 63 74 AF
 7A 90 D1 96 A3 27 21 05 77 9D 08 B6 CE 44 68 0A
 CF 25 67 BC F2 5A D6 17 B0 CC 4A 20 5E 0D 81 ED
 75 C0 BE 86 40 FF 3A 9F 55 BF 78 FA 24 CA E2 64
 B2 AE F0 71 3D 54 1F D6 38 0E C5 AE BF B3 8A 6F
 7E AD A3 FB B2 E5 44 B5 40 B3 93 11 50 5B F4 95
 37 01 42 CD 05 84 CC 41 EA 76 59 46 FF 90 8B 86
 76 D8 F3 66 2A 70 8B 37 69 46 07 EC 8E F8 33 B6
 5E 33 92 AB DB 80 8C 0A 3C E4 3E 8C 84 E4 58 8D
 19 DD 36 48 30 F1 E2 77 39 FF 72 12 24 92 A9 61
 1F D3 F4 93 2E 4A 5D 64 5B 53 D5 E2 7F 9A 37 8B
 12 E4 1E 99 32 F8 28 3A 5A 5E 0D C0 5F B5 F6 58
 C4 F7 6A A2 D1 4C FD E7 83 64 93 A9 FE 49 26 A8
 C4 DE A6 A5 58 DB 95 94 8F 45 82 C4 5D 19 E3 E6
 7F 43 10 B9 F8 40 CA 03 0A 9B 9C 4B CC BB C4 68
 C8 F8 FB 7B A6 29 C8 7A D3 FD 40 E5 C0 34 DE 0E
 1D 92 49 31 5F E0 69 84 DF C8 15 C8 F1 03 20 EA
 DD 25 2A F4 1B 7E EB 22 47 F7 CC 0B 75 04 78 E1
 73 C2 67 C2 93 7B DD A4 DE A1 01 C2 9B B3 E5 2F
 C0 CF C9 7B 94 39 98 EA 1B AC 71 2A 7B 3E D8 9D
 EE 79 6D 2B 84 CC 44 B6 75 DE 6F 5D 69 DF 9E 12
 68 94 55 E6 F3 22 A4 64 7E 23 63 A5 A9 2C 0C 59
 CE 86 BD E7 77 71 8D A9 3A 87 91 20 9A AF 41 43
 0E 2B 3D B3 8F 96 80 60 4E A1 D7 F2 C5 CA F4 A5
 11 C3 37 9E 81 27 95 77 0D 9A C6 DE F7 7F 0D DC
 C1 6D DB FE 3B D4 1B EC DA 0B E3 D8 CD 9E B5 93
 2B 64 AF 6F 1F 97 0D 4E B9 AC CB A2 59 83 32 41
 AB 43 D1 26 9D 3C 77 4E 69 D4 A3 DC E9 EF 50 FB
 0F 3B 9E 63 BB 40 E3 92 6F F2 41 34 D7 75 37 9F
 EB D9 00 71 37 6F 8D 34 EA 26 A0 BE 0A CE 74 5B
 C5 E2 DB D2 5E AA B5 6B 44 7D 31 E4 88 97 4F 7C
 07 74 8D 4D 02 4E 47 0B 2B 76 46 17 6A CC EE 46
 1C B0 A3 85 51 54 D4 FF 16 02 FD 14 8B F8 69 D7
 19 F6 29 CB 08 9B C0 DF F6 6E 95 24 28 94 FB C9
 E4 04 59 3F C9 05 CE EA CF 79 33 13 16 49 AF 0F
 2E 84 84 9D C0 B6 15 02 94 6B D7 61 29 5C C6 BB
 08 AB BB 21 FB 0C 97 CC 3D A5 D4 60 D1 C8 23 13
 AA 77 BB E8 0F 02 44 5A 31 82 BF 1D AF EF 9E E4
 19 9F C8 AF B0 EE 76 94 CA D1 DA 4E 89 B4 6E EA
 D9 26 41 70 7A BC 59 57 54 6F D3 D7 31 97 FE 49
 2B 0B 5D F3 4E 0F 83 80 14 AF 9F 92 69 00 14 84
 4F 7E E5 D1 2D 5A 43 FC EE DF 91 4E 3C F1 CB D9
 3F 6D D8 15 A6 DC 85 CD BD 8F 83 25 C4 8C 4C 7E
 33 13 34 98 08 BD 1E AB 4A 47 D0 B0 41 89 3B DA
 85 16 E1 BE 1A FB 92 B6 E8 21 58 18 C3 55 81 25
 05 18 3A C8 F7 28 D7 7D 07 0E 9E 1C 01 27 81 41
 83 0A 64 F4 3E F3 B6 0B 6F FE BC 91 3F 0A EA D1
 E8 21 33 A6 FA A7 C9 0B 9E 7B 22 E9 71 C9 A8 38
 8C F5 59 53 3D C1 93 DE 91 84 58 83 63 F6 14 EE
 C8 33 DF A5 57 5A 94 29 5F EB CD 79 62 0B 86 20
 60 1D CE 2C 42 01 6E 7B DA FA 19 B9 57 0D 90 B4
 F0 70 6D 61 D6 24 0D 80 F7 F5 3C A7 50 17 2E C0
 30 1A D8 FC 80 66 08 90 B7 9C EC 99 32 03 33 9C
 FF 49 22 59 A2 94 31 AC AC E3 37 06 85 FF DC F3
 7E AD 93 4E DB 39 56 E6 5B E7 D2 E0 98 8A E4 60
 BF A4 FF 7C 13 B9 75 40 39 38 69 9A 19 21 D2 87
 0F CC 87 B3 6E B9 82 E2 89 30 09 FC 6D 2F 65 D6
 F5 DA 72 1E F1 55 A8 C5 A5 12 E5 F5 B3 6B 78 38
 30 80 8F C9 4B 1E DC 2D F1 87 31 59 8A 7D 7D 5C
 19 08 74 15 A4 07 FE 50 1F 08 E4 A1 2C 8C 40 CC
 F9 B1 EC 88 43 50 65 C5 D1 B9 1F B0 36 E9 50 A3
 DB 20 F2 7E 24 F6 3F AA F4 D0 20 F8 87 7C 21 E1
 3E 76 79 B1 54 A6 96 07 E6 5D 06 E3 52 5F 2F CB
 E6 C9 73 2F B6 88 5D B9 2D DE DB E1 4E BF 5D 91
 77 9C 54 E4 64 AD 47 1E 87 D1 EA 13 BB F0 5A 16
 C3 DA 6E 75 83 2A EF C4 5F DD 30 82 64 CA F3 24
 A0 0E B4 2D 93 CE CE 15 35 47 E8 F6 CD E5 8E C3
 57 3B 41 3F A9 8D 12 61 B8 B1 24 B4 D4 54 9C D4
 3D 1C A5 B8 60 D7 F5 7E 4B BC B2 2C 74 8C 30 F2
 89 0D EA 16 EF 00 BD 43 25 FF 45 B1 AB 90 56 B9
 9E 12 AA 41 65 B5 E5 51 1B 32 B5 05 79 8F 24 15
 8C 19 FA CE C2 D3 3C 4F 70 05 E0 AB 6F C2 3F 51
 38 73 F7 D9 42 18 07 D6 32 81 5A E2 DF F6 33 6D
 B1 59 02 0E F1 0B 46 B3 4F AF 44 82 A8 89 77 6A
 02 58 17 B1 17 86 D3 20 92 C5 7C 95 0B 75 87 E5
 EA 45 DB CC 11 38 6D 7B AE D6 54 1C CB C4 B5 C5
 D5 13 3A 17 24 90 EF DE C8 AA 67 72 49 9B C9 2E
 DA AC 99 AF 13 64 28 39 51 7B 49 16 32 0E 87 4B
 CF 7E 72 F0 40 FB 6D FB 1A E8 82 A0 45 33 0A CA
 3A 1D 3B D8 79 E6 C7 CB D2 19 AD 93 16 DC 4E 19
 88 A3 B4 60 88 74 F9 64 84 D3 DA 00 FF EB F7 5B
 01 C2 FF CE E6 CB 8E 37 17 25 45 A9 CB EF 58 55
 F7 F8 4C BE 42 E3 96 D5 E6 46 79 45 B5 44 F8 C6
 E9 A3 02 BA D7 E1 DE A4 76 13 24 A0 FD 06 1F ED
 29 93 32 6D FE 73 7F 40 B0 20 51 9E 61 8B DA 39
 63 08 3F FC 7F C3 69 75 3F B4 34 D4 70 98 02 1B
 46 8B 01 E2 24 A7 20 33 AC CF B7 75 A4 04 BD 4F
 E6 95 0B A9 E8 10 90 99 EB 3E EB E7 58 F5 59 4F
 27 CD 5E 2E 9E 75 F9 01 0B 8F DC 1A 1A E3 9F 09
 24 8E 79 00 C7 B8 AC 14 76 A0 AF 20 0C D4 B6 A6
 4E B1 FA 05 CA 12 99 CF B0 F4 EE 8F 6F 0D 0F 14
 9F 10 91 9F ED 6D 15 F3 58 79 34 AF AA AE C5 1F
 76 AD A2 13 5B 6D A9 B3 EA 93 A2 CA BD BE 39 0E
 4D 12 84 35 B8 75 2B 30 89 79 C7 28 D7 14 E0 2B
 CE D9 10 CE B7 B0 11 F2 E3 7D 86 59 16 2A A8 C6
 DF E4 94 33 0D 82 66 FD BE E2 1E 5C 98 36 47 1A
 49 D7 19 7A 60 A4 59 45 41 37 09 7C 11 36 8A DF
 4D 6E 66 EB 5A 4F 72 AB 5D F7 D4 F6 A7 FF 4B A0
 C2 8F AC 2C D7 26 84 F8 E4 9D B5 07 55 F0 A4 DB
 07 44 A9 B5 44 C3 9C B4 5A 78 92 17 40 BD D6 D6
 F6 9E F6 89 8C 04 69 52 AB 25 AB 1B E6 39 31 7B
 2D 98 B2 33 F0 8D 20 52 2F 05 32 2E 56 EB F7 98
 AD CA 43 2E C0 5F E7 4A F3 C3 74 1D A6 43 09 49
 AB D1 2D 83 A3 59 A4 0D B8 95 03 77 8F 52 2D E8
 97 73 C5 01 C1 A5 1A D3 99 86 96 19 34 2F 34 D1
 82 CD D4 D4 B9 6B 6B E1 81 55 82 9E 55 7F 66 C0
 2E B7 B5 B1 A3 D8 E3 6F 3A 5D A4 E2 A1 C8 97 1E
 25 AC 95 33 5F 84 EC 83 F4 D6 CF 05 75 4E 95 3D
 A4 62 99 37 AF EC 46 BF AC 80 FB 09 14 5C BB 84
 C6 43 C9 7F 17 1E 9F 04 CE 1E CB F9 EB B5 EB E4
 F0 EE BF 2C EB AA 73 AC 8C F9 8E 95 48 88 41 F1
 A3 FA E2 F5 7D AA 93 B1 5C D8 0E BA 7E 5D 1F 78
 D4 2C C2 9E 05 E5 8C F6 F0 F7 EB C7 6F 88 D9 F8
 43 31 5E 2D 5C C0 CA 80 AC 1D DF E7 5D 3F 0E C1
 BE AF 64 64 43 8D 4C 92 64 8E 9E E0 FF 34 4C CC
 FF 9F 42 66 08 B2 B9 C0 DC 1B 2E B5 36 63 B8 25
 52 1E 97 AB 0E 9A D7 F4 B1 21 7E 76 E7 79 48 43
 7A 85 27 2E 4F A4 9A 72 59 E4 95 95 07 87 92 B3
 4F 9D 4F 29 E1 58 21 CE 62 6C 90 EF 85 63 BF 96
 5E 66 25 03 99 97 BF 88 6C E2 27 6A 28 90 42 D0
 90 92 99 35 98 BA 18 53 62 55 CB F3 24 35 6B 13
 7C A6 34 F8 B7 A3 8E 28 D0 52 B6 D9 D0 06 9E BB
 9E 65 05 C7 E4 E8 67 65 52 6F 9B 9F 47 FB 25 56
 69 D0 99 27 2E 46 34 1C 9B EC BB F0 72 65 40 E6
 78 5B 68 A4 53 84 C8 0A 3B F0 BC DC EB 08 AB 8D
 B9 4B EE 10 92 A5 A8 F8 05 D7 AB 9B 51 31 19 30
 92 89 B2 F6 7C 76 90 0F A6 B9 74 C8 FC 4C 1E 56
 F5 EB FF 9F FD 22 DA 2B 7B D8 AB 3D 68 01 7F BA
 B3 58 AB 49 0C 35 46 56 25 D2 C3 99 6C E5 57 BA
 F0 2D AD C5 4A D8 07 41 91 EC 8E D4 B2 FE 39 3A
 02 71 64 1F FD 84 EE BF DC 1D BA 2A 0D B1 53 DA
 5C 0C 53 BB 56 2F 99 07 66 07 31 59 71 C1 9F 10
 1A 14 A7 A2 2F 72 43 B9 C7 7B E7 2F 1B 30 48 10
 F2 E4 60 03 4E AB 6C 61 5A 42 B4 89 B8 0F FF E9
 BE 41 B1 1E A7 3D 11 9B 90 C3 64 BE F7 80 43 41
 6B 1A 46 A0 22 91 05 A0 1E C0 D7 5E A2 79 9E AE
 29 FD 09 85 91 87 68 E9 CC 46 78 3F EB 0A 3E DF
 2C D9 94 46 47 4C DC 48 AD F3 25 46 9D DD D2 AE
 44 93 23 5C 38 42 92 28 0A 65 88 0D 7C 52 63 CE
 79 13 F4 9F 15 2C A1 85 40 15 F0 3F 26 31 1C F2
 0C 25 3D CF DC 9D 22 AE 4F 43 B6 99 72 FD 89 AD
 4E 9E 0A B0 C2 A4 56 DD DA 75 2B E2 13 9F B4 A9
 56 98 85 79 C3 FB 22 43 21 61 AA 8D 2E 37 13 8C
 2D 71 BB FA 13 23 B8 34 FB B9 05 FD E0 34 0B E6
 29 8D F8 2B 47 A9 AC 1E FC 60 F3 92 3B C6 62 6E
 9B C6 94 43 05 DC 7E 57 09 6A F3 05 7F 29 64 32
 B9 E7 21 B5 ED 0C B2 B1 2A 92 41 DA 07 17 6E 0F
 E7 07 BB 96 18 2F B1 3B 36 7B DF 66 6D B0 95 9E
 82 6C 6A AF 0B 45 88 AA E3 DF 60 5A D6 99 D0 82
 CC B5 78 93 7B 7B AB C5 91 4E 02 5B EC 5F 24 EA
 9A 0F 57 0A FA 83 D5 B2 70 30 2B D4 4C CB 42 8A
 8A EB 7F BF C3 BF D9 F7 2A 84 51 70 72 D9 DA 68
 DA 55 68 DC 14 9F A8 E3 8E F6 4D 25 7A D4 A0 38
 8E 0D FC 60 A1 01 76 0D 0B 8D 5E B0 B8 50 8D 78
 3D DC C5 7E AE 12 B6 0E 4F BB 6E 9E 43 0A 64 82
 E3 A8 86 4B A7 42 BA 18 DB F5 1A 70 FB 38 F5 1A
 02 DD AB 57 4B F6 BC 0D BE 4A D0 B7 9B 55 B2 95
 D4 53 EA 5A CF 4F 47 CA 7B DA A7 25 48 C0 51 A3
 57 E4 2F 1A A7 EF 08 D9 16 6C E2 F4 71 21 8D 7F
 CA 1E 77 2E B9 12 0F B1 47 A3 2C 53 B5 A2 65 45
 FC 89 F4 A4 D1 98 8C E6 49 39 17 68 66 04 A2 EE
 6B 2A CA CB D7 97 C5 2F DC 58 5B DA F2 F2 D7 E7
 B6 C1 3C 03 2D 42 A1 92 9D 66 6C 20 E6 1D 20 CF
 FE DA 0E 0F 39 96 C7 5B 7B F2 78 D4 D0 2E 47 4B
 45 52 34 B2 3C 5F 6C C7 E9 0C 91 14 0C 3D AA 30
 00 C9 10 AE E0 F8 60 18 7F 7E 7E B8 AD CB F9 BF
 48 08 27 EA AB D2 70 60 4C AD 59 55 1F 07 BB 2E
 F5 9E 27 8F C2 30 B6 BE 13 9A 87 A0 3B 99 F7 5F
 5D 42 15 D8 8B 79 DE 04 AC 11 90 8F 30 73 71 7C
 8A 72 09 F7 A1 2A DB 20 EA B7 FC D8 72 D1 60 FA
 CC 3B A0 DB 5D 9B 09 18 02 36 83 D9 41 17 73 45
 DF 4F 8F DA D4 B4 73 50 87 1A 3E BB A6 CE D3 ED
 2D 9F 79 9E 6A 46 88 E6 F2 9C A8 16 0B AE A8 78
 A2 FC 57 62 0F A2 3F DB E9 3F DD E7 00 F4 19 37
 B5 85 D7 82 48 B8 F5 E3 1E 2B FD 3D 01 17 D7 A5
 0F 87 40 2D 47 9E D6 EE 8C E4 C4 4C CA D8 19 FC
 92 85 74 57 53 6D 5E 82 EF 91 0C E7 B0 20 FC BF
 70 6A 48 E1 16 56 10 22 3B 26 E9 D6 99 04 7E 74
 8B 3E 35 A4 81 14 23 3A 4A 10 0C A8 98 02 CE 0E
 92 B6 72 45 47 0F F0 85 03 A5 CB BB D5 D0 80 EC
 9B 50 96 47 02 D6 AF E1 5D EB 0B 37 B8 D5 2C E7
 BD 2D 51 7C EF 83 64 BE 20 7A CA 59 BB E8 04 D8
 DE CF F8 01 3D 73 56 B4 15 8B B9 47 3C 22 1B 19
 67 F6 DD FD ED 2E DA 23 AF 76 F1 A7 B5 10 EC 2E
 A2 32 8E F5 B9 12 5A EA A0 A7 EA D0 FA 47 AF 93
 9A C5 94 74 CF C8 BB FE 65 FC F6 20 BB 54 28 A7
 77 72 FF 81 AA 0C B5 3C 41 92 06 28 D3 44 78 43
 49 ED CA 7B 3A BF E1 35 FD F6 31 FE 32 6C 7F 13
 D9 66 A7 E4 9B 5C E6 0C 7B 2C 8C EB 86 82 F0 81
 A7 BE 55 28 65 B0 1C 52 33 24 31 F6 9A B2 07 26
 52 D6 A4 2C EF C8 26 33 13 FE A9 B3 A6 C7 4E 7C
 96 FB 3E D2 F8 AE 70 29 DB 66 79 60 AE D3 18 46
 C7 20 DF 8F 3B 2A 60 08 0D 6B 61 C2 31 F5 1B 6A
 EC 6E 5F 58 F6 6A 3D CE 72 EF F8 23 C6 C5 49 DF
 93 8B CC 9E 17 C3 80 F0 84 1A B6 77 1E 9D 62 3A
 6B E4 A8 3E 04 3A 1E 43 81 74 AF 6C 43 06 FE 30
 8B BB 89 57 FF 57 74 B3 37 CE 8F 08 6A 08 D1 9D
 3C DC 4C EC 47 83 BC A9 17 43 44 55 66 3F 3A D0
 DB 46 7F B6 AB A0 72 F7 72 A1 A3 99 3D 95 CA 3A
 47 7E 9C A0 8F EE 8B 18 62 0A 1F 92 50 D9 99 9B
 B3 75 F6 2B 89 19 B0 6E 5A 4D C7 AD 8A CC 92 53
 73 05 D4 3B 2A 71 9B 47 FA F6 24 14 F8 29 EA AC
 74 F7 DA 69 AC 3A 5B 73 43 AD BE 08 A1 E8 BD 97
 FD D5 BB 12 A7 3A 17 D9 AB E4 C2 66 03 70 B9 19
 13 55 71 A3 C3 C2 7E D0 87 01 9D 20 58 52 BE 3E
 0F F4 1D 3E EC 3D 55 66 EE 0A D5 C1 F0 CE AF 7B
 8F 19 CB 78 62 16 7B 77 1D 38 EB 41 00 68 F5 98
 C4 C1 E3 D6 1B 70 23 10 6F A4 89 23 25 35 48 C3
 3E 1A 43 D6 55 EB CF AD C8 44 6B 2A 54 52 C0 64
 20 9C 62 D8 58 C6 60 4F 09 CA 61 F2 FD 9E F3 15
 A9 46 A7 9F 16 B9 07 99 E5 34 EA B0 56 7C AA 43
 E6 49 EE 8D 78 C1 AC 54 F3 FA 56 8C 87 F6 37 45
 C3 46 A7 12 65 69 50 CD 59 FC AD 27 84 AE F3 1B
 3D A3 20 0F 33 98 46 7D 60 BD 61 FF 32 EF 6B 72
 94 6A 16 00 3E A4 CA F3 0C 6B 0B 04 DD 1A 84 F6
 1E 37 AB D7 71 58 22 10 F5 50 3C 50 A2 81 0D 5C
 57 7D 65 95 92 E4 FA 5F 65 71 E4 50 5C 3D 15 61
 E2 7D FB 5C A8 82 0B B7 52 4A BB 39 50 5D 7B ED
 5C DB E5 EA 8E FE B3 35 1E 96 75 5B 6B 8B C5 1C
 9D 2D 92 F7 89 9A 0C 92 CC 45 6C 6B CB 5A 85 F8
 97 AD 01 6C ED 3B 3C 15 D2 31 3A F8 8D 92 7F F2
 24 0F C3 F9 77 EB 42 78 8F 75 38 AA FF D9 60 3F
 D7 D9 F4 1B 2B 2D 39 4F DA E4 77 D7 BF CA 08 5E
 A5 BC 21 15 39 DC 19 0E BF 59 3D 36 B1 E9 91 C5
 12 03 A2 7E 27 EE E2 D0 EF F2 2E 8A 5E 9D C9 60
 3F 2E F1 95 A3 86 CA EC 0D A2 FF B6 03 F4 51 5E
 29 82 80 E1 69 3E 4E 14 48 87 DD 26 54 89 8F 01
 08 CD D1 E9 EA B8 85 F8 51 85 93 5F BF D3 B1 CB
 2B 85 D9 1E 22 A1 14 FF 86 23 5D 27 9D 18 CD 80
 1F B2 00 D4 10 2E BA 5B 33 26 14 A9 CB 28 29 FA
 C4 15 C5 DA BB D4 1A 8C 48 72 7E 31 B0 09 00 02
 9B 7D C8 23 A3 A0 6F D6 E0 0C 0A E5 D6 B7 96 7A
 64 5C FF 8E 46 FE A7 98 73 C6 52 B9 A5 D1 05 40
 3C 0D 34 0D C7 99 92 80 13 92 AC 04 93 68 50 57
 5A 16 34 42 3D E3 01 7A B7 DE F7 B4 90 0F 58 6A
 43 60 2F B3 2A 01 DB 06 65 43 75 0D 95 72 A2 6F
 E6 7F EF 23 5C A7 08 00 3C 07 2F 45 C0 61 CD AF
 F0 3E E2 C8 53 16 12 55 FD 0E 6F 1D 10 F9 A9 87
 9E 3D 0D 6C 4B F2 18 74 91 30 C8 40 52 D6 61 F1
 02 F9 30 63 D5 A5 A1 54 35 9A 32 C8 82 28 E9 CA
 33 8B 7E C4 4F 9F 27 01 A7 A7 DC 1E D6 2B F4 9B
 55 9D A2 B0 26 00 A6 F1 5C 21 9F 80 2F 02 0B D0
 50 E4 74 22 D7 85 68 FF 50 63 51 0D BA 6E 7F 80
 FF 77 D2 32 95 4B 35 99 B3 EA A9 E4 AD 03 EA 0E
 90 F1 BB 61 39 A1 1B CE 7B 45 E0 68 45 B2 27 7E
 D1 0B D7 32 2D 2D 81 50 51 34 A6 32 7D A0 BA 27
 CD 6B F9 42 F8 CF 0B 30 BE 75 CD 2B CF B2 EF F8
 AD 70 7B DD 01 7D EC 3F B6 4E 17 4C 24 0D 39 41
 8B B8 D6 E8 B6 0F 7C 6B F9 E4 46 C3 BA AD CE 9D
 A0 C3 68 F8 BE 09 D7 42 20 2F E6 C7 23 15 BF 6F
 A3 FC 7F 90 01 9E 15 04 DD C4 D9 3E D5 CC 08 B8
 80 58 B1 22 0E BC 35 85 84 0A 66 F0 77 11 E7 D9
 81 DA 03 D7 87 61 44 F2 1E E9 F5 CB 4F 73 69 D3
 51 F9 C2 82 9C B8 67 3D F6 36 D9 9A 16 C8 CF 7F
 6E E0 6E FD 4D E8 DE 23 9C A2 8F 38 E7 96 1C 69
 30 1B F0 CB 58 49 50 DD B8 F8 FF B5 2B FE B3 D3
 BC 58 B9 3E 0A 7C 86 CC 1F 60 EE 8B 5F 74 E1 A4
 45 95 9D BB 85 A5 96 25 45 2D FA C1 E5 82 B6 8B
 8E 67 E9 C8 9C B8 04 2D DE 4D 98 1B 75 A7 CB 19
 E4 10 02 63 41 DA C3 6C B7 A5 20 41 83 FA DC 70
 CE 8D 29 10 8C EE C9 BD B7 2E 58 BD A2 96 9F 89
 45 08 EC ED BE 0A 9D C6 78 8C 18 36 1B 09 AB 69
 1D 9F C4 E2 BB 11 D2 60 FE E2 ED B3 97 AB 36 8A
 CE FF 25 A1 13 DF 43 4A 98 32 7C BA FA 22 EA B1
 72 27 15 5E AD 62 9F 72 D3 89 56 83 2C 30 26 B0
 99 7D 1C 2F F1 33 4F 8D A1 4E 07 97 28 39 6E 94
 78 B3 55 1D 1B 77 76 54 2B 54 20 5B 29 9B 3A 40
 D7 4F 8C C2 DD 62 55 2B 50 F9 34 1D 98 8E 82 76
 E7 45 B9 F5 03 BE EA 90 26 A2 8D BB 17 C2 86 6F
 51 70 9B 91 38 2B 3E AD 89 2D 04 93 E1 BB 03 A3
 DE 55 2C CD A1 FC 90 1C 09 12 BA 12 F2 AA ED C1
 DB E0 72 52 AC 81 F2 A5 C4 B5 7F C1 35 C9 EC 69
 1B E6 0E 7B 36 6A A2 77 0C 7B 92 98 7C 62 B2 67
 81 E0 E9 8A 51 B0 A3 FC 6C 52 DB 5F 09 9B 02 B5
 57 6B D2 B0 62 74 EB DF 40 86 C4 0B 26 9B 96 E4
 E0 77 2F CD A2 67 45 C7 7A 42 8F 97 6B A8 19 1B
 F8 5E 06 4F 04 CF B2 47 15 29 56 FF 45 2F 61 28
 60 9A 84 B4 60 5D AB 1E AA 15 7E 12 7D FC EA 6D
 08 77 29 80 B8 3A 72 CF 49 72 BF 25 43 B1 01 88
 1A 46 4B 4D CB A9 65 7D DC 4A F3 51 D1 0D 90 85
 44 98 38 9E A5 38 8E 00 9E CC 7E 6F 78 21 2C C3
 24 E9 0D 97 5C E2 11 92 16 B7 E8 85 05 B4 CF 14
 4E 27 4D D7 C8 C5 14 EE E4 6C C1 34 68 4A 0B 49
 02 A9 11 99 AE 14 7A 4F D1 4D A6 03 B9 8B FC 60
 7F 55 B9 2C 60 D1 B4 42 52 56 E6 53 C8 C8 99 E5
 C3 14 78 67 A8 B0 A0 26 06 DD E7 AD 92 1C 49 48
 2B 90 75 54 B1 E7 AC 62 D3 F2 48 EC 52 D3 C7 0C
 A9 F1 C3 34 52 B9 10 4B 05 E7 D9 B1 8A 23 A5 69
 2E 8B 9D BD 83 E2 BC CF 92 7D B6 FE 63 0C 37 67
 F0 98 2E BE 60 63 A1 59 44 9B 42 41 6C 16 A1 6D
 33 6E D1 76 DE 75 FB F6 F4 D5 BA A3 FF F2 DF 4D
 EA 12 0C 75 97 94 D5 07 E9 00 C1 7E 87 D6 8E 8A
 31 12 71 AB D6 52 C8 55 5B 68 38 F3 C4 90 50 51
 DA 7B C7 2D 2D C0 53 D5 31 5E BF 00 50 AC AB B4
 71 AC B2 B1 8F 98 E6 D7 40 4A 29 87 EB E4 BB AE
 3B DE 52 B0 2A F0 7C 28 6A 62 83 A0 CC 67 86 FD
 E3 03 C7 AF C3 68 0E B4 16 64 5D 23 E4 CF 21 5D
 FD 8C C2 20 EA AA B5 23 4C 9E 58 B5 20 12 6F 4B
 26 67 E6 3A B2 40 5D 7A ED F0 D5 8B 06 E7 00 43
 4D 8D 20 1B FA D2 00 EA EC 82 53 4F EF B1 2B 68
 19 8D CA 51 C8 B4 B8 47 24 C6 A4 D2 98 0D 1C 66
 23 10 21 45 D0 0D 85 63 D0 55 AA 08 C6 31 D8 0D
 3F A8 0D 4F 80 46 FB DF C8 A3 47 0F 6D 7A 63 31
 C8 5B 88 F2 EA 4C EA 46 7C 0F E5 C3 83 FE 6A 4D
 AC 34 75 8B 27 C3 1B 28 AC 17 58 9F 7A 27 C4 48
 21 FF 16 8E 1D 01 D2 87 17 9C ED 66 BD 80 59 9D
 00 14 77 37 4E 6E 41 17 D7 6C 79 11 E2 26 80 15
 CD C9 6E 05 E9 6A 9B 61 88 51 61 BB C5 60 0B C6
 50 E9 C6 F2 70 36 6D 18 B5 EE CA 39 D0 90 09 42
 5F 4E 9E A2 0D D2 9A C3 70 03 8C 02 74 BC 9E E2
 A8 78 C6 62 C4 0A BA 8B 61 90 66 5A 0E D9 4C 10
 5A 49 80 7C 1C 47 0C F7 4E 51 B8 60 83 F3 42 4F
 BA 82 E6 88 5C 04 F8 BB 33 65 E1 F0 3F 32 23 48
 B3 A8 FC 54 0D 5D F8 F3 F1 4D 12 46 63 17 72 C7
 9E C9 32 C0 F5 00 2F AE FC 78 48 CD F9 B9 BC A4
 4E 10 01 7B 5A 80 D0 A8 89 7E 04 10 76 61 67 37
 FF A4 4B 08 BE 24 F5 CA 0B 67 DD 1B 52 3A E2 95
 C4 4B 7F DE AC 71 8D 49 55 92 D3 52 84 50 6F BB
 95 58 F2 9C 44 7F BE 66 E2 E9 E0 2B EE 4E AF 81
 07 64 1F B6 85 F6 2B 17 B2 67 90 62 E9 9E 6B 02
 D3 DC A3 35 82 6C 50 C1 F7 91 C2 DD D0 82 67 AD
 47 25 7A 52 33 D4 08 5E 20 1B E3 C4 11 94 E9 4B
 DE 84 58 A1 A9 4F 29 F6 25 C8 4E 1A 40 63 28 0F
 5A 42 9B E2 95 8D 94 BB 92 A9 F9 BA 83 1C 26 8A
 7C 16 AF A0 AF 80 26 56 00 D8 AD DE C1 57 33 7B
 01 DE D0 CB 12 22 7E 2D D0 CD AE 61 D7 2F 20 98
 C6 17 CA 24 54 31 3B A5 4E DF CF F1 98 34 3A E1
 B3 EA AD CA 65 EE A9 9F 99 8D AD AB 21 C8 A9 36
 A2 D1 F9 DF AA 10 30 C3 4A 84 62 05 4F 26 98 A7
 48 02 13 9E F9 FE D3 F9 61 6C E9 3E 44 3A AF 79
 34 37 7C 12 3B 83 18 EF 7E E0 3E 1B 62 7F 07 37
 A7 DD 07 9F 62 52 CC E7 03 27 4F 86 0C 61 DB 48
 17 9F 45 BF 58 DD 67 83 BA EF 8B 7E 30 5E FB CC
 50 EE 9A D8 6C 7F 17 C9 EC 02 57 71 F5 2C 81 49
 BA 68 BF FB 29 E6 22 82 B4 D3 53 13 88 D7 AA 32
 FF AA DA 03 70 90 81 C7 AB 42 D7 A5 A7 CB 77 0E
 48 CD 37 22 59 26 38 C8 B6 0E 6F 09 83 75 D3 23
 3F D9 9E 09 4C C0 09 41 A5 19 9E A5 E3 A1 A8 78
 74 20 F3 4A 44 62 55 FE A4 5B E0 88 EF B3 77 20
 A5 2E AA 10 A4 29 47 23 6C F8 60 5C 44 72 8B 5F
 C9 AE C4 84 AA 08 08 F4 AB 70 87 3A 30 97 25 E7
 DE 25 0C 67 B2 C7 70 81 7E C6 A4 2B 3F DE 39 C9
 39 3E B4 DF CB C2 CF E3 C2 E1 9D B0 0E 85 F8 7E
 E5 F2 F9 6C 16 F4 2A 6C 4C DD 69 8E 51 2A 1F 0A
 B9 EB 77 DF 73 95 F1 82 7A CD 8A 8B 4F FF 13 8B
 56 1A CE 7E 92 30 D4 92 6B D5 31 29 64 2B E4 05
 E6 3B 67 55 CF 62 53 F4 72 CD C9 8E 3D D0 79 FB
 FF 9B 4D E3 1D F2 2A FC 90 8F 5A 73 3A 61 6E E3
 A5 96 CE DF F4 1B 47 1D 32 E4 0C C5 9D F3 FD CA
 A1 25 17 53 48 B2 57 CA 4E DE FD 70 BA AA 1A 3C
 B2 36 15 72 11 CE 31 F7 E6 A5 8D 6C 1E 96 96 E8
 9E D9 3B D2 6E C4 56 55 57 C6 53 E3 09 E2 CA 07
 86 BA A1 C6 D0 28 5E D7 6E F5 3A CC 26 39 E5 74
 A2 A4 50 11 AC 48 0A 4B 86 B9 9F 80 EC EC DA B3
 B6 8E 68 A0 31 29 A9 A0 ED A1 C2 8E 41 60 3D B7
 AF E6 CA C4 63 7E 34 62 FD 8E BE EF FA 17 2A 2E
 31 EA F7 C4 EC 95 08 8E 3D 82 E7 F3 36 BA 03 15
 91 0C 08 EB 18 7B 68 47 FE 9E 3D 2C EE A8 35 93
 80 9D 1C 78 5E 23 58 22 46 45 84 C8 E7 14 7B 6E
 0C B1 6C 72 D9 5D F0 52 8B 10 3D FF 7A E9 91 79
 F9 D2 94 E2 9F F9 85 04 50 99 DA 86 9E D7 6E 01
 CD 4F 8B 70 16 48 76 2D 8D BC F8 CB D0 3F 63 AC
 F5 17 9F DC 31 8C F6 2D AA 70 6C 49 E0 6C E5 F7
 B2 ED 75 FC 53 24 7F 29 EA E3 78 FF D7 45 61 A5
 69 3A 38 B8 6E 60 4E 04 27 0E 26 25 A2 19 12 7F
 89 4A 9A 14 83 7A DA E6 23 DC 42 95 C7 73 CA 9C
 AD B9 F9 B5 ED 40 AC CA 04 35 4A 4A 5B 69 66 19
 0C 78 35 02 3C AA 3A 7C CF 78 B6 4C AC 6E 1E C6
 8D 27 D8 10 73 E0 71 27 24 B0 07 DE 20 67 AA 6C
 A6 7C 77 CB 75 92 0A 17 CA 50 00 AB D9 9F F4 D6
 A7 70 90 14 B2 12 7C 8F 45 FC 1B FB 09 FB 9E D4
 DC B0 94 15 CF 64 8F F1 D6 32 DC 1C 38 E3 28 EF
 E2 63 69 D8 67 CC 91 16 54 6C C5 A5 EA 0E 8C 85
 25 17 6F FF 1F E4 C2 0C B3 C2 64 FD 98 2E 57 01
 08 A9 D3 69 04 49 34 BD DB 20 D4 E8 29 CC B5 C6
 94 40 9B F4 EF 2A 69 27 ED 0C 0C 1C 8E BD 04 36
 43 7C 14 81 A7 68 96 4A 68 0B AD CF 75 98 9A E8
 40 87 32 33 57 9C 63 56 33 1B ED 14 D0 69 C7 43
 DC 1A 52 37 EC 5E F5 B0 45 3D 79 3F E4 62 60 1F
 06 17 DB 9C 3F C9 E4 5E FF 6B DA 2B 18 73 88 3C
 7B 28 D6 B1 98 D9 BE FE AC 75 64 C1 8C 7B 21 6F
 03 52 74 A5 DA 36 99 4D 0A C9 D2 36 72 6D 1E 53
 E9 6F 64 E0 E3 01 2C 59 DA 52 D0 D1 0B 3C CF F0
 1A 0D 4F 10 31 C8 93 C7 89 D5 AB 5F DB 25 78 77
 D8 03 2B C9 07 11 14 AC F8 02 33 A2 8A F3 FE 18
 5C 7E 11 A6 DA 50 21 E0 24 C5 59 F4 82 82 66 F0
 8D DD EE 6C 11 58 FB 9C A0 C8 7D 8A 52 FB 69 82
 60 8C 8F 34 DB 79 0C 68 5F 55 59 42 70 E3 D9 6F
 3E 65 40 90 77 1C BF E0 7D 83 3D 5E 3C 77 FF 94
 CB 48 63 14 6E 0D F5 74 29 E5 8B 5B EC 63 60 5D
 57 6E 21 4D 70 75 8E CB 5E D5 31 00 E3 BB 95 19
 F3 48 09 1B AF FD 8B 07 73 C9 67 C3 31 BD 7C 75
 F3 FA 5D D2 76 F0 56 3F 96 C1 9B D8 A8 C6 5B 15
 87 98 5A AC BD 29 5F 1D 54 C5 F2 5F FC 02 83 13
 E3 B7 CA A0 CE 2C 51 99 28 ED FF 91 87 F1 64 42
 35 9D B6 87 F8 57 C7 F0 3C 40 F3 6D D6 05 79 7D
 FA C8 58 2B 35 68 93 80 02 E6 CD 71 A7 FB EA 4C
 2E D4 1B 48 1D 8C E7 8A B1 1D AD A4 E4 50 BD 37
 C5 E4 FF BE 98 2A 84 52 B1 76 67 1D 89 35 88 C2
 60 69 B4 D5 86 F5 C0 F5 B5 0F 97 73 B4 0E 09 A3
 32 EF 66 F3 18 C7 FB A9 DD 5D 80 15 25 E7 E4 A1
 22 B1 FD B4 AA 3C 5E 82 0A BC 25 40 C5 23 A7 B0
 FC E4 B0 60 E3 41 E6 FB 90 FB C7 AF 6A E4 D9 4B
 8F FF 2B 92 7C 06 C2 B4 DD A4 28 30 C1 C8 05 0A
 39 C1 D0 14 F6 0E 07 B0 83 CA 7A 85 EB E6 68 96
 EA F1 B8 C3 9E ED E5 A0 42 D3 1F 5A 54 15 BA 5F
 16 6C 8B 4E 50 64 A2 08 C8 39 C1 A3 18 EF 6A 19
 0D 46 AF 13 AB DC 6F B7 9F D6 5F F0 F6 9E 34 ED
 C5 4B EA 3D 65 5E E5 66 F2 1A 6F 2A 55 A2 AA 20
 D2 7C 7B 89 30 F1 57 D0 A1 59 30 FD D1 83 12 C0
 41 34 31 4C 5B 37 6A 69 DE CB BB 28 DF F6 BC EF
 A2 43 C7 1E 8C 15 20 80 80 BC 25 53 61 29 57 C3
 E2 FF CA AA 71 C3 6D AD 8D 86 FE B9 F7 7B 1F F1
 2F 3D 57 3C 11 3E 38 0C 64 00 EB 7F 69 D4 F6 AA
 38 87 F0 7C 34 8A 42 3E 1E 8B 26 3B 59 F7 53 4B
 84 B9 16 DC 73 EE 7B 3A CE C8 36 08 37 7E A1 9E
 87 9B 55 64 6F AF 90 BB 00 E9 99 B9 8D FF 2E A0
 E0 E0 C6 04 D5 DE 82 26 10 66 A0 FA 3F CC 36 8F
 06 56 79 79 40 C8 12 28 F8 32 FC 66 8B E9 93 9E
 01 7B 43 C0 E5 EF CC 10 CC D5 32 F9 09 1A 68 8E
 5B F3 69 1B 11 10 BB 93 0E A6 09 05 69 08 0C 9F
 F5 8C C7 5D EE E1 53 ED AC AB 7F 6D B2 E5 DA 26
 A7 15 6B B9 B1 B4 5B E3 A1 0D D7 CF 5D EE 89 43
 9A 0A ED F0 41 EE 7D 0C F5 C7 3A 29 BA 3A C5 8D
 0E D4 41 0A 71 BB D9 69 8B DD 1E A4 A3 ED B9 48
 77 98 F3 FA AA 49 36 13 B5 80 3D 56 0C 30 A3 7B
 0A 76 BF 2C 9B 31 2E 06 6C C5 EA C4 72 E6 42 7F
 B9 9B 55 08 2E 98 0F C9 82 CB BE BD 77 C5 91 AE
 44 4C 21 DC ED FD C9 26 66 81 B6 AE 35 E5 35 E4
 78 D6 B7 F3 49 A4 29 00 AF 1B 2D 66 98 88 78 B9
 94 84 DB 0D 03 93 6C C4 62 61 17 EC 4A 47 F8 B3
 0B D5 8C 88 D2 44 AE BA AB B2 06 3B 3A 98 58 0F
 C0 C5 23 F7 C3 77 EA 3E F0 74 BF C0 3C 08 CA E5
 84 C0 DC 08 07 39 6F 69 87 63 D2 6F 46 FC FE E8
 9F 38 48 B8 EC F5 48 3D 8B FB 9C 88 5D E5 2B 8E
 4C 27 23 29 2F A7 09 DD A0 6E 9C C6 91 C5 B5 E1
 D2 A1 BF 31 99 B8 62 0B 0D 39 D5 3F 19 A0 55 C9
 65 67 1D DE 44 2D 7D 73 58 78 27 53 29 A5 18 B8
 34 8C 0B C5 EE AF 51 5B BA 50 05 28 25 9E AB 4F
 8A 54 8B 31 76 9F DA 55 F5 ED D5 D5 8F 84 AC 17
 17 1A 4E FD 82 93 7D A8 7E 9E 6B 5B 81 74 3F 60
 93 90 A8 BF 69 E8 E5 ED A8 CE 38 6A 7E 55 07 32
 7A 86 88 07 C4 77 F8 B4 4C EA B9 B8 7A DA 43 4D
 09 49 F8 34 F8 92 6B D3 85 B3 E2 BC E4 26 7C 0D
 4F 69 7F C3 5A 9C D3 0D 31 02 0B F4 29 54 46 2B
 16 0C C3 55 16 93 7B 50 A1 6E ED D9 3F 76 48 F9
 19 F1 23 37 12 12 1E 04 7C 37 FE C3 83 8D 3A 2A
 E3 9F C9 5D 31 0A 43 8F 53 9D 44 0C 91 60 43 22
 30 5E 29 62 DA 5A 69 61 5A DD 05 0C A6 71 49 1B
 C0 9F 78 7F 9D 0F C0 2A 9B B5 AC 95 94 99 EF AB
 BB B8 09 10 75 D0 31 F6 C9 32 D8 DE A1 00 8F E4
 31 72 76 CB 51 50 1A 17 FA 23 7A 64 53 E8 6A E4
 4A 8A E4 3D 32 AA E2 F3 FD FC 11 72 DD 04 E6 5F
 46 C5 F0 9D 39 8D BD D0 4A B4 E9 A5 13 E7 9E FF
 9A 95 C5 41 CC 74 39 A8 A5 0A 40 59 B8 0B C9 AD
 5B 92 13 3F B4 DE EC 2F 3A C5 79 4C EF 9C 0C D1
 04 51 B8 91 ED 95 96 89 E8 7A 33 81 F4 6B C4 8F
 69 4D 07 AB 8F 3D D2 F6 BD 96 31 F0 B4 32 E9 6E
 1E 05 5E B1 6A BF E9 A3 AC 60 7B 66 EB 47 D4 0D
 05 56 A3 77 49 3C 3D 47 0C 5E 0C 1F E9 6E ED AE
 47 DF A7 CD 2D 17 BA 35 10 EC 1D 05 90 7A 29 CF
 B1 85 F5 58 55 D7 73 4E AF 8A D8 37 8A 54 40 72
 2B B1 6B 3F 4C 6C 51 D3 E5 2B C8 DD FD D7 78 60
 E3 13 25 36 49 A1 6B B7 8A C5 39 98 0C 04 42 FE
 22 12 93 BD 92 04 5B 3F 54 30 38 63 A6 01 89 6F
 CC F2 1F 3F BB D0 B5 5B 2D 84 6C 67 D7 5C B9 8C
 65 93 B7 9E B5 14 01 32 33 26 6E 2F 31 20 1A 27
 3E C9 1B 44 B0 03 7B 8F EA 0E D2 64 4C C3 82 FC
 6B B9 71 A3 EB 78 4F 67 A6 A0 6F 5A D8 85 19 06
 21 64 6E 12 97 00 2A 78 47 5C 9B 96 98 6B 8D 83
 6A 6B 3E 1D 68 27 AA 89 29 69 FA 90 0D 00 DE E5
 D6 D5 BA A1 FF DF 79 58 08 D4 4B 23 87 7A 8C 58
 27 DE BB E9 D5 70 3A 44 28 72 B7 FF 6B 91 B8 3B
 D0 40 6A 15 4E 27 E7 C7 D5 FA C1 30 75 E1 D0 9C
 CE 66 8B 62 3A 03 13 5A BC E0 06 59 2B 86 D6 6E
 83 A7 EE 57 CA 93 63 EB E9 A4 59 CC 4F F3 9C 4A
 24 41 8E 4B 44 22 73 84 7F 3E 4D 8B 93 92 0B 58
 D0 BD 33 D1 9F 56 71 9E FD DB 33 1B 82 3E FD 52
 88 6A 41 59 CF D7 B9 C1 97 26 C9 A6 55 73 92 DC
 35 63 27 AF 11 E7 0B DC 90 96 A9 51 3D 13 B0 36
 1F 97 B8 3A C8 9C 85 DA CB 57 7D 83 9E 8E AC 5F
 F9 3C 6F 94 64 DB 5C 0D 6B 00 58 BF DF 9F 37 0E
 32 15 5F 9D 62 50 DA E1 46 96 9C FD 2B 16 28 87
 7E 2C 3B 13 67 DC ED 18 67 F3 46 6C 19 0A B4 79
 DB 67 CC 9A 6C 38 4B 80 4D 68 FE 2A B3 37 E1 53
 CE 31 77 52 FE 99 D6 7D 8C 9C 70 2F 8D F7 5D 45
 16 2C 17 3E 3B BE BB 47 25 18 9E 60 C8 47 65 5A
 3F 9C 9A 64 85 A5 62 98 39 8C 3F 4D BB 80 5B 3B
 F7 CB F9 EA 5F 9A 03 39 4F 31 4D E7 A9 F9 21 17
 64 19 CE 26 CE 72 86 2B 22 67 13 20 42 48 B1 C4
 38 1C 69 A3 DC C5 42 31 CF B1 55 A4 01 F4 0A AB
 00 06 EC F5 15 0A 2C D1 B5 60 96 FE 04 73 38 74
 00 27 06 6E 51 CA 9D 78 8D 8A FB 7B B6 11 3E BB
 EE D8 B8 2D 1E C4 E9 C4 7C 7F 62 7D C6 7E 79 09
 8B 03 18 C1 61 CB 8F A3 F4 DC 42 7D 78 22 8A 3C
 F3 5F 41 E1 B8 42 A6 4A A5 47 AA B5 05 42 35 89
 62 8A E0 B5 57 92 0D 00 AD 6A D9 79 F3 27 46 A4
 94 45 0F C3 50 FA 7B 95 B8 40 18 2E F2 28 34 84
 DD 2B E5 AE 4B 41 A2 A5 70 40 46 D9 EE 9C C0 8B
 AD A3 ED 63 FD 5D F6 DC D1 DC FF B7 F5 A5 5D A3
 50 C0 4C BB 57 65 56 1F 29 2A 4D 48 63 EC 88 C4
 81 04 2A F7 6E D1 4A 0E 8A 38 3A FC 71 D1 F2 F1
 E3 FC 73 0F 4C 27 3E CC A7 DB CA 2A B5 BA FF 61
 6F 23 1B 89 BD DC FB 48 4F 52 6D 2E E1 09 7B E1
 F2 00 3A 5D 63 8A 3A C5 6A E1 BC 7A 27 3D 14 42
 B4 87 21 FE C3 9B BD 67 09 C4 79 B6 06 9B 88 D8
 28 D1 1E F1 1A 86 01 B0 58 A8 6F 73 1F A2 50 DE
 F2 21 70 7C EC 27 99 5E 3B 1D 80 4D 74 FE D3 1E
 60 83 6B 1B D3 82 22 50 5C F7 9F 90 60 36 53 B2
 37 81 98 C9 F0 8F 35 01 96 B0 04 61 6E 6C 87 B2
 BF B2 AE A7 F7 6C DF 09 89 DF B5 CC DC 85 A9 A6
 45 47 E1 BC 3B 73 32 3E 56 77 FA 35 0A AE F7 03
 49 F8 09 A3 BD D0 91 A7 DB B0 E8 C0 C4 39 FC 54
 66 46 C7 3F 9A 96 DB 90 D9 D4 32 03 AD A8 B9 B0
 7E FE D2 19 DB 73 95 48 C4 23 47 DF 35 57 5A 31
 A5 D8 CA D7 B5 53 AE DB BE 6F 28 98 B5 81 C8 15
 09 8B 06 D4 4E AA 29 BD 63 BF 50 99 EE 4F FA D9
 E6 1F D7 6C D4 F3 67 3F 2B 00 E4 12 4E F7 D1 D2
 47 EA 84 C9 53 17 9A 40 94 1D 89 0B 64 B0 70 91
 EF AF 6B 50 F7 0E 6A 49 3A C8 47 41 04 46 32 AF
 CD 14 07 F8 DD E9 58 F2 8E 0E 72 31 97 7A DA 06
 5C 1B 8D A6 C7 6B DD 17 66 69 9F 87 36 87 EB D5
 8E DC 13 3D BE 78 74 C7 D1 24 30 A3 EB 88 1C 95
 CB 00 B5 05 E3 38 C3 F6 17 C9 D5 98 67 F4 FA F6
 36 50 B3 22 85 F8 1F 4A 1C 83 6A 24 EA 38 55 E2
 6B 36 48 80 EA 21 02 F9 18 49 2A 25 46 F4 4F 15
 53 C8 8A D2 C4 CA CC 65 F2 73 6F 42 26 6B BE 46
 49 A4 6C 0D 8D 41 AA C9 F4 A7 1B 26 82 E9 BE C3
 F2 45 E6 DC 55 6B B9 BF 47 97 F9 83 AB E5 4A 82
 1F 7D 66 92 85 85 72 5A 01 E9 61 BB B2 90 39 0A
 B7 DF 9A C1 71 53 DE 03 D4 88 7C 89 C7 DD ED 20
 8D 14 3C 11 29 BF 42 D6 87 E4 24 43 D6 A6 E7 0D
 C3 D7 E4 8F AA 58 72 C3 C0 1D 97 93 9B 16 CD D1
 9B 79 78 80 35 DF A8 2F DB 50 BD E8 8D 91 B2 E6
 1E D1 D1 E7 9B E0 C0 64 7F 95 23 3B 0A C3 E1 3B
 DC 4D 6D C2 62 B3 EB 8A 5B 3A 8F 5E 2E E4 F4 53
 8A 1A D6 15 FD 84 6A A9 33 C8 36 54 B8 E8 9C 95
 E5 18 86 B6 BA 4E D6 28 E4 C7 5F 6A 77 CD CF 02
 24 98 E2 38 FB 03 9E E9 B4 5F 39 F1 84 E8 6C 46
 55 B2 BF 51 AE 86 62 15 E0 25 4E F1 63 75 3A 0E
 CE 55 EA F1 B7 E0 E3 2E 63 E2 E6 51 CF 92 23 22
 4B 91 E3 90 06 AE 6E D1 D7 96 33 9F F0 3F D9 2E
 25 30 BE CD 0D F1 DA 5B 67 3C 82 09 9B 5D 32 DA
 BC 05 2A 51 AB AA B9 E6 F8 3B 1A 87 CC 97 51 78
 C6 64 F1 F6 16 79 BC 43 46 D4 75 83 EF AB EE C7
 2C CF 4A C0 2E A7 93 DC E3 C7 B4 D3 CA 3A CB 55
 4B 92 72 74 FB 67 D5 F9 7B 26 90 3B F6 94 50 48
 FF BB 40 C7 54 D8 FD 45 8D 6A 2F 3E 69 22 41 1D
 7E 2C 67 CC C4 28 F5 35 1A 17 33 93 3D 44 79 A3
 CA C1 1E E8 BF 0C 82 64 D8 32 1F CC C0 60 61 4D
 1F E2 6D E7 22 D5 9A 8A 2E CF 32 51 58 52 40 B5
 FD 61 5D F1 9E 57 C2 3A 99 72 83 A1 04 D5 02 94
 13 1D 8C 22 B0 53 57 9D C2 84 60 65 15 78 D9 35
 0E 70 8B 47 03 08 21 C9 F7 E3 A5 B5 B3 17 72 5A
 77 23 0E 0E 79 85 BD 38 2C B6 75 70 4D F7 A1 AB
 B1 C0 DE 38 7F F9 D3 41 9F 55 23 17 54 0A 2F B9
 7C B5 A0 B0 4A 85 0C 97 D9 57 B1 A7 9F 98 C0 46
 F8 ED C3 A2 BB 52 B2 F3 28 34 63 85 A5 06 F8 43
 55 1B 44 FE 00 D0 D4 8B D8 3D CB 5A 23 17 36 8C
 7D 56 5F F0 1D 52 0E 1A 28 10 F1 A6 E1 47 91 5E
 E9 4B 7A 4C 70 1B 99 A1 39 F6 D3 AC 28 BA 17 10
 E4 B0 9B AE D4 05 E4 9F 2E 85 6A BD E2 49 7C 89
 25 3B D5 B8 23 FD 27 9B 58 F3 6D 88 8B 06 9F 94
 1B E1 9D B0 0E 82 A1 8D 12 E2 2E D6 74 4B 62 6B
 37 29 63 D7 BD A6 66 BC EB E6 2F D3 2E F9 32 11
 CB 66 13 A1 46 45 EB 46 F1 66 FA 9E 27 13 10 53
 A2 7D 59 1C B3 3D 68 F1 C0 4D 49 43 2D DC F2 F5
 8B B6 C7 5E 49 00 A1 48 90 9B 92 5B 61 38 65 53
 47 D8 90 5C FF 8D 3A 71 2D 95 78 40 4C DA 75 C7
 46 74 17 5B 37 51 D0 FB 25 4E 69 8A FC 60 5A F3
 EC 4F 2A C3 2D 77 2D 6D 22 1C 18 1C BE C9 51 F1
 A2 77 C5 62 70 2B 1A 71 87 7A 88 79 99 E9 1C E0
 54 7E 74 A5 CB 5A 52 BD 66 B3 1B 15 E7 D5 5D 60
 39 4A 4E D1 A4 7B 3F CA 06 50 87 B4 E6 BE 08 43
 D2 86 32 8C C3 B5 14 B9 5D C9 2C 6B 6E 7A 61 55
 70 29 E0 F5 F9 37 CC 56 B6 69 BA 37 4E D3 C5 11
 9A 87 A8 8E 02 FE E1 0A 12 BD 81 58 7F D8 FD AA
 98 2C 10 BD 96 7D F7 C9 1E 76 86 EA 9A 81 C7 C3
 31 0D 39 F0 B4 F0 3E CF 0B 8A 4A B7 6B 06 92 7B
 45 EB 7D 0C 9F 1C 80 0D 0D 72 25 BF 03 3A C8 C3
 C6 D3 70 DE 5C E3 7D D1 75 F8 0E 29 F3 72 61 83
 76 03 CF 7D D4 90 9C 36 99 6C 37 20 EE 85 AB EF
 B8 02 A6 F8 EE 33 92 00 98 89 10 81 29 FC 13 EB
 76 8B 26 4D 40 9B 57 7E 20 50 25 CD 2F DA D9 2D
 82 6C 24 C1 04 AB CF E6 89 5B 63 9E F0 42 34 04
 15 B7 A9 6D C1 A1 BB 3C 64 2F 87 91 05 F2 D9 39
 F7 B3 C2 CE 19 23 D9 53 96 9C FA DD 03 A5 F4 0E
 CE F9 2C 72 47 C5 60 C0 7C 6C BB BC 68 30 78 AE
 55 DA A6 87 ED 95 93 F8 9E 80 07 E6 42 69 B7 B7
 EA D9 C6 60 BF 9B 91 75 AB 79 F4 C3 0C FF 93 FF
 F5 95 5E DF 2C FD 99 C3 F6 68 A0 75 0A BD F6 67
 06 6F 99 9C 67 7D 84 5E F1 64 FC BC 1F 37 70 39
 79 B3 26 58 C6 88 C0 96 41 65 FD 78 7A 35 24 2A
 A2 37 E3 17 8C 37 E0 C3 16 34 81 0E E7 87 30 BA
 2A 3A CE 06 C5 23 C1 F0 A2 AA 37 FC 6E 72 B7 E3
 2C C5 C8 3C 8F 0E 95 23 A9 CF B1 0C 52 A8 99 52
 A7 1F BE 21 EE 49 D5 B8 B7 D2 BD 48 A6 F5 C6 11
 3A 3A 77 0F 5D 9D D8 77 69 A9 40 9F 8D 53 40 32
 FB D8 79 A8 70 D1 0B 23 DA 52 CD 4F 8D AF CA 7E
 A2 90 3B DB 80 D9 25 5B 69 73 B7 82 FE CF 17 9A
 92 49 F7 A5 69 7F ED 77 C0 B3 DF AF AF 3D CC 1E
 06 41 19 A6 3F 06 67 DC A4 30 8A 0A 9D 2D 2B 95
 CC 9A 67 3C 72 4A 1E 78 A9 DD F0 68 DA 3E 96 33
 EE 62 52 1A A5 AB 9F 1E 2E 1A 2D 84 56 BB CB 96
 E5 A3 B7 03 FC E3 13 9B 09 E9 1B 54 99 18 E4 5B
 9A E7 D8 60 67 4F B1 AC 5D 62 0E 48 B5 40 14 AF
 43 56 40 23 A6 45 CD B3 9F 3B 90 98 67 E7 FD 4C
 0E B9 11 BC F4 E7 B8 B3 EC 31 B9 3C 0A 84 D5 28
 EC 97 DB C9 43 97 C2 43 F6 83 AB 53 99 35 08 F8
 36 14 8C 86 DF AA 7B 28 5B AD 29 A0 CC 20 A9 AC
 62 80 10 52 F1 63 17 0A 8B 99 9B EF F4 50 BE 6C
 DA 91 6F 84 14 CF 4A 32 DC 44 9A 5A 08 23 CD 72
 33 B4 B0 EE 18 4A F0 AA 6A E1 C4 FB 7E A8 A0 91
 78 9D 9E 4B B9 23 06 BC F8 A5 1E EE 2D 74 5E C7
 A4 9F 1C 2D C6 1E 20 AA 19 8E 80 85 7B 86 FA 97
 02 DC 04 F9 E8 62 96 BB F4 78 C0 F8 02 09 EA 79
 7D 55 C9 97 48 25 D1 C1 03 1A 75 F1 0F 61 46 AC
 D1 D2 41 EB 2D 7A 76 14 3E 8C B1 A9 08 36 9E 1E
 A5 A7 7E B7 21 81 AB 0F 79 7C 6D D5 7B 7F 8D FA
 64 C5 91 5E 55 FA 54 7D 65 41 6A BD 3B B7 F4 F1
 27 ED E0 73 B2 A2 C6 15 B5 1C 81 2E BE C7 0A 8A
 97 09 A2 CE EA 59 55 A7 94 01 C2 B3 A4 E7 F5 1E
 64 5E 4E 70 98 AB B2 F5 51 31 64 99 D6 48 B4 AB
 A9 0E 08 33 03 BC E2 5C 17 5C 8D B2 D6 05 E9 31
 FF A3 63 6F D3 2E 81 B7 B5 32 92 20 65 74 93 17
 77 FA 7B 1C AE 5B 76 38 42 C5 F9 5B 0D CD C1 25
 66 A4 76 A0 5C 89 35 8A DA 60 9B 56 85 0B 2A 03
 0E 07 8F D6 CE 7B F3 16 9E 63 C2 8C B1 93 BC D4
 55 F5 69 06 06 7E 56 85 DD A9 59 E2 AA 47 8C 22
 C1 93 AB 55 02 A6 87 75 E5 C9 C7 78 5B 81 02 B8
 F4 55 42 4B 7E 88 D0 1A 6E 40 D1 4A A9 DB 2C 17
 B9 16 70 9B A3 C4 15 64 1B FF 77 7B DC 41 BD 42
 D6 23 74 42 02 40 D3 C5 6C 7B 84 A9 81 8E 59 4E
 B1 79 9B 23 78 4B 56 2D 77 BF 86 1F A0 99 F1 07
 4D 51 48 37 7C E4 7A 34 45 90 27 AA 34 0A 22 0F
 4E DB B1 6D 02 86 DB A1 39 B6 69 05 D7 FE 12 03
 39 6F E0 81 35 27 B2 42 4D 96 C5 4F 20 EF 47 22
 64 6B 2E F3 EE 72 BC 0F 81 61 10 D6 55 4F FA 01
 EE 5D 6A A1 C0 3F 88 4F EA 22 86 44 7C 10 B5 7A
 76 A7 EF AD AA 84 78 1D 22 2F 89 84 E2 1E FD EE
 BE 56 64 AE A0 86 1B 69 A6 8B F8 50 AF E2 F2 DC
 CA 4D 10 37 BE C2 C8 6B 5C 08 CB 10 BC 3F 57 E2
 03 ED 67 8C 77 79 69 85 1F F6 47 10 DB 25 49 17
 FE 15 36 51 7A 68 4C 25 69 9A B7 C8 73 6F 11 33
 F9 A4 78 F0 6C FD 72 24 76 42 88 A8 2C D6 54 7C
 02 C9 37 54 CF D3 84 B0 91 E1 BE 46 70 3D 67 5F
 CD 38 8F D0 90 9B 3D 49 4F EF 2D E6 E2 87 3C 47
 03 98 00 12 17 D8 90 C5 B1 C6 31 9D 10 DC BD 5D
 BB B8 F2 BF 8A EF 39 5E FF D9 4A DF 56 79 B7 12
 C7 C2 8E 11 14 F5 AA 39 57 6B 1C F5 99 DA E4 CF
 49 6F B2 14 B6 96 CD 6C 5C 94 2E B1 08 F0 B3 54
 C3 8A 9A FE C4 AB D0 DF DD 36 FD A8 35 AD DF 7C
 83 B7 A9 7D 45 C7 5B 79 EB 74 56 22 D8 CE 18 02
 9E 44 5C 34 8B 37 89 E5 11 8B 77 E9 24 B2 92 0C
 A9 00 24 30 53 33 58 DC 38 57 95 AA 1D 7D AC AF
 F7 30 F4 78 74 78 8F BF EF BC 94 0D F8 33 76 C4
 DD 10 AC DF B2 82 87 BA 96 44 3D F4 F2 18 6D A3
 38 18 04 35 F9 A4 F1 B0 5B DE 3E 14 0D 2A E6 57
 7C 7A BE 9B 92 D2 09 4A 8B 36 69 6C CA 24 F1 F4
 D8 16 A0 C8 A9 05 80 C5 E8 A2 03 F5 05 0D E1 98
 15 DA 67 00 BA F0 C9 7E AF E2 1D 30 26 FA 03 62
 4F 19 E9 12 F5 E9 61 E2 FF 7A CF F3 E7 04 46 F7
 7C 45 32 14 BF AD 7E 59 90 41 11 C9 E0 78 4C 85
 FA 17 04 65 E0 D8 AB 01 D2 B3 D4 6F 4A 0E 15 06
 5A B2 E6 EC F0 60 2F 00 37 06 B7 30 59 F6 6F 3E
 6F BD E8 CB 2A EE 11 EB 48 55 8D 9F 14 D2 22 CA
 B3 22 5F EF 21 DE 45 4D 7D 1C 6C AD D6 5E 1B B8
 4B D4 66 5E E1 B0 FC A0 44 5B 19 02 88 AE 19 8A
 D3 3A 2A D3 13 3C AF 64 CF 4D 23 4C 6D 3C 30 9D
 24 A7 9F 9C 2C A6 31 D1 A5 4E 11 F4 C0 6A 97 A2
 D7 78 61 A9 CD DA D1 3B 1D 28 15 6C D3 10 4A 49
 A0 34 33 E6 B5 90 03 AE A0 4A D6 9B 23 0B B3 0E
 7C C0 3F AC 9F 42 D5 6C F6 11 2F 42 EF 4A 50 58
 3A 4B 16 D5 AE C3 FA E8 60 76 C7 F0 B6 3F CF 44
 09 0A 2A 12 05 DF C7 D9 6D C1 66 A0 7D EB 01 15
 C7 FE 70 EB 38 D4 68 F9 B3 03 52 4E DE A7 D5 FF
 1C D9 CC 95 16 AF 26 A4 AE EF 69 6A CD D0 0B 90
 AA 19 76 66 93 C0 4B 89 EC 26 08 7B 09 5D 74 A5
 3A 09 E7 97 9A 95 00 28 93 17 CD 44 D4 8D 78 33
 CA 37 16 28 3B F6 61 42 DE 05 7D EF 80 DE 14 4F
 7D 8F 8D 35 BA E3 A3 A2 07 0F 36 66 32 6E B6 C7
 10 E6 79 5D FE 34 51 CF BB 4A 60 E6 20 F8 11 01
 5B B7 49 8D D3 D4 31 3E EF 7F 89 66 82 45 EB 6D
 55 7E 70 B3 B5 E8 C3 75 E1 48 AF 46 09 A7 88 B8
 32 E8 21 9F D8 7A FC FF D5 6C EA EA A5 BB 15 86
 F8 E4 BA 84 87 9A 97 00 9D 3D B1 ED 46 31 D9 80
 B6 29 EF 1D 86 7E 45 E8 80 2B FA 33 12 D0 A2 95
 30 73 8A BF 1D 8F 16 5F B7 B4 CE 99 C7 B6 39 78
 54 18 5B CF B0 09 1B 8B 42 C8 90 92 9B 2F 30 97
 48 E7 BF 9A 02 6A AA 6F 6A D9 3F A3 5E 20 F9 48
 C2 77 F5 F8 5F 8C 07 63 37 3C E2 04 60 BB D3 40
 BC D6 C7 54 1D 05 28 A8 B4 C6 03 4F C0 6F 45 96
 B0 24 6D 87 42 84 1E 3A E8 8A 22 CD 5C 07 24 CF
 78 03 1B 72 FE C8 0B 14 80 54 76 B5 CF C6 A8 8C
 64 37 76 1B 0D 71 9E B0 4F 29 83 3F DE A4 8A 8F
 9D A5 8F 4F 79 31 12 00 6B AF E8 9C B8 DE DE 7E
 59 71 95 EB FA A4 75 4B 6C 17 59 4A 1A EC E7 D3
 17 C6 64 A6 01 CA 77 A1 61 1F A4 5F B6 29 F9 94
 68 50 0B 47 E6 7B FC F9 01 E2 AA 17 1C 6D 35 0E
 59 EF 36 7C 81 25 C6 D4 E8 FE F1 7E E3 28 58 18
 BC D5 0B 90 84 0D 6B D0 5C C1 27 B8 B4 DB E1 37
 59 B1 68 67 EE 5A 7A F9 35 B1 7F 3A 86 CB 07 5F
 D6 F6 52 4A 4D B2 CC 05 8D B2 11 23 2E 77 4D 43
 33 E7 17 3E 03 72 D3 FB CB EE B8 E8 A3 AD B2 61
 5E 72 F4 02 BB E2 69 C2 3E D2 91 86 AB 32 6D F2
 82 48 F5 ED 67 6B B8 D3 AC 7F 47 C4 D2 98 44 06
 B1 91 D1 46 61 11 2F 07 B6 2C D9 DF 8B DB FA D2
 ED CD BE E9 69 87 42 E3 AC 12 34 E5 D4 7D D3 EA
 39 16 D5 DB 41 60 96 D9 D5 3B C3 F7 B2 45 2E DF
 25 84 2B F8 E4 D6 2A 31 2A AA AC D4 22 07 51 D0
 C7 A6 07 22 39 CF B1 DF A3 78 B6 3C A7 AB 21 F1
 62 E0 41 E8 9A BF A1 31 96 78 64 66 2A 7E E9 CC
 2F 2C 8C 8D 39 93 F6 37 74 A4 B4 39 E1 BC E1 33
 05 1B 4E 91 68 72 54 4F 24 E9 65 7F 9D 2E 11 63
 1D C8 3A 4B 63 02 59 59 AD 74 D1 65 DA A7 48 12
 18 33 BB 01 FA BE 44 1D 6F 6E 6D 50 D1 40 56 D1
 02 D9 C9 F7 A6 32 92 A3 A5 4C DC FF 21 1C 5F 87
 F9 A4 65 D7 F6 C7 FC 7B 7F 01 8F CE BC 79 2D 00
 16 47 65 C1 8A ED C7 4C 28 0C 43 DA 6E BC 7A 6A
 96 F7 D9 D3 D5 06 52 8F 03 6F 49 40 98 5B CC D2
 B0 18 48 77 3C 46 70 CB 8F A8 49 FA 1F 66 48 99
 D6 1A 98 BC E8 FF D2 76 05 31 D6 3C 03 C1 07 39
 D0 D8 3B 39 63 B1 1B A7 C5 85 84 3C 5B CA FB DC
 C7 08 04 40 83 EA 8F 8B 3E D8 6E 82 27 34 02 5B
 F9 ED F0 91 F6 E8 48 C5 1F 69 19 E5 68 BA 37 04
 59 48 08 0F 7B A4 89 58 60 1E FD 9A 12 69 22 75
 28 0F 01 38 DF 1F D7 B8 78 40 BE 35 2A DD 96 60
 97 28 32 F1 B8 45 C4 3E E4 19 74 2F DD 7B E8 B7
 93 62 B5 85 0F 7A 46 26 4D 2A F2 EB 09 0D C6 46
 C5 35 59 6A 8D 80 E5 6F 7A D2 75 1C 05 CF F3 33
 B5 D1 6C 73 A6 1C C3 4E 64 F8 F0 10 D5 B5 64 59
 1F 4E 8A 52 90 28 8B 6D 5C 9D A4 9D E9 16 59 CE
 C0 8E AB 0A 4A F3 41 34 1E 14 A7 88 51 34 A5 30
 3E 25 03 1C B9 C3 55 52 B4 85 B8 C9 AC 43 F3 51
 AB 0A 15 EE 44 40 F4 18 49 2E 82 49 B5 53 91 20
 0E B0 FD 6F F2 82 66 13 36 18 4D 0A 11 1E 6C 30
 F9 33 66 0A BB DD AF 46 60 0B 46 5F 67 0D 9E 71
 8A D7 15 C7 E4 72 8C 77 72 D9 7D 3E 64 A2 99 28
 10 3D C3 7F 58 37 18 D8 DF 88 9A F3 4D 31 C4 A8
 8D 69 21 35 46 3C 9D 00 56 97 DC C5 EF 82 16 27
 D4 64 86 BB D5 49 28 D3 F2 45 38 60 2A 96 42 C0
 71 85 60 9C 0C 5E 28 55 66 D3 F0 62 37 E3 7B D8
 B3 1F F9 FA 87 22 F8 73 3D 24 20 FC 7C 26 82 B2
 34 2A 95 CE 4E 3B 4D 3C 36 0E 0E 6B 34 7C E1 7F
 3D 0A 48 3C 49 50 BB 02 C0 38 80 D4 18 09 59 88
 EB B0 04 9B E0 9F D8 67 A2 D9 5B 4B FA 4D 09 89
 6F CE CF 7F DE 54 8A D0 D6 07 F6 DE 32 35 E7 10
 29 36 56 CE C9 C6 9F 1D 9A 5F 84 DE 15 80 63 23
 BE A8 AF 96 AD 21 C4 25 D3 26 43 52 0E FD C8 7B
 F2 98 94 77 69 BD E0 72 AE 2F 27 2A D5 2F DA 77
 43 1A 9C 3F BE 87 AC 97 F3 B8 1E 12 AB BA B4 4D
 53 70 D6 4D 8B 93 0A 23 95 2A 0B A9 C7 33 33 55
 D6 E9 14 10 84 EC C9 E2 AC 42 74 3F 9C 1B CD 6C
 65 9D F2 92 A0 CC 63 DA 9B BE D4 25 00 57 9B 3F
 F4 3E 44 8E DB 1C 46 EA 02 3A 24 F0 F6 54 DA 14
 E4 F8 43 B4 2B 71 4C 1A 1B 8A EA C2 0E 54 AB 0D
 9E 07 2B 39 4A E6 42 E6 06 05 C1 F6 4E DA 2A 3E
 6D 44 16 8F 5C A7 BA 80 14 36 37 BF F3 C9 5F 29
 FA 55 5A 82 A0 DB E7 10 9B C1 32 19 F9 43 C7 92
 91 F5 A9 B3 D8 7B 8B 48 0C 30 D8 07 8B 3B E5 67
 55 A2 A4 D7 96 00 CA 83 42 13 E8 C4 D9 2A 83 FB
 47 D0 8A 48 BC 43 20 48 CA F0 B0 F4 3F 04 E5 D7
 F0 A4 39 2E 2C 2F 97 B9 1A 7E 53 6E D4 EF 4A B3
 BA 5D F5 0E 6E 1C 3C 93 74 A5 F8 CF D4 98 AC 9E
 FD 6D D3 16 61 44 31 CB 18 6C A9 CF A7 36 64 6B
 21 EE CB 15 29 A6 C8 FC EF 8A F4 69 52 CB F0 29
 26 37 BC A8 D3 67 9F 53 49 F8 48 8A 77 C1 3D 48
 01 D3 BA E7 D7 4D 5E 97 E7 43 08 10 AF F8 1D 4C
 86 77 6F 6A 6E 64 38 16 D7 26 1F C3 DB C0 EB E1
 B5 C1 15 91 00 3D FF FD 4A 25 3E E6 E2 03 44 BF
 58 F8 60 C9 AC 9F 25 90 7E 2B E8 E8 19 F5 14 2F
 4D 69 FA 26 12 65 0A B8 AD A4 8C 83 5F 39 B5 63
 66 A4 26 F1 FB 4A 15 12 19 F7 65 E2 61 38 0F 97
 8C BE D2 86 31 F9 83 40 C7 4B 46 96 8D DC AA B9
 B9 59 3F DB 97 5A 7E A4 44 B3 EF 36 D3 9F 95 1F
 6B F4 19 36 00 68 34 34 7A 04 63 21 84 09 81 0B
 27 B7 C7 49 49 9D A1 6D 85 A4 D7 5D 2F B0 46 CB
 B7 94 40 C0 B6 1D CB 09 42 AF EA B0 6E E4 70 44
 C2 39 7A 82 8E 68 66 FA 2A 43 73 C9 90 2B A4 40
 88 81 E4 13 0C 91 EA F0 C3 FB D1 9E 07 3B 57 EF
 82 13 26 62 51 53 59 7A 55 0E BC D4 15 A1 8E FC
 FE 74 E2 13 17 59 48 D5 08 0C 05 DE 8F 79 92 FE
 B8 34 5E 94 43 6C 39 F3 27 B7 48 09 1D B5 CE 65
 9E 45 6D ED AC 46 59 20 7A 7A 3D 21 D7 AF 13 8D
 5C 3E E2 A4 A6 58 D8 D0 9D AF 81 77 33 C4 E6 02
 6D 24 4C C8 C1 55 A3 82 E0 52 9F 33 62 41 8E CF
 2F EC 51 3A A9 F9 65 21 69 6E 57 39 28 68 88 DE
 91 E9 01 ED 4C 65 A5 3B F8 BB 6D 28 3A 8B B8 D8
 17 7A AB 64 1C 29 05 93 5F 92 D3 72 B1 1F 73 67
 99 13 DC 66 A0 ED 16 F8 9F 55 14 F7 D3 84 1A 0C
 82 49 AF AF A1 51 F6 84 A5 C4 95 62 CC 6E 6A 94
 66 93 B6 9E 83 EB E6 0A F6 E1 D8 40 E4 75 A3 B8
 08 2E 81 C7 C5 E7 C2 85 78 CE 09 22 B5 37 7A F5
 3D DB 10 35 E8 28 26 6C 7A B7 1F 99 39 5E 07 70
 A8 AA 7C B8 41 2C 9C 06 7F 8B 69 DF 83 D5 8B E6
 BA 10 8F 3F C0 81 97 68 6B 64 72 D6 B6 52 B4 6A
 67 57 3F CE 86 F3 38 26 F7 01 B8 F3 F6 CD 96 E7
 79 8F A2 B4 3B 31 38 EB B1 3A C8 CA DE 4E C2 57
 D5 EE 1E BF 7D 18 D7 8D 49 A4 20 3E 40 2D 8F 81
 39 C2 78 DB 9A FE CB F3 5F AD BC CD 7B 34 71 61
 7C 74 71 36 14 51 87 3B 02 CB 60 23 41 EC 44 9A
 1E 1F 42 62 C9 E0 A0 A9 77 5D 79 53 94 3C 05 F4
 F0 D9 8F E7 41 0E 89 96 D0 7D 4A 51 63 DC D5 6E
 A4 48 40 97 0E 2A 13 CF 9E 4A 6E 69 1B C4 89 04
 36 3F 99 07 10 B6 04 69 16 4E 22 37 15 15 6B C4
 89 22 0C F7 6E AC CE 9C DC 1B D4 74 1E 7B F1 93
 F3 4D F4 D9 6D 16 10 3B CE 87 20 F4 33 04 89 06
 A1 3B FC 62 83 1A 32 B8 5D 2D 4B AF CE 2C BA EF
 24 F2 6C 0A 5D C0 23 F7 B3 BC B8 DB 58 C8 B2 8F
 2F 27 C4 90 87 7E 41 68 10 EE D9 A0 97 1D 6B DD
 39 D2 73 45 20 2B B0 91 69 95 F9 4D FB 78 85 67
 2B A6 C7 BC C2 4B BF A9 39 72 E6 33 A6 8C 7D 2B
 9F B7 D4 8B F1 63 2D 52 6A D1 8E E3 57 D8 9E B0
 B9 CB AD 29 1C 9D 08 79 69 D6 D4 DB 1C 91 02 C1
 37 D3 AC AF 7B 40 DF 41 BB A7 6D EC CE 0E 80 F6
 82 4D C7 70 2F FB 2B 7C 6E E4 BF B4 60 8F 54 D5
 F9 B8 2D 42 77 F2 5A AC D0 38 65 C7 90 23 9E 21
 D6 B6 84 63 97 BC 18 68 C0 1E 56 47 80 56 42 77
 28 B0 7F 31 11 4D CB DF B3 5A 06 82 4A A0 1E 38
 5D F4 D4 46 6F 23 DC BA 70 37 CE 9B 12 C4 EE 7E
 D6 EB 54 E4 F8 A4 31 7C 0C A9 F8 D1 53 7C 2D F3
 E5 6C 80 F3 AD 25 C4 52 6E EF B0 AC D6 8C DB 9D
 91 60 95 B2 E3 AE 0B 4D 30 C8 29 97 6E B5 F6 05
 9D A2 D9 3D 78 27 A3 A7 7E A1 C8 A2 DD E0 BC DB
 6C 25 D2 9D 1C 48 94 CE FC F6 C9 D8 55 23 97 B2
 F4 CA BF 5D 53 0F 35 D8 7C FE FC 13 BF B5 F6 CF
 3D 1B CB CE D2 EF 38 AE 86 AE CF 64 82 C3 E0 8F
 8D 52 D9 5A 63 2D F8 C1 D4 A8 56 FD 89 D4 50 FE
 FA 14 25 D7 CD DB 6F 59 23 7F EC BF 92 86 AB 56
 3A EC 7A DC 8F A6 CA 02 F8 82 09 BF 50 3A CA 86
 B4 B5 60 BA 44 6B 2E 65 6F 6C 09 ED 04 BD 07 14
 05 5B E8 C8 40 8A 76 37 E4 B8 AC 07 9C 53 E7 62
 24 0A 11 11 9B C2 64 64 B5 60 00 D9 83 53 5F DE
 4F 97 72 64 AE 98 4B F8 7C 6F 33 B1 DC ED 3B 03
 F5 2A 57 60 60 14 44 6A E5 87 76 72 B7 85 96 4F
 8C 59 9E 93 B8 FA 7A 07 CE D0 5D ED 17 D1 8A B5
 73 2A 79 B7 F8 FF BF 70 7E E5 D5 89 F9 AB BC 4F
 02 EA C4 D9 6C 15 7E E7 D3 90 37 79 7A 5D 0A BE
 56 F4 D5 BF 14 0A 33 F3 AA C1 F1 57 7C DE 0D 52
 D1 5C 13 A0 AB 7E AA E6 1D 41 60 1B 46 24 B8 B9
 64 87 03 42 81 31 53 77 36 D4 09 36 02 3A E3 4E
 2A 28 6E B3 F0 A3 0E 9D 4F 1B C6 8D 24 74 81 9F
 BF A8 39 68 0F D4 1A 41 7C 49 C6 E9 24 A3 3D 3F
 72 82 29 1B 70 BA 5F B4 D5 9C C4 03 1C F2 8D C9
 77 CF 6D 9E 2E 28 83 2A E4 2A E4 C1 B8 21 14 DD
 76 D8 0D 64 0F 86 B9 B5 14 2B 91 32 9A B9 AF E2
 14 9B DE 61 3F 0C 17 51 9D B9 40 FE 48 5C FC 97
 6F F4 EA D7 98 4C E0 C1 64 07 80 8B CD D5 E3 31
 64 A6 F7 6E DD C7 35 A6 CD 3A 73 D3 D2 7B D6 7F
 79 CB EC 90 8A 0A DE 52 10 F8 60 0F 42 69 78 AB
 C5 3D C5 90 C5 D0 59 88 23 AF 80 CE 62 CE B8 11
 0D 72 FE CC F8 01 84 AE 70 D1 B6 F3 05 07 67 45
 E6 78 13 E2 D0 5C 8D 30 AF 7A DF E4 C5 D3 71 EC
 50 09 89 F0 42 09 3B 20 06 34 23 19 00 07 29 07
 F6 00 31 64 90 64 EA BC 09 D1 C0 A0 51 7D 2F 96
 53 33 32 3B FC 8B B4 0F A1 54 E1 AA 4F 18 57 34
 E2 71 4B 51 65 B8 F4 AE 4A 5F B8 69 1C 57 21 59
 F9 FF 3E F7 10 AC C1 D9 43 BE 32 C0 E5 4B BC 03
 CE B0 73 D3 52 05 13 34 E7 B2 45 0B 70 19 DD F0
 D0 24 D1 8C D4 2E 09 C4 A2 F1 47 F4 59 1E DF 40
 BC 8E 3B 06 05 61 E8 75 BC 2A 29 05 C7 05 B8 73
 FE CC B9 D5 AD 3D 77 15 08 B4 B9 B4 18 99 E6 13
 7F 44 11 F7 60 D0 D3 13 DB A2 CE B5 00 B2 61 79
 0F 5A 21 F5 2A 70 EE B0 EF 52 C2 96 6B 7C B4 C1
 98 72 BF 24 9E F5 45 04 DB DE A4 AA 89 7B 55 73
 F5 FC 54 08 A3 0B 48 2E 20 58 3F 22 C4 19 BC 5F
 6C 3A A4 2A 48 57 37 57 84 CD DB 32 86 5B 5D C4
 17 BC DB 5E 29 23 BE 12 80 76 24 E0 4D 34 8F 04
 98 2A 38 29 7B 24 42 32 4C 18 98 53 AA 0C EF B0
 97 23 32 C9 71 0F FC CE E3 AC 80 90 2A CE 59 5A
 3D 95 2A 0F D3 C8 78 03 80 9C 0C 94 CB 92 4C 97
 01 AA 84 47 7E CB DA B3 1D C9 E2 22 56 9E A6 E9
 A5 B8 03 8A 2C 0E E0 71 DA F0 FC 8A 96 BD DE A6
 5E 09 EC 91 6B BC DE 31 03 96 F5 62 5A A0 47 D3
 74 FA A9 3C 2A 57 C2 8C 52 F4 D3 1F 85 0B 88 87
 FB C9 A1 F4 E4 14 B6 BF F8 17 40 D9 D1 33 B3 2B
 0D 2F CA 77 C7 43 7D 4D F4 77 22 95 9F 59 2F 98
 75 1F 73 03 B8 66 7F D8 3B 51 81 D8 B1 FE E1 8C
 B8 BC 33 C4 92 72 7F CC AC F4 86 8D 1F 0F F2 75
 DB E9 81 7F E5 39 A6 E8 0D 47 16 DF FF A9 56 76
 58 F7 17 93 10 54 F0 A7 FC DD 71 54 FD 84 64 29
 A9 73 D0 C5 02 24 B8 ED 73 BE C6 28 F9 16 81 78
 2B 85 D9 01 1C F9 37 88 CB 5D 32 6E 32 F4 64 A7
 00 CE 07 6F C5 C8 FE B9 A3 4F 4A F0 4F 39 54 64
 F1 6D E7 A0 73 8D 62 63 5A A8 05 DD 5E 6A E6 42
 6A 5B 74 B9 1A 3C 83 8F 09 A3 F6 0B BD 2D 44 C1
 CE EC 46 66 86 61 87 98 13 98 2D B9 7E 8A 20 06
 C1 FB 6E E1 CD A3 10 FE 21 6E 6F 7F A8 62 D0 17
 D8 76 36 30 CE 30 37 3D 76 E5 C6 CD DB 0D D2 16
 BA 1A 09 AC DF 7B AD 73 D3 20 C2 D7 9E 25 F8 34
 01 5B C4 B7 36 F8 BC 7F C7 56 13 52 B6 0F 99 9E
 C1 8F 2F 65 24 92 8B 80 63 CA FE ED AD 84 59 B2
 CF 21 21 EA A9 C5 A2 CB 7C E9 6C D7 D5 91 B5 4D
 DA AD 20 0F 11 6F E0 44 A8 E7 B7 C3 35 1C AA 95
 8E BB 14 F2 68 53 F8 E6 B9 27 32 08 16 95 0E 6B
 6A D6 1A 78 46 70 F3 60 78 96 AD B4 EB 79 63 44
 CF 70 A8 C2 25 A1 41 82 27 AE F6 5A A7 31 46 09
 74 60 26 E5 7A 02 54 BF BF 02 F5 76 04 2F E0 97
 B0 7A 8A 85 7E 16 80 DC FE 1D C8 45 75 6C 3A 63
 02 A9 4B F3 0D E0 43 10 9A 46 64 6B CB E1 98 88
 3C 3E 3C 00 AD 4A 4A 2C 10 0E 38 61 94 65 E4 23
 33 10 9A 0C 03 8A 66 37 8B 3C 79 B1 C5 0A 13 48
 2D 92 4D D5 8F 81 16 60 C6 54 49 BD 3E 18 5E 8D
 A5 9A 47 D2 F1 CD 88 44 56 C0 0E E0 F3 DD 93 9D
 11 F1 24 10 F9 94 40 2B 2A 4E CF 2C FB 4F 61 2B
 AB 69 36 69 9D 3A 91 43 7C BB 13 28 43 7F 70 B8
 90 D4 1F BD 93 87 FA 01 A1 6F F6 E9 4D 09 CB 57
 06 7D 0F 4F FA E0 7F E3 52 0D A0 AE AD DF FA F2
 27 CC 42 D1 42 82 C0 16 63 C9 93 B2 17 5B 73 06
 6A 16 94 75 0B A8 03 F2 84 D2 75 EC 62 17 ED AF
 55 33 20 28 71 63 5A E7 AC BB DA 96 FF 67 8D 27
 8D D9 DB 33 C9 3C 2B BE CA 84 8F 6A 2D 41 C1 AA
 3B 43 B8 79 B3 C4 05 01 35 FC 05 BD F5 9C 7C 95
 D8 F7 B7 86 0B C4 7A 30 B3 52 27 40 CF 4E 0C 2B
 C8 44 82 1A A1 9B F3 BB F2 6E F1 1E 17 83 CC 02
 94 99 62 A7 F1 32 94 1E 5C 4F 3E E1 0A 93 15 DF
 10 D6 05 A5 6B A7 C7 C2 EE FB 6B 89 F2 02 24 25
 57 FE 96 84 C6 54 04 8E BA 69 09 EB C2 5E 12 DB
 7B B2 5A D4 C7 18 40 26 76 2B DA 70 8C AD 66 7C
 B1 7A B3 45 6B 69 B6 84 BC 94 EB 38 18 6C 2E 25
 7A 73 48 FE 84 45 41 57 05 8B 0F A1 E4 1B A7 63
 14 FE 58 77 F9 39 DC 66 93 3F 92 47 00 DA 52 C1
 40 5B 97 C4 C3 23 3E 1E 61 0A 1F B2 F0 57 A8 EF
 B8 4B 60 98 13 8C 01 06 43 61 17 D1 09 8F 87 05
 21 CA CA 8E 68 FC 3F 29 43 C9 99 47 FD 98 18 A8
 8B 92 20 AD 7C 64 75 1B 8F 7C B4 E3 AF DF A3 25
 D0 2D B6 5C FE 3A 9E BF 76 02 A6 2D 0C 68 77 CE
 A7 19 F0 55 05 18 0F 36 80 5A 71 47 91 FB D7 F7
 02 4E 80 41 88 90 A2 FE 5C 27 77 0C EE D3 61 C6
 40 B6 A5 28 1B DD 2C E5 19 59 C5 AE 05 C9 F0 5C
 C9 A3 4D D1 A7 5D 3E 3B 70 F7 AC 64 8B EB A4 A7
 20 6C 64 52 10 A1 CF D6 6F CB 44 A2 A6 46 C2 75
 CE FE 3C 16 25 D4 F7 1B 4E F0 E5 5E 1B AE 02 F2
 FD D4 8B 59 A0 19 89 D6 25 E6 7A 1F 79 89 A6 19
 A3 6D 96 B6 87 C2 40 F6 47 CD AB 49 5F AC CB A5
 FD 2F F7 D4 1D 8C 2B 34 9F 4B 8E EA 82 27 B2 71
 96 E5 90 0B BE 1B A8 73 F4 DD 47 E4 3B 0A 2C A2
 EF A7 BB B2 8B B9 99 0A D2 75 27 62 C3 25 2D E6
 4F 62 70 1A 2E 30 B3 2C 01 29 42 F1 BE 18 29 CB
 57 74 B0 2E 5D CC 9F 50 DB 8F 01 B1 D0 5A 37 4D
 A5 6F 5B BA D7 9D 25 62 79 DA 16 D8 1A C3 A8 47
 B9 7F 4B B0 E2 21 99 FF 7B 25 D7 3D FE 77 F3 C8
 0A 79 B8 70 41 7A 41 7F 19 E7 B7 48 A0 66 08 7B
 8A D1 86 C9 D7 67 95 C4 4F 91 CD 7C 20 FA 73 EB
 40 C1 E9 F1 80 4F 7C 48 E0 D9 8F 71 0C 5D 5D 6A
 B8 76 A3 F5 53 0F DA 89 21 C4 05 5B 64 B2 B4 01
 97 59 6F B9 80 D4 3B 24 E7 53 AF 49 5B B5 23 DD
 A4 41 84 F9 CE C3 CD B7 65 59 1A 5E 9D 3D 4F 51
 25 7E 4B CD C6 A5 40 00 D2 7E 2B B9 6D 50 CF 17
 12 9C 41 24 7D 7B D6 6D 90 ED 80 6E 3F 6F 81 43
 6A 5D DD 43 99 56 C2 1F 1F AD C8 67 82 90 6D 26
 CE 90 88 D9 68 74 4E E5 8A 6A 74 65 DC 66 56 DD
 38 4C 81 B0 7E 27 FC C1 0E 46 8B 97 C2 F6 71 99
 37 75 59 38 15 16 9A 43 37 A2 66 33 DC C9 6F CF
 3A 4F 6F EB 53 09 C1 54 BA 06 BC FE FA 6A 7B DE
 B4 2A 7C B6 0C 05 4C B9 64 42 05 3B 5D 89 98 8B
 89 EB AA 44 CD D6 D9 89 72 25 B3 A0 43 A2 97 49
 10 9A CF 86 6E 0D 80 F0 25 F8 13 F6 CC 82 18 E6
 AA 63 D1 0B 37 1C 07 C5 85 C0 2B A7 5C C8 CE 5F
 0A D1 9C 5A 38 FB 39 34 C9 1E 8F 86 01 32 EE 13
 A1 2D 16 CC CE 24 6A 04 3F C6 D6 8F 2C 0D 4A 56
 54 33 3F 69 75 32 7B BA E2 B9 74 BB D5 32 E7 49
 00 07 A5 0A AB 3E 1A 0D EA 07 E6 A4 22 BC 1B D5
 EE 6E A0 66 99 8F 50 42 C3 51 A5 85 E8 F2 2A 06
 AB 8E 65 C1 BA 47 29 50 9E E2 79 3E 94 72 DA 85
 5D EE 48 06 C9 81 87 7C 6D 77 2C 47 35 93 71 2A
 38 AC F3 04 2F 39 A9 BB F9 24 72 B0 60 86 46 58
 E0 4D 5D E9 F2 1A 81 BA 06 9D E4 B7 A7 6B A3 46
 14 18 CA B1 35 BC E5 C0 0E 4E AE 33 B7 09 6B 44
 72 F3 73 F9 DC 19 57 6C 8A 35 6D 55 47 51 AC 39
 C7 46 B4 1E C9 4D F3 71 53 DF 10 8F 2A C6 DC 61
 D4 9D B5 8F 86 FF 20 D1 E1 1C CC E7 37 5A 5D 54
 8B A5 B8 72 A9 20 32 D6 09 0F 90 68 08 9D D4 D6
 A6 93 C8 51 36 BA 82 F1 9B 9F 0E 1C B1 95 F4 FC
 D0 15 CE 5D 20 9C 01 62 C3 A6 57 6B 21 B0 34 8F
 3D ED 43 9B 26 39 42 82 25 E4 A4 11 A1 6D A3 7F
 4F 97 67 3E 95 F1 EB 5E 82 6E AE 71 28 7A 08 BC
 82 0B 05 9D 4B 48 FB 76 12 64 33 D2 88 AA AE A5
 17 C8 EE 28 5D 2A 60 24 1D 2A A3 59 E4 A3 D8 63
 15 2C 7D FC 02 53 F0 03 3C 05 67 B2 44 60 D5 34
 67 07 49 D4 EB 03 B8 1D 43 F6 DE AF C0 F8 66 47
 C6 EB AE D4 BF 7D DC 8E 46 EC 1A 01 2D 8B 00 4B
 CD BA A4 E6 43 47 3C 35 E3 79 4B 2F ED B3 AE 0F
 8E AE E9 68 58 42 37 E1 87 FD A6 94 73 95 5A F6
 29 6B 0B 6C 00 03 ED 87 95 80 AC 6C 2D D8 62 00
 F6 6D 1D 9A ED 07 B1 1A 96 34 C3 77 63 64 B6 C7
 86 D4 A6 D8 4F 37 2C 5F 60 E4 9A DC 6C F7 36 BC
 C8 48 B8 7E 40 69 E7 13 9A 1D F2 CA FC F6 5E B2
 29 81 FD 66 68 82 E5 82 F0 7C 0A FB 35 DE E6 AB
 7B 12 54 2B 7A 09 B1 7A B7 5F 86 31 37 CF D0 C3
 74 4A 1B 20 73 96 1E D9 C5 AB B6 DD 60 8F 3E 50
 FE B0 50 12 B2 65 AB AA 33 91 85 BD 35 EF 74 33
 43 3A B6 B9 70 CF A9 A4 73 2C A4 6E 31 AF D4 11
 88 DE 46 12 BA 96 5C 08 86 22 6F 6C 9C BC D4 BB
 9F 07 55 C7 0A B8 5B A3 B4 8D C1 4F 0E A6 27 EA
 B6 A5 AD 9C 55 C9 4D 0B 54 74 1B 10 02 D9 1A 07
 2A A4 E0 48 BE A9 BE 5B CD F4 DD E3 E6 EE 81 55
 DE 58 2D 82 D1 EA 25 DB 3B E5 6E 96 03 D8 2B CD
 D1 6A 32 CE 85 F9 89 0B 04 95 F5 E2 F1 C6 8B 6A
 C2 91 44 01 04 47 C6 D2 62 12 D2 80 70 DF 51 9A
 40 56 FE C3 03 2B CB 6D 91 3E 51 AA 2F 43 5D CF
 C4 D3 6C EE F8 60 70 F1 92 9A 4F 64 F5 24 CA F9
 1A EB 0D CB C4 6E E1 31 E1 9D 14 42 DD 8A DF 6E
 2C 18 03 A3 5C 40 87 9B 24 31 54 0F 79 CE C0 16
 7F 68 D6 C1 F0 96 73 5E 35 22 59 2D 86 CB 3B 8F
 78 83 D8 61 D1 DC 78 A5 BB 73 A9 4A 4A 8A 78 2B
 65 08 C7 71 1E BF C3 2D B7 92 58 98 C9 64 21 E9
 A9 C0 6E 12 A5 B0 37 C2 27 2D 21 5C 5E 48 C4 AF
 CF 3C 56 68 B7 1C AE 3A 49 93 ED 28 58 35 8B 21
 3B C6 9F B3 22 98 AE 15 F7 C6 12 AD 82 B7 D4 84
 60 85 4B BF 1A 87 FB 5F CC D9 47 E9 E6 D4 8D 1A
 95 4E BB FD 46 82 F1 60 1D 20 72 9F 2D 38 67 47
 75 85 24 7F AD DF CE 2C 41 0B A3 43 80 64 BF C4
 C1 9A 34 74 70 D6 DB 30 DB 8F 93 52 20 9A 23 C5
 3B 0A 66 90 35 0F 00 35 40 4C 2A C2 58 44 55 F9
 5F E1 4B 1A BD 26 FB 3D 70 41 D0 83 E5 70 77 43
 65 2A B4 C0 A0 74 71 C9 2D F7 F2 45 07 2F B5 B5
 7F 55 AB 66 3C AD 1B 5B 63 F7 DF 95 C5 A0 D7 B4
 0C 05 13 A0 74 AC 3D F5 94 11 6E D3 61 80 99 34
 36 D4 65 4E 0E 35 DC 5B 8A 01 A6 A9 38 29 D4 3B
 81 7C 9F 85 2A 0E 59 A0 BC 33 E5 FB 95 39 19 A8
 1F 04 AF FA 75 64 52 B7 5D 81 DD 6E B0 42 E1 C8
 C1 40 DE A8 8E 2C F9 56 D8 92 2E BF 3D 22 1E BF
 AC B1 D0 E7 D2 74 32 52 31 7D 2A D2 A3 D2 6D 23
 50 A9 1C 34 4D D9 22 FC E1 D2 AD E9 FA 09 D3 5A
 B5 06 6D F7 95 82 0B 32 A9 AF 35 A8 5C 04 83 1E
 AF C3 F5 D1 F0 DE FE B6 E9 12 11 5A 74 5B CD 1B
 6E 5F 98 71 DD 69 7F B9 71 19 F2 04 1A 71 D6 2A
 FB 49 C6 A9 36 2B 28 C8 27 B4 0F 42 9C 87 50 2F
 7B A8 D8 F9 21 6B 81 D0 44 BF 58 96 E7 F7 21 53
 63 0A 35 14 CC D8 42 86 05 3A 00 F0 91 11 0C 9D
 26 71 9C 09 8E DD 9D F4 DF 18 1A BB 2B CF CD BA
 B5 4F 5D BA 82 6F 3A 3A 6D 53 9C DD A8 56 48 B9
 73 F6 49 EC 21 9C 4D FC 46 DB 00 AE E6 4B 05 B2
 58 38 91 9A 48 F6 CF D0 B7 F1 CB E6 D1 5E ED DF
 BF 1B 14 60 B1 6B B2 01 83 F1 6F 0B 7A E7 51 A5
 03 E3 C5 BB A0 3F A2 1B 5E 6E 79 F0 2D 3D 68 40
 F2 57 99 CC 13 F6 AC 78 99 FE EE A2 D3 6C CE BC
 72 DB 03 99 94 B5 24 BB 4A 65 34 5E 8B 2B 9A E1
 A9 93 C8 9A D7 F5 1B 42 BB 2F 9B E6 EA 29 BA 74
 AB C7 3B 55 B5 41 4C B0 BD 74 D8 BD 2B 9E 46 B0
 CD 14 76 0A 43 45 15 28 AB 23 EF E8 A6 B5 2E EA
 5A E5 0F 1B E7 D6 85 E5 D8 98 3C EA B6 C0 FE 6D
 8A 8C F5 46 37 FC 6B 8F E3 43 3A 3B FA CA 55 C7
 96 F7 45 8E D2 76 25 16 71 B9 11 91 AF 9D C1 35
 18 21 FE E6 DA 96 AA 5D 44 AD 6B D8 9F D8 00 C2
 2B 33 FA 67 C7 B4 9C 91 E5 FE E5 30 35 30 C2 6B
 99 9F 56 73 5B 09 27 5B 28 0F E5 5F ED 49 65 6E
 33 45 A7 4D A9 E9 28 4A 1B 8C E7 54 BF D0 9E 3A
 76 CF AF ED 1A 7A 0E DE 9B 4F D5 5E E7 71 74 E8
 7B 98 62 3E 18 23 34 91 FF 81 FD 4A BC 65 2E C1
 CE 96 CC D6 C6 D9 EB 87 0A 5E BD 15 EB 7A C0 C0
 CA B9 93 37 C2 34 A4 6C 5E D0 41 76 7C 9A 08 22
 27 E7 04 7A D8 7F 5E 12 42 87 7F B4 29 F7 3C 93
 17 D4 D8 92 89 2B C1 76 0A 84 8D D2 C9 C0 E8 81
 26 AB A6 8D 58 66 EE 93 9D DC 00 0E A2 C3 83 71
 21 3F 2A 28 E1 92 57 E7 06 01 EB 87 18 05 27 74
 34 E7 2F 4C 52 D9 EC 5D 3B AB A9 C9 55 7F 61 45
 4E 8D 75 A5 0F C5 EB C5 9F 9B 46 6F F7 ED 0D 70
 3D 9E DA 6D 7B 5E 6E 88 F8 C0 FE B4 68 41 D0 8B
 BB 37 5A 27 35 BC A6 AE A2 DE F5 68 4C 5D 9E 13
 C3 18 3C 83 CC 5E 91 A9 FA 2D A9 79 09 34 42 E0
 BD 16 C3 10 D8 71 46 A6 A3 22 A5 5A E9 69 25 A5
 3E 1C A5 F7 20 93 5F A8 CB E6 AC A1 A2 AE 32 6F
 BC 86 A1 E6 1B 4E 0B D2 4F 22 DA 8F B7 A9 33 4E
 D9 D1 96 AF 14 1D B6 63 C8 47 EF 94 DC 10 5D 10
 30 8B FC D9 1E 0D 01 CD 64 F7 A5 11 DA FA 90 0B
 1B 1E 7C 73 F6 E3 A7 D2 8A 51 C9 48 0E 73 ED E4
 66 BC F9 E2 EE 1B 41 E0 30 EB A4 6B EA 39 6F 1C
 89 C3 56 F3 C4 69 79 D0 EF EA 4A A5 8B BD F7 0A
 B5 67 3B 00 4C AC F0 FB 8D 30 04 52 3E 7C FE AE
 2C 96 15 F5 82 91 4B 1E 24 03 04 19 D1 3C 35 BD
 06 35 31 A5 E3 4C 6C F8 D9 07 B3 10 A3 70 79 A9
 D6 46 F8 F4 E8 4C F3 4D D5 DE 96 0A C6 55 8E 79
 A9 81 6C B3 FB 0F AB F5 2E 05 85 6C 48 1C 54 24
 E0 AD AF 9B 1C D7 E9 0B 92 28 3A 47 F2 D1 70 F7
 8D 03 DC A4 B2 17 72 22 B5 FC 62 92 C2 25 72 30
 36 4D D8 06 39 20 BF D2 B6 06 3D B9 14 2B 7F 83
 FC 17 E2 AC D9 F3 25 07 A9 F4 28 7B 3C AE 90 DD
 B1 AD B5 7C 28 17 21 24 82 01 1B 8F DD 31 C1 F7
 F7 04 1B F3 23 CD 02 2E BD 86 E3 EE 24 9F 7D C3
 01 22 A7 09 8F 0C 3C 92 75 DE F3 84 59 01 3E BB
 16 7A 2D 2A 5E CD 3B 79 DB E8 38 86 21 1D 80 93
 CE 1A 28 1E 8E AE 18 33 F5 BB 53 C0 A0 98 AD A0
 CA 8B 53 22 C0 1D A8 48 89 51 7A 5A 97 95 AA 27
 57 00 1B 1D 30 F2 E2 F1 1F 9F 4C 42 CF 67 D3 57
 6D 34 D3 83 34 51 7B 4B FA 9A 43 5B CD 6A 55 E3
 CD E7 C0 72 C3 10 BD 4A 19 09 94 E1 D9 CE 4B AE
 D0 14 A8 50 30 DD 8B 59 82 6E 7B AD 3E D6 4A 8C
 E9 00 41 D9 7B EE 80 AC 17 96 63 66 B2 C5 76 D6
 D6 CB 18 20 DD 52 01 2E 97 D1 63 9A 9A 48 1F 9E
 8D 33 B0 F7 39 F3 4D 13 62 99 5D B0 8E E4 BC F9
 A6 63 25 44 9D 92 71 2A 4B 7E 08 FA 3D 82 23 8A
 4A 93 1C CE BF 52 12 D8 DD AE 99 88 67 2A 86 1F
 E0 9A F7 0E B3 8A 48 64 77 69 B8 B8 F3 99 A4 C1
 70 37 FD 11 58 00 90 BA 3C 56 7F CF 72 36 E3 D9
 9D 2C 89 E1 AD A1 81 F5 C3 96 50 17 5E CF 85 DA
 71 7D FD 2B E0 86 34 7C 22 92 E9 21 9D C7 25 86
 47 38 CB 0D 97 47 A3 33 A6 92 00 55 F3 10 2D 5F
 3A F8 34 96 7D B0 C5 70 F0 46 A7 BD 10 FD BF F6
 E3 33 50 C4 F2 F5 8E 8D 29 37 59 63 19 5D C2 80
 7C 67 48 7E F6 8F 85 5B 3A 70 C9 6C 75 34 9F 5B
 3E 1A AE B1 A0 79 3A 83 48 1C B4 CE 30 28 9A 64
 40 BC 00 BD A2 53 3E A8 48 F8 4A 8B B8 7A 2A 26
 A2 A4 65 4E 2D C3 24 F1 3B 0C B2 D7 4C D9 19 31
 1B E8 21 6D CD 3E CB 67 7B B2 03 D7 63 15 D9 E0
 50 F7 B1 0D 65 62 D4 04 FE 26 25 DC 83 47 8A 83
 23 9B C3 56 44 64 4E 90 47 4B 58 47 4F C4 1F C4
 FA 4E 3C B6 1D 32 0F 8C FB 44 81 84 2C 20 2F 39
 0F DF A6 A2 DD F0 1C DF E5 D3 B6 23 5D 1F 71 FA
 88 43 50 79 40 9C B9 3D 4F E4 6D 97 5A 52 98 C8
 68 AF 1F 17 3C E0 A0 15 BB 22 4A 6C DF 8E CF F1
 B6 33 79 1E 12 EF 34 C9 4B 43 C3 E4 97 9C B2 D4
 5C 43 A3 D9 4C 3D E5 14 40 20 6E 49 07 8A FA 35
 44 59 3C 93 28 77 FB 88 62 B8 7E 01 51 65 FD 7E
 88 DA 58 E5 8B D3 1B 24 76 E1 B7 7C 4D D6 18 99
 00 B9 43 60 F5 BD 4D 91 AC D3 F8 53 F4 54 C7 79
 A5 9F CA 24 53 79 0F 2B EC 24 47 30 C5 56 B4 48
 22 B0 8D 8B 49 BD 8F 47 0D BF 47 9D C2 13 3A CA
 F6 4A 2A 52 BA CE 7E 5E 1F 21 67 F7 AF 1D B6 24
 AC 2C 61 10 20 43 AC 9D 62 99 79 C6 84 C8 B1 58
 4D 7A 8B 2E 1C 7F D4 C7 A8 E1 48 E9 DE B4 00 CF
 18 7A 6A 0D 45 4C 85 E4 32 1F C6 C1 80 61 C8 17
 B2 32 FF 17 F7 CC 8B 29 E4 21 66 83 6F 15 66 09
 CA FB 49 69 0F D3 AF 05 66 8D 0C F7 E0 B4 F2 9B
 0B 2C 35 EC 91 3C 47 B3 AA E4 FB AA F5 B0 1A A5
 71 82 50 4B 7D 2C A1 AA E7 E7 C8 66 62 03 8E 73
 57 A6 C3 99 91 A0 E3 70 27 55 02 23 37 AA 58 12
 96 96 32 4B 11 FC 98 9E 24 B8 CC 21 F4 E7 ED 76
 2A 79 81 57 81 05 6A 59 05 63 EC FC D8 27 1F 1F
 9F 80 5D D7 36 C0 39 12 FC 13 9B 66 8A 52 72 58
 39 2D 07 B0 85 39 B3 DA 7A D5 E3 8C 18 AA 34 5E
 79 FC 63 94 8F 8B 9F 36 55 3F A0 36 CE 28 DB 77
 C3 2C 89 A6 2B BA CD 9F FA 8D 1D 9B C7 BF 58 83
 DE C7 B5 EC 57 94 3E C0 1D 0E A7 DD AB 10 08 80
 D4 AA F9 D7 6B 16 63 01 22 88 B6 9F 88 0F 3C 6A
 FC 2D 88 6C 6F DB 36 28 46 A2 E2 BC 9E 4F A6 01
 9F 77 12 B6 1B 33 BB 0F C4 31 B8 52 1B 90 C2 4E
 C0 BD 7D CF 11 8F E7 61 9E 59 F3 42 AF 98 18 E8
 7C 76 81 F0 33 9C C0 6E 06 D4 68 D3 F7 38 C2 AC
 44 C4 B7 CB 75 C0 8E 30 70 96 17 C4 6C 41 D2 A0
 E2 01 AF C7 52 60 06 55 39 E1 5A EE 3A 3C A3 E0
 FD 06 F6 19 F7 0A 7B E0 57 A6 DA 01 B8 12 7C 61
 33 4B 28 4B 3F 14 E6 C5 A0 02 5A 20 AD AB D3 0A
 31 FB 66 16 1E 68 D5 89 99 B8 3C 76 21 73 33 20
 CE A7 CA CA 42 80 A3 FC 62 28 02 91 26 59 CB CC
 66 A6 1D 5A F8 75 8A BF 5A B4 88 B2 C0 41 F0 64
 36 BB A4 46 D6 4E B4 A2 02 8F 3D CE C2 E2 AF F0
 87 EC 86 22 CF 9C 60 15 E9 EA DB 94 FC CD 82 4D
 EB 3A 53 1A A1 9E C9 15 DD 15 13 1D BA 0F D5 27
 5A 3D BB 3E EC FC 73 10 A9 3E 37 28 E6 3A 2F 0E
 A4 7C B2 3E 87 47 E5 46 62 CB 3E 9D 35 A2 3A 0E
 35 6D B7 C1 D7 CE C2 D4 D0 E4 34 44 03 29 92 19
 F0 91 81 64 E8 E5 01 A6 B5 1C 00 19 49 02 84 D3
 C0 6E 6A 2E 63 6D 99 87 02 85 D9 87 AE C4 DB 54
 52 02 F6 9B 31 B0 A8 2C 65 9A 96 47 BE BC 1F 97
 B7 03 B5 BA 92 78 7A 45 BD 26 55 94 65 45 69 25
 9B BF 1D 6B 2D 95 0E C6 71 69 B4 FE E7 EA E7 F5
 23 38 96 A5 B6 58 02 3B 74 04 B0 65 48 A8 AB 44
 47 21 F7 58 99 57 43 75 D7 E0 48 84 5D 73 B9 9E
 A2 9D 7C B0 70 FE C2 E5 DA 91 AC F6 54 AE A7 E7
 BB CA 04 DF 5E D1 22 45 8B F7 A0 90 B3 01 74 58
 C2 2B 23 14 58 EC 17 62 67 80 B4 BD E1 B6 89 1E
 84 5E EA B6 38 17 1D D9 95 DB 78 45 F2 D4 C3 26
 2B 77 EA 46 4A 09 0F 81 97 BF 51 56 51 5F F2 FB
 2B C5 6A F5 44 35 17 D7 CC C2 36 4A F6 C6 11 28
 94 9C 75 9F 09 C2 F9 E8 35 C2 F5 7C 63 DA EA AD
 98 BC 75 76 83 B7 32 09 54 BA BE E1 95 B8 97 46
 B7 30 A8 6E 5F 7B 43 09 6E B9 94 9B C3 C7 34 73
 4C 3A 95 F7 CA 62 FD D7 A7 E5 9B 04 DB DB 19 23
 7F 84 4E 48 60 B8 AF 65 72 38 10 43 1D 99 55 16
 25 06 72 A8 35 31 BE E6 E2 85 FF 67 E3 3A 1B A0
 22 76 4E 0B E1 E1 8F 73 53 CC F3 7F F9 35 67 F6
 A2 34 4C 73 19 06 99 F0 B9 CA 30 6A E1 67 BF 26
 CE C4 1C EE 86 26 82 D0 EC AB 97 17 5F AE 32 6B
 5F AA F2 C4 FB F4 E8 45 62 16 A5 B4 F9 FE A7 90
 3B D6 14 45 20 29 14 CA 94 93 DF 60 80 24 AC DC
 A2 C0 D3 BE 39 9D B9 89 84 7A 97 94 0C F8 43 66
 66 86 D5 2F 67 3D 1B 28 F8 AC F2 0D EA 4E 40 8A
 EB 44 93 C8 6F AE 7F DB CA 38 36 1B 30 0D 97 0D
 CF 13 E2 38 CF 25 CE C3 C9 7D A4 A2 B9 6E 9E C7
 86 0E 81 0C CB CE ED 83 2F 36 04 F2 2C A2 89 B7
 3A 92 8A 46 43 18 EF 2D 15 15 18 D2 5E 68 E9 03
 BA 47 45 F7 B5 8B E6 B1 8C 1A E1 D7 E1 3C 45 71
 92 6F 76 64 47 4F 45 EB 6F 73 1E 30 C7 82 45 0D
 A7 7A F7 4B 7D 3B 94 85 93 D7 2C 09 0B F9 EB 3A
 B5 75 F4 64 69 AA 33 1D 06 27 DA 18 0E 14 4C 84
 15 0F A3 BA 5E 78 03 2E DD 97 05 B2 A9 38 0A CB
 44 D8 A4 08 87 39 93 60 C0 28 B9 23 6F BC F9 52
 66 A8 DA AC 11 46 83 CB 7E D8 8D 5F 97 12 B3 2A
 BA FD EC B2 03 93 95 D8 69 06 4C BD 1D 71 14 08
 AB 1A AF A8 77 D3 9C B2 90 2F 70 CA 60 80 99 13
 8B 9F D5 69 45 C2 BA E2 AA AE E5 EE 47 F4 55 2C
 9B 73 CB 14 45 CF 31 E4 9F 84 05 06 DB 30 53 82
 3D 66 00 5B 88 51 0F B1 AB 2F 56 59 A2 E7 CB 61
 2C 95 11 E4 E5 C3 57 5A D8 D8 1E C0 F6 F4 76 44
 C3 21 CD B4 FF C5 D1 2A BE 89 EF F0 9B 96 CF AC
 48 2C 16 DD 25 6B 17 BA 7B 4C 21 EB 21 49 CB 4F
 DB 99 CB 5C 39 23 5F F6 D1 B0 37 94 9B 09 F1 BF
 85 02 14 EF 0F D8 99 5E B1 87 7A 25 33 43 F7 88
 32 89 92 32 6E ED 5B 1F F1 D4 D1 FD E2 A3 5E 22
 D0 FE AE A6 19 E3 A8 FF 24 0A 6E 74 7F 67 5E 42
 2A 35 88 36 4B 75 10 56 7E A2 FB AD BA 54 B1 FC
 58 8B BB 34 A1 78 42 76 E8 01 FF 0C 5D 2A 93 39
 66 F1 52 F5 73 62 71 A5 DA 17 A1 56 61 46 CF 15
 0C B5 F7 9F 3E 43 F6 15 A3 88 92 B4 C9 3C 5E 38
 A4 3A 8F 0E AB EC 4C F6 F5 0A A0 B8 28 94 47 07
 6B 50 DB D9 81 58 10 87 EB 93 51 72 EC AD C5 1C
 0B 55 34 3F 5C D7 EE AD AB CF C7 DF 0D DE E3 7C
 F8 25 72 15 D2 B4 3B E8 C0 97 F9 2F F7 0B 7B 2C
 F9 AF 31 3E E1 C7 EF 19 75 B9 69 8A CD 11 56 8D
 D4 3E 67 09 1F 63 AB CD 23 C4 3F 54 FA B7 3A 3A
 EA 60 0E 0F AA D9 4D 18 E6 7E 28 FC 48 A8 E8 B7
 88 33 30 3A F2 B5 BE 3E 2D 06 18 93 72 53 F6 9E
 9B D9 3C 7E 34 AB 2E 4C 79 1D 6E FD 12 CD 5A 77
 EC 3E 4A 4D 88 0E 0B 93 6D AD 46 26 58 A7 F2 AA
 91 AD 9F 89 BE 0A 02 D2 EF 92 87 4E 6D F7 71 65
 6F 98 E6 6A A8 E6 29 66 28 24 87 D0 7C 24 C5 8F
 F8 68 51 2C B8 AF 6D BD BE EF B3 F7 D1 5C 2C 6B
 B2 54 4A A0 22 4C 0A DC 52 2B B5 BC 88 9D 61 3F
 AB 25 A7 DB 68 4D 0E 3B 6C 34 CE B5 7A 1E B9 47
 F0 6D F8 AC 74 6D 87 07 81 6E E8 02 D6 BE 12 6F
 BB 7D EA 40 A6 1A EE 5E E8 14 22 94 C3 7C D8 CA
 FE A4 C6 C7 EC 4D 13 8C E0 97 06 88 45 1E EA CA
 B5 A8 76 B2 33 CC 57 E2 8F B1 69 77 18 A0 8C 74
 46 E5 8E 84 93 FD 3F A0 F1 14 13 88 20 39 CA C5
 6E AC E6 55 39 4C 1E 05 3F 66 D3 C7 10 8C 62 47
 72 C9 CD AB 9C E9 4E FD EC 4A 6E 0D 4C C0 3D EF
 97 57 95 62 09 A5 67 D8 74 12 F8 D8 73 67 CB E8
 05 19 39 81 3E 3B 14 7C B8 71 91 22 C1 AE 1C 34
 8E 15 80 E2 3E C2 19 EC B8 6A EF 2E 5A 53 31 C8
 C7 68 9B 1E F3 BF EC B7 E5 86 E9 0C 02 E8 C8 F8
 8B 3F 8D 86 DE 7E C1 0B 1C 43 E7 31 48 9A FD 52
 51 14 DE 2C 71 55 34 E8 6B 1C 1E D0 68 55 59 A5
 BA B9 BE CD 3E 07 F4 CE C0 EC C2 E8 9C BC 04 74
 91 18 41 90 C5 59 10 C5 8C F1 79 42 95 15 5B E2
 FD 46 04 68 21 56 B6 CB BA 24 BA D4 9E 74 C3 AD
 C7 AA F7 32 F6 7E 7F B8 4B E8 1F 19 5E 6B 1E D1
 06 D8 D4 8A 44 06 8D 20 50 C0 6A 96 21 0C 88 25
 B6 C6 00 7D 07 6D EB CB 84 5F 5E E8 60 EE 04 56
 72 74 B2 5C FA 4B 00 FB E8 09 89 75 57 1C 19 4D
 E0 44 95 1F A3 93 5E AB 10 F4 72 1A 52 31 97 3F
 AE D6 4A EC 5D 93 AA 81 0A 10 C0 7F 08 19 33 DD
 28 BD D6 13 BE ED 8D 28 D8 D2 E0 62 7E 52 70 B8
 25 22 EC 9D C9 B4 A3 29 5A FB 85 52 79 39 C5 98
 C2 29 AE 46 D8 0D 73 EB 66 E9 FF 33 D4 2C 77 E8
 1A 76 BF 74 2C 7E 7A 89 B2 8E 73 84 D3 EF 82 1E
 73 E9 47 54 F1 BE B0 6E B4 4A 1B 35 1F DA 79 FD
 50 9C 07 94 3B AF D4 B3 6C C2 30 D9 46 CA C6 F8
 D8 11 36 81 4A 37 E7 D5 50 FD 1A B4 E7 C0 19 52
 36 23 52 84 8E 9F F2 12 E0 CA E7 D5 38 6D CE 96
 C8 91 00 0D BF CF 06 15 8E B1 FA A8 24 AD E7 1C
 77 38 2A 28 4C 69 6C B3 24 60 7F E4 D3 B6 AE 2C
 48 22 8A 1E 9F 5D 44 72 76 C9 B5 6E 25 1B 4D BD
 E7 0E ED B6 A9 F1 C6 83 03 91 E8 3E EA D2 FA 4D
 A1 3E 90 39 EA F0 C1 F2 D2 89 0A AB 63 E0 23 70
 48 DA 36 28 6E 0C 51 EE 93 65 39 AF 7E D0 B3 B0
 73 24 8B 60 EE 61 5C A2 90 FD 07 F7 69 5E F3 64
 C9 B9 37 E6 C8 2D 13 74 EB FC AA 9D 78 8E 8D 30
 CA 0D E4 17 D5 7D 3A C5 FE 01 B2 63 6E C0 79 64
 DF B8 DE 80 A0 0D 6A 54 EC C3 20 8E C1 DE BE 57
 32 0A 9D FC 71 83 3C D8 D3 34 A1 AE 15 9A 15 B1
 1E 53 16 0B 56 C9 B9 DD 35 84 6A 58 4F BB E2 36
 8E 6B A6 8E 9B E3 3A 7D 82 C2 70 66 F3 65 F7 C5
 24 0C A8 11 C2 F8 13 73 02 79 D3 C8 49 97 4F 0B
 D3 4E E1 F4 52 2E 9D F9 93 88 11 45 C1 2F BE 16
 00 7D FD 33 49 D5 74 2D 6E 4E F5 07 94 A7 3A 3F
 FF 60 85 8E EB 64 AD 47 BB 9E 82 76 FD 6D 2A 60
 F2 80 F2 82 47 12 64 F2 F7 18 B4 A6 18 8F 1D D4
 D3 E0 3C 2B 02 AF 4F E1 1A 79 95 96 0E 21 AD 67
 AE E9 91 67 B0 6A 9C 92 34 D4 A8 74 56 5A 6D 47
 2F 95 AE 44 DE 03 E6 7F 5E EF 78 77 11 03 FE FF
 94 1A A7 C5 17 52 51 60 77 9D 53 18 DB C2 0D FA
 C8 9D BE E6 39 8D C4 A5 8C 77 22 AB 38 D2 B7 BD
 EB E9 F2 E6 09 D5 0E 35 31 8A 74 56 5F 33 93 41
 C0 28 01 24 AE 55 41 77 56 68 0B 82 8A C0 6F 87
 B7 05 5A AF E8 E4 0B 17 FA 32 3B 46 9D 21 D8 12
 48 DA 12 03 CE 2C 08 93 08 10 EF 12 D2 7A F7 C4
 D7 B3 15 A0 90 28 67 B6 19 A9 23 E6 DD 93 8A FE
 7E 50 62 9E AC B4 81 65 F5 C4 8C 60 20 94 E1 D3
 A4 35 56 C6 74 A0 CE 72 D2 9C D1 D5 EC 2C 1A 49
 53 27 46 92 3E D4 6A 3B A4 93 DB 84 11 0E E9 88
 EC 16 B5 18 DC 72 C1 BA BE EF D5 DE 1E 8B 98 D4
 C6 86 87 BE 1C DB 15 D7 6F 37 0A 51 CA F2 F7 11
 0D D7 C2 6A 77 5E 74 E5 B4 B8 44 2F 54 6C 88 DA
 BA 0D 5E BC F6 E5 F0 47 C0 E7 A7 BB 6C E8 D2 D4
 8E B2 0A 12 B1 6D 41 26 E1 61 53 05 C1 02 14 DA
 D1 B6 A5 61 85 46 DC E2 29 FF 28 63 76 04 E6 BC
 6D 55 3B BB 7F 57 8A 21 11 D9 AD 2C B8 F3 36 00
 0A DC 4F A1 12 DF 58 FD 1A 70 49 A3 A6 70 DB 3E
 1A 0E DE CD ED 30 6F 95 C4 7A C0 89 97 F4 E5 09
 33 00 50 5C D4 99 2C 67 62 E0 FD AE 52 EA DD 84
 41 FB 3A 2C 44 D2 22 72 8D 35 91 3C 90 A6 2A 41
 C8 8E 9C CA 8A 08 BE 64 F6 F2 D5 DF 2D A1 00 E3
 28 8F 45 FF 74 54 84 93 08 9A 67 4D 05 A6 5A D2
 00 A0 6F 03 C2 0D F0 85 3F C8 71 2F 8A 59 C1 2D
 17 7F CB 61 CC B3 91 5C E4 99 C0 DD 94 65 41 79
 2C C3 61 CF B3 FF 1F 54 F8 32 38 1E 06 2F 0D E5
 51 2A 08 08 F9 35 48 94 4F 63 4A 64 44 16 4C 88
 E4 F9 CE 8E 63 6D ED 21 0E 6D 5B BC 0A 82 0D B4
 F1 9B CB 0A 8D 82 9C B1 A7 FE 9C 4C B9 3C 8C 4C
 71 4D 2B B0 6D 83 93 50 68 20 F7 DC E0 AE 1B 3C
 57 D2 B6 A7 93 B0 8E F9 C8 04 78 84 C5 55 EF 3A
 FF D4 BF 9E DD CB F5 F9 63 81 70 AC 99 1D 6C A2
 1C 31 18 8F EF AD 8D AF B1 4D B5 66 80 9E CF B5
 C1 40 36 BF 12 E1 6A A7 5C 84 1E 45 80 64 71 51
 38 3A AF D1 80 18 3E C7 37 80 E6 C3 C1 1E 22 E9
 28 BA 3C 20 25 38 D6 BA A4 9E 19 42 0B 37 56 93
 D8 0C E5 9C D4 8B EA A1 D3 9F D8 00 31 A0 00 14
 AC 03 CF 82 C1 C9 E9 7B 06 93 52 BE 98 E3 83 13
 D7 20 8E E6 00 F2 41 4B 50 57 60 22 33 FC 15 6D
 FE 99 87 1F 5F E0 57 E8 0A BE 78 70 01 0D 16 A6
 01 A7 EC 8C AB 33 F9 3D 08 E9 A9 E1 4D 71 B7 2C
 6E F2 D3 C6 7E 0E D7 28 EC E5 28 08 60 2F 95 E4
 75 C4 38 B8 DE 50 F0 82 DD EF 23 0B 63 2B AE 46
 63 47 3B AA F4 43 02 76 89 89 6F C4 89 CC FD 21
 B9 3F 36 15 F9 FF 66 56 7D DA 3A 61 80 D5 60 A6
 F1 96 E7 BB 63 D4 B3 B9 EC 3C 14 ED 23 DC 9F 07
 30 37 6C 99 1B 15 C1 DE E5 D5 4F 8C E4 F3 EC A9
 AB 06 60 6D C3 9C D0 11 3E 8F 8A 57 E6 C4 18 08
 1B E5 9F 29 C4 62 44 F1 14 D6 5E EA D3 AA 35 DC
 D3 22 50 4F 70 67 2D E9 45 5C 58 83 32 8B 24 68
 7E 58 4B E4 A6 8A 93 AD 50 B5 31 BA BB B2 87 2E
 67 75 5B 2F F3 8D F0 86 DF 0E 32 58 1C 3B A3 1F
 4E 6A ED 3F E5 8E 27 C3 06 47 D2 45 18 16 13 C2
 01 1C 35 86 96 73 26 D7 BD 64 FE 3B 57 55 0B A5
 BB 20 A2 4A 02 7A 00 18 B5 55 76 04 F0 93 CC 53
 1F 87 2C 92 C8 F4 B2 96 D0 7D 7A 32 FA 52 BF 5F
 32 21 70 44 39 F4 1C F9 08 51 31 1B 05 05 73 BF
 0A 17 29 61 46 39 A3 0F 8D 0D BC F7 E4 DB 55 7E
 5F C2 08 47 64 46 A8 F9 AB 4B 33 98 F6 30 E4 57
 01 3C 70 49 E2 C3 E8 44 B4 49 48 4B F6 C9 CF 73
 B4 91 3B C8 0D 10 0E 00 AC F2 4C 59 CC D4 30 AE
 FD 7F 7A D7 BB 75 4C 59 A7 2E 6E 7F D4 4C 5F 42
 EB 05 B7 43 46 A6 FE 37 34 0C F3 9C E5 A0 DF 54
 8D F1 08 0E AB BC A3 80 97 D9 96 95 4A 09 2D BF
 CE 60 DA 87 31 DC 2B 0F E3 AD 65 8E 95 2D FE 52
 9F D2 73 E8 B7 0D 0A 05 85 84 16 AC 63 94 EF 17
 1A 95 C9 8E 96 E4 BB 20 7F 94 01 1C 20 A1 58 92
 F0 72 1E A3 94 A3 CB 02 42 59 6B FB 82 2F 0D 02
 B6 AB 86 73 5D 45 E3 F5 57 76 5B E7 35 CC 4F 65
 99 14 47 80 5F 24 9C 1E 22 88 A1 8B 48 FE 48 2B
 DE DF 30 A4 2F E1 D7 26 8E F1 DD 6C 08 53 22 17
 6A 44 8E 49 09 04 91 69 9A 3E 31 19 FF F5 6E 00
 08 4A 60 85 46 A3 0C 05 A4 6D 72 44 5B 27 E0 42
 BF BC AD 14 F4 E2 6E FC C2 61 92 74 49 B2 7D CF
 93 E2 B9 1A 9D AC A6 C9 2C 4B 4A 53 D1 43 EA 58
 CA 7C 07 7E 91 74 B3 6E 9C 20 76 93 89 1C FE BF
 67 1C C8 16 8A 5C E4 98 71 D8 AE 1E 3D CB 97 79
 F3 A2 9E DA 0F CE E0 64 FF 47 F1 00 8C 4D 57 28
 E6 24 D2 A9 B9 AD 80 20 49 10 45 B7 F3 CA F2 BC
 A6 F1 09 24 FA 30 7E FE A9 22 2E 61 93 B2 4B DE
 AA CB 31 EA 58 84 19 77 84 33 77 09 EB 5B BF E0
 6F 00 25 F5 A0 E5 F0 CF 7B 90 C8 2A 2E 9C 00 C9
 C2 41 B3 11 82 48 2D C5 FD F2 A8 BE DC DC 9C 1B
 CA 53 75 42 57 CA 43 42 9E 22 FF F6 A6 2C A2 08
 5D 40 04 58 9A B3 AA 21 4E 64 1E 20 C9 C0 E5 0E
 86 ED 8E 8F C5 AD E1 1D EB FA 06 69 EA 25 6C 95
 3B F4 F0 7A C7 40 F3 7F 91 04 1A FC 20 47 43 33
 F9 2F 67 01 6C 47 1B 61 C2 AA 25 DD FB B3 4E 7B
 21 1B 8E B2 A9 B8 61 CE 5B E9 85 1F 6B 2C 00 AD
 11 EF 89 C3 8C CD 72 F5 71 C1 C3 57 37 EB 9D 92
 09 C8 01 DE 7A 92 06 43 97 72 4E 11 B7 64 AC 17
 D4 62 9C DF 45 BD CA C6 5C 7B E1 27 B5 CD 88 BC
 F7 F4 AB 52 14 7B 93 54 FC 3E 0B 4E 71 1F 9D 3F
 00 CE 2B 59 40 82 CB C8 C2 17 D3 11 71 DF 46 53
 C9 FC 1C 71 2F 83 EC 7C C4 B8 E3 99 93 90 F8 FA
 1E B5 A5 75 0E FD B7 C8 62 0D 13 C6 CC 68 E8 DD
 22 EA E6 07 9B 67 CE CB E9 4A 41 D1 9E 05 97 E8
 E9 21 11 E7 D1 5E 8A 4E B6 DA A7 46 1C 98 E2 69
 73 92 33 A5 9F 9A 11 CC 6F 9A 4A 46 7C 73 03 92
 52 C4 06 0F E0 9B 7E E3 BD EF C8 A8 E6 B8 25 69
 EB BC 83 A9 5A F9 9C F0 2E 55 45 99 45 BB 31 5A
 C3 DC E2 7E A2 BF 52 43 63 51 FE 61 7F 9F AF 23
 5A C5 17 9A 9F E6 DC EB 0A 08 2A C9 19 82 87 A0
 9E 21 AE 33 F0 FC 7F 67 51 3D AF 18 9F 44 CA C4
 0F 3E 56 9E 7C AA 4D 89 4C AC 4D 09 65 A2 13 17
 21 4D E8 C9 5D B3 4F 8D 70 89 BE B0 E4 E6 93 D5
 43 80 A2 10 E6 37 05 83 43 32 52 0F E0 C6 48 F9
 1F F6 A4 9D B7 A5 E5 39 FF 8F 4B 62 A3 66 1E D0
 B2 41 D3 C6 39 EB CC AD 20 6E E7 CD 07 C3 D9 4A
 DA 01 C9 09 E5 90 D2 C5 3C 7C 18 87 D1 DD C2 6A
 41 FC C9 D4 0C AB D1 56 AB A3 B1 9A 0F 0C B8 5C
 30 B6 31 32 0C 7E AF 94 76 8B 93 FD 65 2B 3A 8E
 C1 11 AE 8D 02 E3 48 FF 41 F5 63 91 34 72 5F BA
 36 62 AA AD DF 68 0F E8 8C 58 1D 19 60 F4 E6 EE
 3D 42 7D 9B 72 EA 7A 6A 5D 33 A8 77 0B 65 3C 34
 BA 0B 09 FF D8 AE CD CB 81 89 86 1E C6 A1 05 31
 2B E0 0D F5 FC F2 83 D7 1A 71 40 25 39 9E D8 B2
 07 87 2A 99 7F C9 7F 26 89 9E 88 4F 13 58 1F 1C
 6A E6 A1 B4 3C 6A 7F BF C9 ED F1 49 CC 8A 95 69
 1B 62 8E 6E DB 4D 19 E5 93 7A A8 08 CC 12 FC 9C
 98 41 A8 01 17 79 AC 7A A7 92 C1 1C 51 14 D0 B2
 91 0A B1 66 6E 72 A5 B7 2F 8E 65 5A 2B 07 0F 6A
 B9 C1 56 7E 8F 1B 71 8B 6E BC F6 1E 12 32 09 43
 BA F5 1D C6 A8 45 38 67 5C 3D 11 6E 23 56 3B 6D
 9F D5 9D DE 73 3E 3D 74 72 9D 16 7D F7 27 52 45
 0C 61 89 49 7F 71 D7 22 66 FA D8 C6 91 58 E4 F0
 5D F3 BD F3 5D D9 72 B9 83 86 DC F8 16 D6 EC 2A
 37 1F 89 BF F5 9F A4 D4 C5 77 80 5D C4 EC 6A 95
 52 16 98 13 76 99 5E 5D AF 9F D1 F0 DD B9 76 5C
 8F 29 E9 A7 FC E4 78 31 5F 2A F6 97 7E 3B A6 F0
 F3 5B CE 8A 19 22 F5 D4 28 3A F6 A9 03 63 71 D4
 9B D7 7B A0 36 01 22 77 F4 43 5F 67 5E 25 E2 88
 84 93 87 5B B5 B4 4B 92 FB 94 5B D4 F7 F9 F8 B2
 9C E8 03 72 5A 74 73 41 F7 A2 96 ED 93 C3 30 7C
 C5 4B FD 72 7A 31 2B 1C 17 B4 44 97 C1 81 E5 E9
 63 4F 41 C6 7F EE 54 EF F5 A1 C4 4C EB 41 B1 3D
 24 C1 30 2B 3F 66 8C 4B 0F B8 F6 7A 2C DB CC 7A
 34 99 A7 09 AB D5 17 06 1A 8D 5B CE 68 B4 B7 50
 71 5E 5C 66 27 19 05 1A DE 8F E9 E5 28 1F DB 0A
 3A 78 D7 B2 3F 29 81 8B 6E E9 ED 15 0A 5E 7A 1B
 3F 93 DB 5E A2 A6 D9 EA FF A2 47 99 E0 F0 00 A5
 71 C2 D5 B6 6A 49 C4 ED 48 A7 60 E7 6C C6 F0 AC
 86 5B 4D 41 4B 2A EA 40 0B 5F 54 6B 0F E3 21 53
 85 F8 CB 7D C8 0D 70 10 A5 E6 08 F5 87 8E DC F4
 4B A1 2B E8 41 75 6D 17 8D 7E C6 39 F9 B5 47 05
 B9 5D AC DE B3 80 69 F3 3D 33 46 C3 84 7E 27 DB
 55 8E 9D 50 23 B6 AB ED 7B AF 43 77 B7 E7 F8 2D
 00 07 B5 B3 49 74 3A 4F AC 88 17 65 F1 FB 81 CA
 58 E9 AC 07 4A 9D 06 70 5A B1 E5 83 2B 86 6B CC
 75 21 CE 78 7D 84 CD 0A 9E 12 2F FB CE 76 34 53
 E9 80 9A 3B 95 09 EE 17 39 CA 91 69 F6 E5 5D C5
 48 A5 3A 2C FD 78 28 DE EF 0F 31 F8 86 27 66 80
 1B 55 23 7D 1D 43 D1 94 2C 92 B7 42 97 69 A4 74
 AF A2 5B DE 9E 7D 0D 88 ED EE 3E 19 91 89 AA FE
 6F 62 EF 89 13 0D 56 6C 27 5F 4E 48 6C D9 EA FC
 4B D1 7D 93 7A 7A 2D 7F B9 67 AD 94 53 9F E1 A3
 BB C3 85 CE D1 54 39 C6 DC 2B 5A 52 F3 FA 53 66
 27 81 A6 D4 FA 17 39 99 DE 97 3D 6B 5C 4B 28 3C
 DA DF 72 4B E7 82 53 8A B3 62 83 AF E7 E2 D1 CE
 7D 1F 02 39 7F F7 1D BA 15 AE 68 D3 6F 23 C6 A4
 E6 4D 2F 47 3C 62 AE C5 38 96 FC B0 6D 5F 5E 19
 B7 9F 4E A5 51 D4 6D 34 DB A8 30 F9 F2 9E C7 F8
 DA C1 98 2E D3 66 96 F7 B7 F0 BC F7 82 8C 52 EF
 A9 CE 2C 30 D8 77 E8 CA F7 24 55 1C A8 84 3E 69
 3D 5C 03 1F 93 DC A9 15 79 8A 40 C5 27 65 1A DD
 29 7B D1 44 19 56 F4 B8 4F 22 31 B0 30 4F 75 FD
 B7 00 3C 76 EC 1D D6 CF 14 63 0D 7B 72 69 A1 8E
 54 B5 E7 E9 BC 3F 60 24 77 3B D2 3D 61 32 B7 B3
 2E A7 4E B5 FD 07 BC 68 F0 5B B4 AE 26 C5 7D CF
 4D 2B 3B 95 6D 06 1D 84 DE BA 0F 60 F9 73 F6 01
 48 7C 6B 3A 35 17 D4 BB 74 E3 F2 09 C2 5D 84 B3
 39 A7 42 3E 7A F7 C8 91 8B 1E 59 C4 B0 10 32 ED
 E8 F2 16 12 FB E4 A3 B3 26 7D 6C BF 6D 83 F7 3C
 33 FA F2 89 3F 42 E2 50 88 7F 4C DD 47 B2 25 EA
 8F D8 29 65 4E 38 51 EC C8 1E DD 0C 54 13 35 F6
 29 12 B6 F8 CB AB 81 DE 8C 3B FA 79 24 00 D6 C5
 7E C7 D8 D7 84 4C 0F 14 E9 B7 EE 07 8F 9B B5 4E
 38 16 48 E8 DE A0 D4 98 E1 C1 7F CF 0F 7D CA E7
 BD 65 F4 8A 66 2E 53 9D 7E 11 5A 4F 44 23 9A 42
 1A 8C 98 F5 88 6D 9B FD DF 43 26 3F E8 FA 98 5E
 25 E7 DB 19 4A B4 ED A4 2F FE EE 67 E8 69 12 DD
 E4 E0 B2 B4 F7 99 5A 8F 41 41 49 3A 90 A2 FA 4E
 52 16 78 00 62 CA 34 90 63 E1 22 39 D4 70 2F B1
 EF 27 11 E4 57 FE DB C4 C2 7C 1E 7F 1C 2C 05 9F
 F5 EB 7F B0 CD A4 30 7F 6E 78 D7 91 DD 3E 3F 39
 ED 52 26 15 C7 28 33 7F 9B 99 04 5F D3 C6 D2 EA
 5A C8 8A B7 0F 62 4B C6 E9 6C FD 32 B0 F3 E0 CF
 EE 99 B2 CD F5 99 DA EE 08 93 BC 12 CF 46 77 66
 CE 30 03 14 6B C5 B0 0C C3 B9 39 7B E4 F8 9A 62
 44 95 58 A4 8C B3 18 6D C9 4B C0 37 0E B5 5C 22
 BB C7 7B 29 9F 25 17 93 25 81 1D D6 DC F3 AA 83
 7B 3D 88 C2 0E C1 37 F2 08 E8 C9 BA D8 82 B8 3B
 80 CC 66 AF 54 2B 1F 1C D1 31 B0 DB D1 D3 7C 76
 C2 BA 76 8A CB 51 B3 C0 A1 C7 26 0F 8F 51 03 DC
 ED 48 E4 FE 76 8D 91 AD 31 0E F3 11 BB AE E8 8A
 31 E5 38 F1 CF 1B 32 B5 55 18 35 1B 9F B8 E0 50
 2C EE EB D1 C1 FD 80 DF FC 43 DB C1 79 7A 63 B1
 9E 13 76 7A BF BC 8F 3F E7 7D E2 F6 E7 3A ED 0F
 26 38 27 9E 9E EF 59 6F BD 46 AB 2D B1 67 36 B5
 0A 07 9B C7 CB B1 F8 F0 0E 38 AB 6B 7F 74 F8 DC
 7C B9 15 43 E2 9C 00 A0 24 75 B0 0B 26 24 0E EA
 73 C8 9D 44 0C 85 95 47 55 AF 21 7E 92 5F 48 0B
 5A FB 16 48 7F E7 A7 36 DF 75 B9 98 CA B9 AD 21
 43 94 E5 DD 73 A9 7E 82 C2 44 B4 B2 DB 0E 47 EC
 F8 E0 B7 33 18 6E FD 14 8F 78 7E 54 FB B0 4B 1C
 62 FC 72 8C 41 30 D2 EE 6B AB 12 36 1C 37 E5 03
 4B 67 2A E1 EB 2D 06 54 0C 97 39 09 C3 13 20 34
 3E 68 83 BA DB 3B AA 2A A2 2D C2 0C C3 6C A4 12
 19 7A 6A 5A F5 4D 68 37 A3 AB B6 CF 77 22 3B F2
 1C 26 33 58 2B 47 DA 87 C2 41 63 CC AA F3 38 F5
 3E A9 EE 47 DE 7F A8 A0 C6 36 03 64 49 74 77 E9
 9A 04 4E AB 13 A5 CC BF F2 14 BE 68 A2 6B E8 88
 81 87 A7 96 68 64 A0 16 04 31 5F 86 5F 2D B3 B1
 90 1A 41 47 A1 9D 6C C2 47 5F 65 74 74 3E AA 2A
 9A 05 D0 8B 1C 26 D5 D2 BC 89 A0 B4 34 B1 37 FB
 BA E1 2A 37 06 78 65 63 71 E6 00 89 30 B3 65 49
 49 35 62 A6 8F 05 55 2B 66 21 28 30 30 9A 80 B6
 E7 BA F7 F7 5E F0 D0 B1 5D 37 36 2F 14 22 B9 EE
 D6 56 63 6D AF 7A 5C BC 1D 5A 0B 42 98 3F 4D FD
 34 1C 6C E7 A5 FD A6 98 4C 68 E5 D7 D9 34 71 92
 92 AC 31 5E F2 16 15 70 C7 5A DE DB D2 56 48 18
 27 10 1E 9F 62 1E C5 BD 96 C6 D1 9D F2 FD 7D EB
 23 9B 1B 0B 46 3C CA 39 5A D0 27 C2 8F 53 80 3A
 27 0B 73 D5 24 BB 7A 9C CF FA F4 82 14 9F F0 9A
 BF A8 D7 E2 46 29 95 4B B4 F0 6E 65 C7 53 67 5E
 46 DC E1 F3 16 A4 9C 74 01 E6 E9 77 DD E1 CF ED
 9B 87 DC 1D 0F A8 A3 57 24 0E 60 71 12 B5 81 0A
 76 05 91 22 8D 74 5F D7 D8 A5 E0 42 5D CE EC 94
 DE C6 FE EB 7D FF 88 C2 4A 6E 40 E7 81 52 3F 9A
 1C 51 DF 73 52 BC BA 99 25 04 31 4C 3B EF 26 A8
 29 79 CE 42 C0 46 EA 4C D6 FE 2F 66 CC BF F4 43
 48 0F 8E 8F 25 47 E9 14 C7 5B 1A 00 4E DA 08 D0
 C9 77 3D 10 BD 43 68 13 A1 9E 3D AF BD 0C 37 64
 33 76 F8 80 AB AC 44 42 82 83 11 C1 C3 A6 3A CD
 48 7D 9A 4A DB 40 F3 F4 F5 8E C3 9D 14 F5 EE 2C
 48 BC 98 6C 46 C0 C3 AD E5 51 19 6C A9 36 4F 0F
 DD 9C 76 1E B4 B2 FC 2D 1C D6 26 AB 46 77 2D 50
 96 36 BD 8B 81 DA 08 83 93 09 07 E1 5D 4C C6 02
 1F 19 C3 22 EF 5F E3 74 76 17 40 F5 37 37 18 AE
 F6 13 22 32 73 63 69 4E CC A1 7E 30 3D 07 0C 3B
 CD D8 CD 41 3F 00 13 6E 44 DD 71 5A 43 D2 14 51
 9C C8 32 EC 02 38 BA 00 4F 23 BA A8 78 CA 5D 5D
 17 0D 3F 30 25 DF 37 5D 56 2A 63 54 AE 22 3A D7
 F8 8E 03 1E 21 60 9A 04 C0 C8 CF 54 50 A6 28 CE
 57 21 12 4D A4 C6 25 CE CB 97 11 7E 31 24 38 ED
 3C AE A3 32 1D 49 F8 91 F6 D5 15 93 EA 1D CC 39
 70 76 8E EA 79 8C C6 83 41 55 2D D2 8A 61 69 3C
 86 E4 5C 3A B2 79 B3 60 B7 29 2E 94 58 10 B5 1B
 4A EB D4 B7 54 77 2B AA 21 B5 05 22 DB 28 2E 6C
 36 3C 9A 29 40 78 8B 10 9D 6C 92 A8 7D 9D 97 D3
 B9 DE 91 64 76 47 1B 02 87 FD AB 97 AA 5D C2 27
 2E CB C0 B4 8A 1E AA 14 F3 81 7C 00 3D 25 D5 4D
 49 C3 98 F4 57 42 79 65 38 53 5A 2F 00 94 90 1D
 72 FE 3D 49 5C C2 EE 5C 42 39 F5 B9 B3 DA 41 29
 3E 96 D6 92 04 22 77 07 70 A4 E4 5B DE 31 85 D1
 E3 45 BA D0 16 A6 D8 C1 03 9B 65 76 5B 3C 74 D8
 AE 99 8A 75 89 72 89 E4 2B A6 46 9F 51 E0 1E 64
 5C 91 C2 CE A0 5E FE 36 17 F7 3B B2 45 86 90 D9
 12 3F 2C DE 77 A3 24 6B 18 EB 96 2C C2 3D 9F 15
 04 3B 59 C4 34 BA DE 80 F4 C7 F1 16 E0 5B 4E 92
 79 B8 73 7D 3F C6 4F B5 7A 55 4E 91 1C E7 3C 87
 A7 7D 30 0D A9 7F DD 8F 8A 90 F8 AA 0F C7 40 8A
 A7 31 B5 6E EC 71 0B C9 09 EF AD 32 34 18 39 65
 89 31 4D 86 F4 CB C6 84 3D 19 FD A7 F0 FC 1E 66
 6B 2F B2 A2 56 7A 7A 27 40 E3 90 F0 B3 E8 EE AB
 C7 61 1D 88 FC 64 DB 84 34 35 75 A5 76 9F FA 69
 B1 EE 10 D5 24 C5 B8 A3 A4 A2 BD CD E3 E1 2D C1
 2A F2 3E C6 FA E2 25 F8 CF CB 9F 17 66 84 FF 33
 6A 32 80 07 89 6B 70 DE 3A AC CF EC BF 2B 9D 4C
 77 5D 9C 23 CA 1E 4C 33 50 4B 35 FD 0F 50 A9 7A
 43 37 E7 91 AE 24 F0 9A FA 69 E9 63 83 54 7D 12
 A8 EA 89 F5 F6 25 2E 4B B4 C2 00 ED 67 6C 75 AC
 E2 D6 A9 49 0F 4A D8 52 EC 56 0C D5 84 75 65 67
 A6 3F 9D 32 26 4C FB 46 2A F9 33 48 36 5F B0 00
 CD 5B 4B C0 FA 85 3A E1 23 1D C6 FF 6C 17 8B B9
 F6 8E 35 BC F1 94 D3 71 D8 21 1C 20 C7 82 6B 4F
 33 30 8D 2E CB 2F 36 1E C4 D2 CB 8E 00 96 94 09
 AA FD 16 9D 12 D3 CB E0 66 9D DC 28 73 11 9E B3
 D2 DA 5A 91 00 58 F9 2D 75 6A 31 55 2C CE 68 D0
 7D B3 9F 31 09 7D 19 87 23 35 D6 49 DB 8F 6E F5
 2B F8 AA 79 9C 03 BF 4C 18 A3 F2 17 DA 94 87 9C
 9A F5 AB EA B8 63 0A B8 7E DA 16 97 D9 2E EC EF
 4A F1 8E D2 7C 09 76 C0 07 49 B4 84 FB 29 0D 88
 26 2B F8 83 B1 03 10 BE 40 64 84 F7 A3 C9 2B 2A
 16 11 1B 37 D5 83 27 6D 8C BA F1 AF 13 00 E6 B4
 8E 95 E9 26 B9 38 F2 D6 48 83 EE CC F7 F8 C4 0C
 ED D4 C5 FC 38 42 2C FF B5 5D E5 39 EA 43 75 9C
 B3 60 C0 02 9D 21 BE 76 30 52 7A 2B 50 7D C5 35
 16 3A 19 68 1A 86 D5 22 2D C0 F4 39 99 C4 9C 3D
 45 29 8F A6 6B 30 7D FD F8 89 FA 6B BA 58 26 7F
 89 9B D5 01 7C 37 6E 7F 1E ED 38 CD 3D 07 CB BC
 63 FB A0 C0 D1 ED DB 97 F2 04 BF 70 49 C0 CD 7B
 85 E8 CB E7 21 A2 F6 DB 9F 3C 01 CC D0 13 51 14
 6B 04 A9 9F E3 8A 62 94 AC 33 A8 A3 D1 7C E4 97
 7E F9 AF C9 44 42 60 0C 4D E3 C1 92 D9 9F 0E 0D
 48 82 F8 9E C0 E3 DF 5E 04 92 6A B4 B1 76 E8 3A
 CD 50 2F 81 53 E0 43 7E B5 C5 BD BD D4 B5 2A DC
 E6 D6 D8 5C 54 20 9D 19 75 0A CA B0 60 07 A6 BC
 0D A1 BB 7A E5 8A 2E 5D E6 51 0F 9F 9E 3F 3F 44
 71 D6 52 F0 37 20 E1 8E 07 22 97 EF BF 35 BB 0A
 16 30 B5 BC 2C F3 54 CA E3 44 DD 08 7E 9C F2 41
 EB C5 0C B1 0A 49 EF 0C AC 88 06 AB FA ED 29 24
 D2 9D 4F F5 71 33 F3 29 8D CD 49 0B 8C D4 5A FA
 C2 0F B4 1E 92 28 CB CD 3F 21 D2 CC 28 AD C0 10
 F3 3B 0E 9C 70 E0 74 2D 34 5C 47 08 64 1F E9 48
 4B 02 1F F8 F0 F4 A1 22 E1 6E F7 70 08 49 2D 7C
 24 C9 AE 11 FC F0 41 BF E7 AE 5A B9 57 4A F2 4C
 89 1E 3D CE BD C2 2E D8 34 0C 08 21 BF 95 81 EA
 FC 56 53 84 26 10 48 E0 64 9D FA BC 1C 43 06 B1
 A7 4B 9A 00 DE B5 77 67 CC 31 44 9A D6 95 96 89
 F5 95 1D 0A 9D 4C 5C 04 9F DF 03 9A B8 61 18 0A
 74 01 BD 62 BE 02 B5 E9 47 FB 90 08 EC F6 77 9D
 B4 70 28 7E 60 9A CA 9C D0 96 B6 9F C6 80 B0 52
 CA 82 36 2B 94 5D 13 47 40 A8 30 11 1B 71 E8 AA
 BA B0 EA 8A B4 67 80 F5 5F F1 74 58 3F 6E D2 54
 F0 C7 DA 57 BC 6F A8 3A A6 2B 82 21 90 B4 D8 4B
 D3 DF B3 52 C6 4C 54 44 BC 81 28 70 A4 7C 1C FE
 E6 0A DB C6 0E B6 8D A2 87 C8 DE 0E 27 72 C3 33
 25 7E 5B 51 5B E3 36 2C E9 B9 C9 CB 25 E0 AF 0F
 E6 6D 87 68 8B 50 5B 4D F2 BF 25 B3 09 D6 64 D3
 34 6A 82 1D AA 30 79 34 3D 98 8D A7 30 2A DC EE
 3C C8 F9 7F 20 F0 A4 77 11 6E CF 63 FF 90 22 73
 DD 49 B2 D1 70 4B 49 DE 2F 74 8F 70 16 60 32 D1
 A8 35 0E BC 90 DB A5 1A 4E CB D5 00 6F A4 3F 80
 C5 13 26 A1 BB 73 65 8E 65 A7 58 C6 14 96 87 DF
 52 FE 28 FC 69 1E F7 C1 14 68 FE 27 41 7F 0F D1
 7B 59 CB 81 EC AD EA AD E5 2D E5 B0 10 5A 95 9E
 BA 66 F3 1D 83 AC 18 A6 D1 51 20 A2 81 BC 72 06
 8C F8 3D 1D E2 EB 72 40 ED 21 3D DD C6 29 A4 43
 AA 40 78 66 33 F8 9B 39 56 E1 98 1F 23 BE 89 4E
 5F 10 72 0E E0 6B FD 6E 14 85 05 12 AC 08 85 B7
 EE 70 7F 26 4E BE E2 13 54 78 3E 9C 80 FA 7A 58
 32 BB DA AA 07 73 27 C3 6D A3 67 FE E7 80 1F 49
 99 9F E3 D7 43 B5 22 FE 77 64 28 3F 1E 54 A5 92
 F5 BA B7 16 FF F1 39 1E 08 9F 39 A0 C5 FB 0F 6C
 BA FA 51 D7 0E E7 92 5B FA 72 3D 59 FF D1 9A FD
 58 74 2F F3 AD 07 C7 55 27 D8 33 10 45 3C 29 70
 F2 D0 0A CE 4D 2B 93 3B 14 36 FD D9 37 B9 D1 F7
 94 DD 78 58 DE 85 19 0A 2C CD E1 BA 0B B7 02 46
 6A 98 83 0E 63 B2 1F 69 C3 7D 98 AA DB 6D 75 F4
 A2 DA 66 A1 F7 63 9E 8B F5 19 8E 04 6C ED 50 81
 9F 05 48 03 74 06 FD B3 95 73 55 55 B3 65 A6 22
 87 CE E2 FC FB 88 D5 72 D9 35 AD 5D 29 15 22 C9
 C3 EB 69 97 B0 6D A1 F7 1F 0D 6A 43 20 BD 52 85
 D4 DF A5 7B B6 4A 4B E9 29 76 45 16 84 1D 63 94
 58 C0 5A 29 FB AC 10 72 19 9F B9 DF 26 5E C7 A6
 B5 89 C9 7F 3A A8 A2 FD AC 8D 51 8C 08 C8 1B 58
 0A A3 F0 3C 24 6E EA 4B EA 7C AE A2 20 FC 4A C0
 B2 04 CE 79 14 66 16 D0 D3 58 87 87 C7 7A D7 96
 C6 16 59 66 AF 48 4D 8A 5F 5B A7 1C 56 E5 62 47
 A5 DA 10 A8 0D 46 A2 C2 42 05 C4 3D 19 FC 86 98
 37 1F 98 D1 CB 92 AD C0 37 8C EA 9E 4B EF 34 AE
 E0 02 E1 C2 D1 94 32 DB 11 C9 1F 1D A7 A3 05 4E
 74 36 6F E8 17 39 54 03 4C 73 23 92 4A 21 42 26
 F2 C6 9F 04 D9 E4 A0 D8 3E AE 83 EB F0 05 64 E6
 CE 82 EA 92 74 24 79 02 9F 67 E3 25 C8 3B 99 8D
 79 3D 9E E6 B9 17 6F 80 E5 B0 E9 67 92 C3 3E D7
 DD 41 33 21 0A E6 DF 69 DE F1 DD 98 9F F5 D4 3E
 AC 75 72 72 87 BF A0 05 45 3F 19 B2 21 64 70 4F
 E4 C4 2A CD 01 4A 65 16 84 3B 7E C0 86 94 A8 CB
 EE 7C 60 84 8C C4 F4 81 16 57 1D DA 69 05 EA D6
 0A C2 5B D9 59 90 A8 6E 13 BA 1F 56 B1 EC B7 00
 F2 1B 0A EA A8 42 D2 79 98 0B DE 81 60 D2 B5 44
 8E F2 62 66 A2 1F 76 28 7E 57 DC 67 DC F5 05 D5
 CE C8 78 CE 23 DE 35 40 8C 6E 48 28 F5 AE FB E2
 1F 38 54 85 50 3F 67 AB 5C E6 FB EC 6F 74 2B 27
 07 4F 8D B9 92 E4 10 35 CE B1 49 63 2D C3 3A DB
 44 9F 1E 47 AF E7 81 5F 65 47 3F A6 46 58 C0 2B
 DA 98 55 A4 83 82 4F 5B 0E E0 49 1B 3B 7D 88 C6
 87 87 26 4B 63 A2 04 B0 D1 CE F8 EA 41 98 FD 2B
 89 4A 18 D8 CA 78 BA ED FC D6 D6 3B DC 7D 16 FF
 C8 33 4F B9 8C E3 25 79 54 55 A3 BE 52 60 EC F4
 C0 3B 6A 25 9B BB E1 36 80 94 C8 5D 42 8B 33 80
 DF 88 F2 E7 15 C6 B6 0A 01 AE 81 6C AD DC 1D 0F
 1C 55 9E BE 2C AD DB D1 A2 6D 47 49 14 37 42 A2
 FB 26 4A BF 46 63 32 14 48 1E 44 41 D0 A0 86 72
 25 83 E1 98 7B 79 2B 36 C0 83 9E 83 4C 3D 70 8C
 FE 53 F4 CD D0 72 C2 D7 A5 DB D6 3C 52 3B 5A 1E
 36 ED 9A 8A CE 04 4D 78 30 37 A2 C2 81 AC 52 46
 E5 22 C2 6E 8C 45 7C 2A E4 F3 38 ED 96 C6 47 93
 D3 A2 F4 D3 33 93 C0 D8 2B B5 F2 91 76 C4 C5 4E
 55 74 69 06 BF 3C A2 E0 D3 A5 52 AA AB 76 A8 C0
 FC 5F E4 4A 31 B6 5A D3 30 14 54 7F 47 DF A0 0E
 4E 15 DF 90 B4 31 69 4B D4 8B B5 86 72 BA 11 CD
 76 64 03 97 51 7A 05 2D 36 D8 9F 74 D8 60 1D 7B
 15 16 0B DD 1B 53 CB E0 36 DD 8F 60 27 03 CB 63
 AF CD 2F D9 1E 99 43 64 F8 D5 5B C4 BC 95 20 9C
 5A 9C D5 8B C5 13 50 82 24 C9 12 70 0E A2 CC 9D
 21 FE 25 C4 11 9A 3B 59 65 A1 71 B3 DD F6 EB 8F
 82 01 83 BE C5 70 79 08 DB 62 02 B8 5D D2 BF 15
 56 56 ED 16 77 CC 3E 58 E7 BD E4 E2 89 84 E5 17
 38 DE 16 6A A9 DF 1A 02 D8 C6 80 10 72 CE 5A 1A
 6E 5E A5 47 41 E7 79 D5 6E 55 FF EE AD 1E 97 3D
 0D 37 36 C9 3A D6 19 A0 D1 8C 58 7F 44 5E C1 06
 CA 56 E0 B6 A2 61 53 FC 2E D5 04 D8 90 46 08 B0
 55 26 E5 5A F9 74 96 88 B3 68 CF FF 59 9C 6A 98
 6B 0E 7A D1 95 61 41 37 1C 88 58 8E FC FD 43 2B
 EE E2 6E 51 89 26 8A 9E 3B 62 A3 0A F5 92 23 AF
 DD EE 68 7A A8 BE FB 28 F6 90 7C 03 26 6F 2E 1A
 C2 19 8C 9D 4E 22 87 18 09 55 71 96 7A D5 A9 77
 C5 DE CE 69 5F DB 88 A5 39 16 6B 54 57 00 B0 0A
 D5 55 70 5D 32 74 BB 1E 35 8D 98 FC 17 FF 72 D7
 2F 98 42 1C 08 6C E4 89 37 A5 9B 0A 76 A6 95 9A
 E5 78 40 83 F5 44 F1 E3 F8 2D 8F A3 4C 9C 3F 51
 0E 50 A5 D2 E1 C5 C1 4A 46 CD CD 32 64 B6 C9 5C
 A1 EC 9A 3E D3 66 67 13 D9 E2 C8 5B C4 62 2D 03
 FA CD E4 15 78 37 FD 66 37 DD B9 A1 F0 56 5F 14
 01 07 17 0D 6D 1A 54 B1 00 60 A9 A9 24 DA BD 19
 19 84 D6 0B 87 29 E9 85 05 4A 20 32 4E C8 FC B6
 D6 D3 EA 16 E1 B9 0B 64 69 FB A1 52 11 D5 F2 85
 0D C6 6A 4E CD AA 02 1F 69 A1 D8 6C 44 A6 F0 FD
 45 53 46 88 0B CA D9 D2 4F 7A 6E 2A 88 C5 BC C8
 A4 9F C3 56 2D 4C 9A DA 99 5D DB 58 23 E6 8D 86
 5A AF 41 39 74 C8 CB B8 B2 29 EB B3 25 FA DF 0A
 DF 21 DF F9 57 9B A3 D6 50 29 C6 5D 60 C5 98 93
 F8 5E 78 25 43 1B 5A 75 5C 2C EA 5B 18 35 4D CC
 5B 19 37 C0 E2 FB 68 0D 62 87 D3 34 D4 BA 19 56
 2D 96 BD 08 2F 1D 5F 00 DE 12 18 2C 01 45 76 49
 D2 C0 C2 CB 86 00 AA 67 D8 E5 68 FE 7A 2B 0C 97
 F2 42 41 A9 F9 88 35 11 7B 79 62 E9 DC FB C6 40
 58 BF 48 5E 49 BB 31 B4 35 6D 73 19 79 49 1E A2
 61 C8 A8 43 C0 D2 54 27 60 2B 2D 2A B8 32 BE 1D
 79 0A B4 7B B3 37 61 A9 E7 D8 89 67 60 69 03 44
 DB C3 37 AD 87 D0 3D EF 4E 93 85 CB EA 31 BE F0
 4E 2E A8 47 D5 5F 2D C4 F8 FE 9C F5 AD DB 6F 63
 22 9F AB F7 A2 3A 6F E4 6B 65 B8 1E 13 AD B8 B3
 C3 D4 F7 22 FF 72 FD 68 B5 D5 27 2F 37 60 4A 55
 D8 32 7D 22 A9 D6 22 78 7A B7 73 DA 17 DE 20 C4
 FE DB A6 FC 3E 4C 25 A1 26 CB 53 66 98 CD F0 A6
 F5 37 D4 8B 3C 33 3D 6B 10 7C DA 8A 0E F7 CB 63
 68 97 3C 13 F4 0C 97 CB 7E CE F7 D8 DA 0F 9D 89
 68 FA 87 7E FF 8E 51 33 FB F4 EB B1 49 18 1D 72
 C2 3E 33 B4 6B 75 D9 23 AF 47 50 15 B6 4E 9C AC
 9E 90 A1 0F 27 20 4E 02 50 3A 1C 38 90 FD 70 55
 9C 5F 21 88 97 B9 B4 DA 89 E7 A6 CC E2 1B 4F 03
 8D C2 DB 97 1A E9 99 2A 3B 02 C5 18 8D E3 66 4D
 1A 0D 66 27 07 B4 7A C1 04 40 A4 DF 32 B8 9F A2
 C8 BC F1 CE EA E8 8F F9 62 44 8E 2A 1E AF 4C EF
 96 C7 C0 CB 4F FA BD C5 C0 3B EC 7E 5A 7E 2E 65
 A1 27 65 37 B3 33 20 58 05 E6 A2 65 39 F9 C0 E7
 0A 28 81 11 47 38 B1 FA 37 8C D4 74 5E FC 7A 94
 E2 D3 96 BD AF 9C 1C E7 54 D3 70 95 2B B4 0D E0
 59 DF A4 BA E8 F5 EB 72 60 CA 34 88 B0 CA D9 A0
 76 00 DC 98 72 1C 34 C6 C6 21 69 91 13 11 4C C6
 3C 7C B7 08 0F F5 D9 0A 51 0E 04 8F E2 90 17 B4
 8F 86 2F 1C 51 9E 3C 42 DD C0 DC BF AD BB B3 A1
 C1 46 9D 2F A6 56 1C 38 75 D1 06 D6 24 64 C1 7D
 0C 6F FD 3B FB E5 43 A6 2D A3 D5 0F 25 8E 25 90
 A5 F9 37 36 60 9A 9A 04 40 60 C4 C2 54 B6 69 D5
 42 A5 62 F7 AC A5 7F BC BB 46 AD 13 B9 0F 00 75
 DC 3F A2 D0 8C B5 FE 0D 7B 61 48 31 98 C8 C4 6C
 05 E7 55 BB 46 D3 68 C3 D5 79 7F 9D 91 D2 5C 33
 C4 1F B4 78 0D 8C 83 21 7A B8 A1 16 84 29 3C 04
 53 68 6C D8 C8 65 1F B3 FF B9 B6 49 77 72 4E 4A
 80 B8 30 CC 41 CC 92 0E 73 1E D2 FA 6D 27 30 E1
 9E 6A F5 85 8E AE D6 C8 D9 91 FF 8F E5 B1 F4 C8
 89 9A A9 16 36 2D 7A 42 94 E1 26 E8 B4 07 E2 2C
 92 FC BC 7F A6 E6 B6 1E 9D 07 13 40 2C B4 30 91
 4C 26 BA B3 59 B1 E5 9E 77 37 6A D9 77 DB C6 57
 5D 03 9D 0E 2E 08 C6 17 04 52 32 9C EB 8E D1 3A
 0D A1 1F 4D 74 FA CC 85 EB 4A F8 EA DA 30 9D D3
 92 AA 71 6D AC 4A 30 B0 BA F4 07 9C 29 E5 A1 71
 5C 55 AF 3A 35 05 13 BB 9F 42 CA EB D8 B6 C9 CB
 F0 2A 09 5E F9 BC 0D 46 40 33 7F DB 38 95 3F B7
 EE 0C 0E 83 2D CE 0A 05 41 C4 D0 CC 4C D4 5A 28
 19 21 11 7F E4 83 09 CC C7 78 D8 D5 02 41 C2 0E
 6D 92 FF 66 FC 70 D8 81 A4 8D 95 2A 4E 1D 76 C0
 83 AE 15 A0 13 C1 CE 31 84 3A 39 9C E6 7B 20 F3
 A1 AF 8D F8 8F C8 34 97 D3 A2 11 5B 2B 1F EB 07
 06 08 97 30 81 B8 FE FF C1 3C B6 4B 68 2F C3 07
 E1 E0 AE 0E 8E 49 5E B5 0C E5 E4 F0 C9 0C A8 75
 D1 40 EC 57 D8 15 9B 48 05 DE F3 F3 C9 04 CF C4
 82 4E 7D 43 6B A4 3A 5B B7 51 8E B3 44 CE A3 41
 BD 49 1F 08 64 51 08 D6 38 C2 17 F8 A9 64 E8 62
 7A CB 96 9C 15 87 B2 7E B4 6E BE D1 B5 6A FF 36
 69 3D 1A F2 D7 73 C0 A1 BB B1 95 0D 49 A0 A7 56
 18 91 B2 6A F2 A0 0B 08 EE 98 BB D0 40 6F B6 B7
 25 D3 C8 A3 FD ED AE CE E5 5D AA 4F 38 AF 11 B8
 7D 9C E8 3B F6 F1 2E 13 01 D5 23 43 07 48 99 C9
 35 62 44 2E D5 EA AC AD 8B 2F F7 B3 31 C4 A1 C6
 93 40 4A C5 3E DC 8F E7 3F B0 61 A2 04 25 B6 F5
 77 E5 F3 B0 89 B4 65 DB 54 16 F8 5B 38 5B D5 C8
 ED 52 75 47 76 E2 BC C3 3B E3 C2 69 09 86 B1 09
 10 1D C0 03 5C 24 D5 D8 AD D9 DD 18 0C BE 92 A0
 E8 D2 92 F2 64 AD D0 24 8F 6A AE E7 5A 93 9D 3B
 22 1A 53 D4 69 D4 F9 95 9C A0 AB 70 91 E7 72 1E
 EB 40 DC 06 15 50 2B 9C 2D 9B 5C 5B A9 ED 56 DA
 62 38 6C CC B9 66 42 1B 51 0B 98 41 FB D8 05 7C
 CD BD 02 A6 BA B3 9F 09 C1 C2 55 67 1E 60 09 36
 10 97 60 84 76 65 0D 93 97 61 AA 7E 51 41 BC D4
 77 A2 1E 3F BA 58 FF 47 19 51 6A EA 34 52 58 45
 80 34 BA C3 18 E9 D1 6C 67 1A BE 5C F4 94 17 97
 1D 6F A6 2F AC 7B 7F 06 C0 5E 0F 35 7D A3 01 71
 6A 64 F5 54 E9 48 A7 B0 77 A6 B0 39 07 5A 6C FB
 BF F8 D2 DD 18 CC EB 69 67 A2 BF 43 04 91 7F FB
 E7 A8 00 BD 6E 11 C2 D8 7F 6B 12 02 C3 24 88 B3
 1E 22 66 EC 50 78 A2 47 0D 72 99 11 F0 03 C2 C1
 22 B4 C6 F1 D7 6C 9D B6 2C 65 5F 2D 3E D3 16 B4
 70 29 A3 38 57 7D C7 3B E0 ED 42 24 0A 5F 1E B6
 F7 1A EF F9 87 B9 AA 00 79 A4 D6 3F 65 AA 80 0E
 20 B0 C0 A3 4E 18 04 C1 9D A1 EA A5 7E 33 15 2E
 2A 1A 87 5B FE 99 F7 AA 88 61 1E EF E5 E9 2A B1
 65 E9 DC 1E 05 B5 A2 56 21 FC 2C FE 54 67 22 67
 55 1C E5 1B 55 D2 33 68 57 6A 51 D0 D8 AC 18 97
 A8 4A 14 2E DC A5 3F BB 1E 59 F5 0C 10 E5 7A EE
 6B 93 1A 62 2E 4F 20 D5 A5 9B 18 6A DD 3E 1B 7D
 E6 DB FF 99 A2 A3 BE AB 6E 06 66 56 D7 20 B4 3D
 C9 7F 27 C4 67 41 3A 3F B7 2F DD 93 B7 4A 77 8C
 A5 69 C8 48 0D 11 CC DE 34 01 F2 9B 78 8E 4B BC
 43 B3 D0 5F 7F 40 6A B7 9D 51 29 92 19 05 16 02
 BA 9F 48 F4 17 48 3E 1B 84 69 7D 8F 10 4F 6B 93
 79 DC 4A 34 DF 52 5B A2 AA A7 EC 36 61 1E E7 02
 DF 18 4C 61 8D 36 05 E7 26 B2 71 3B 76 62 A7 1E
 11 B0 5F DC DB 56 2C 88 FB 03 DC F5 BC F8 E0 94
 D5 93 79 9E 3C 91 FB C6 04 21 9F DD 94 9E 0F 8B
 03 AB 71 0A 5E 15 E8 76 F3 01 42 6E 7A F2 8C 6A
 43 EB 95 51 74 99 44 5C 9F 88 E3 BD A4 FD D9 CB
 2F BE F7 54 2B E1 7B C6 37 C2 AB 7C FE 91 9C B4
 50 4A 0A A7 8D 09 8C E6 25 06 F0 0C D3 DD 34 7B
 DE BF B2 C1 3E 2D B5 F7 25 C9 BE 8D 79 53 D7 DB
 FE 68 01 35 BD FB 24 F7 32 CB 7F 01 57 D7 FE F6
 11 DE E8 92 CF 09 76 30 BC 55 8D D7 91 C1 35 04
 06 1C EA CE 24 BC D2 FA 20 84 12 F6 37 74 92 93
 DE F4 F7 D6 A9 4F 2D 10 89 DE 1F 63 B4 24 DD 2A
 49 5E CC 69 E2 04 C8 5E F3 BC 96 DA E1 59 11 86
 C3 00 CF D9 52 35 64 09 D6 61 75 B2 D3 31 BC 95
 0E 93 42 1F CC E7 D5 2B 88 01 8C BA 44 89 BF 27
 A1 6A 5C 9E 36 48 CB 47 61 9F B2 32 5E 9B 9C 30
 9B 9A A3 C4 E6 F7 8D D6 10 5C AE 18 0C 65 9D A7
 D1 FF DA EB 1E 48 40 7C 4A 0C 99 DD 76 CC 37 3D
 04 9A 49 93 04 AF 7D 30 12 07 05 35 73 11 F3 55
 71 CD 1D 03 9E 00 A5 92 0A F4 AD 45 9A 49 C3 F6
 AA 30 E3 8F 78 84 C7 2A 79 59 0A 97 10 C6 0A B3
 9F A4 C8 96 9A C4 8E 7C FC 22 4E 6F C7 69 72 C6
 DA 1A B7 5C 80 4C 77 8E D0 6C 76 4A 20 D2 21 A4
 52 E3 76 8E 24 EC 18 DE B3 C9 F6 06 C8 9D 10 B2
 19 FF D2 80 6B 19 95 30 37 AA 26 58 BB 5B F3 0F
 09 2E BF EC 8B E7 51 4F 26 7C DE CD 5B 6E 05 53
 CA E1 2C 05 92 BA 80 C4 F7 A0 13 20 5C 95 E8 03
 C1 C7 6D 19 A5 26 C9 00 CC 22 15 20 DC 2F 77 AD
 4C 5F B4 C5 52 4F CF F5 31 2F D3 26 D2 F9 C2 92
 4E F8 E0 48 33 FC 60 D1 1C 13 ED 64 76 85 4B 75
 B8 EC F0 CC 00 31 1F 0D D2 D7 44 4E 07 EB F0 D7
 27 EE 32 D1 75 15 0E 14 4E 26 41 AB 3B 2A 00 00
 40 E5 16 13 6B 98 26 60 39 BB 79 51 6C 2C 31 C9
 2E C2 6A C6 B7 C6 5B E7 76 83 4A 36 9F 58 F4 FD
 E6 02 2B 1B 97 1B 4B D5 E4 7D 22 30 C0 62 5A 55
 28 EE C9 3B 88 EE 2E CA EA EE E2 52 D0 51 D1 38
 0F AB DD AE 3A 58 9B 9C 92 F5 10 B6 3F 03 CC 56
 9F F1 AB 5A 4E 2B 51 4C D0 A1 87 12 55 C8 1B 38
 96 11 3F 47 88 8F D9 7B 8E 4B D1 D1 1E 7B 0C B8
 07 57 9E 09 70 4E 00 CA 85 9B 7A 23 7A 35 22 2E
 A7 3B BC 46 2C 0F FF 08 FE 20 57 BD D7 AD 3E C8
 6C 2C 77 1F E8 26 97 D5 74 B0 83 69 25 2D 00 E7
 E0 88 E4 B8 B4 1B F6 F2 9C 96 B1 60 4A F1 09 88
 65 8D 91 D7 27 4F 01 B4 86 C3 67 89 57 05 47 BB
 7B 8F 6B 3D 69 46 A8 08 FA B2 95 59 71 6A F6 2E
 6D C7 26 CD FE 9D 70 B5 2F 67 7F B7 8E 98 33 E0
 8A 3B 59 FE E8 AD C0 1C F7 24 44 BE CF 91 72 76
 D9 23 92 D7 79 41 05 4C 47 DA 6F 34 6E AF F3 58
 8A D4 6E B4 6E 8D CD 0F 15 84 5D 5B A3 5F 86 91
 4E 2F 83 6A 26 71 10 15 71 87 21 66 39 5B 01 76
 42 D4 55 DF 71 06 22 E5 5F 7C 93 F1 FA 5C 7C 5D
 05 E6 72 E0 A0 D9 A1 BE 73 67 B9 CA A7 BA E7 38
 FB DC 05 DD 53 C0 66 24 4F A5 48 BF 86 2D 86 12
 BA E2 39 4A 40 82 68 E2 B1 F5 1C 09 D3 CC 40 D5
 76 A5 67 89 22 D1 5D 8A 4E 92 10 55 B8 8B D5 71
 2C 1C FB A5 58 9C 90 D0 0D 1E A1 39 0A CB 54 46
 93 DC 0E 87 E9 47 35 B4 AC BD DD 29 B1 79 4C 76
 B7 F0 04 EC 5F 73 A7 06 DF B6 0D 67 A0 D7 A0 93
 D6 AD A3 04 AE 01 9D 02 DD EF D9 61 C0 3B 0C 55
 B8 E6 0E 58 4B 3F 1A 35 97 AA 8D 52 5E 6F 9F 79
 E2 A7 49 C4 B7 14 FF 3D DF 96 CD D5 A1 11 CA 99
 A6 2B A9 B4 10 99 61 AA 04 35 A3 49 33 DC 01 B7
 40 90 C2 33 D8 3F 8C 38 1E 80 41 68 96 C7 CE E2
 6C 69 60 1D CC AA 2E 00 BE 7A 5C FC 40 35 B1 FD
 8B 19 BF 4F 63 A9 85 87 87 5A 92 ED 59 D2 77 0E
 56 D5 25 76 C0 4B 53 3B 4B DD 8F A0 54 83 9F 74
 00 5F 7E D9 71 80 8B 17 98 4E 0C EC 40 69 DB FA
 5E 7E 64 3A AE 1F F8 CB 27 A1 BF 3D 2B 26 BF 5C
 33 01 30 3D 90 D5 2A 20 AB DA A6 A6 1D 20 F5 71
 C5 1E 99 55 8F 92 16 85 79 1F 3E 92 46 D8 09 2C
 4C F3 92 F0 07 00 CA 79 48 52 00 6D 5C DB 08 56
 D7 0B EF C4 93 87 34 C4 A1 E4 D0 30 78 91 7D 7D
 41 89 03 F1 D7 CB B1 EE 5E 7E 16 F2 0D 8B B8 11
 6E 1E D2 E0 80 F1 D5 91 BD D2 F2 B1 00 BE F6 67
 42 94 22 B7 46 0B 9E 9E 17 24 A7 48 34 DA 24 6E
 2E 79 17 A8 AE 6B C3 52 75 7D E7 B0 74 A4 4F B4
 15 09 B4 EA E2 FA DF B6 E4 03 D2 63 73 38 22 EF
 DB 04 B6 E6 09 13 87 90 C5 3A A4 AB 57 4A 73 E5
 7A 50 B5 B9 32 EA CE 9A 9B 2D 98 2F E0 71 96 B5
 19 BB 27 4D F9 D4 12 06 C3 1C 19 CC 18 7C 15 B1
 5C 5B 2F CE 57 FF 74 FC 37 49 8E 93 D3 48 F3 20
 5C 88 01 DF 82 10 19 89 DC 8A CA 41 B1 24 95 7C
 31 6A 29 99 6A C8 D6 36 3A 84 53 DF 8B BB 34 F9
 11 F3 ED A3 94 AE B0 45 05 38 C4 C3 63 5E 96 23
 0C 25 BA 36 65 D6 BC 40 07 E2 70 4C D5 48 4B B7
 0E 9B E3 A7 33 74 9F 83 DD B3 44 BA A1 F4 2C DC
 9F B7 A3 92 3A D0 EE E5 C1 EE FB 57 F0 78 70 AA
 39 A2 8D 9F BF DC 7D A1 44 34 48 4B 11 27 BC 9A
 42 91 90 8B 01 D5 94 89 1D 35 92 8B 7A EB A5 4D
 BA 4A 88 81 FF 8B 1D F0 DE 52 67 94 8B 06 AB F9
 A2 74 DA 8C DC 69 A2 04 A1 28 A1 2F 86 B6 1B 2D
 F7 ED A5 74 09 41 E8 DB DC 6E 07 BC 22 72 29 92
 69 7C 57 F3 E5 F4 30 D7 77 8E 09 AB 0E 6E 7D F0
 4D 72 4A 65 BF F3 87 5E 2C E8 DE 16 C9 67 CF 8A
 09 E2 67 D3 EB 1E 2A FC CF D3 99 DC A5 ED 3D 00
 2D C2 DD 8D 4E 9D 53 3D 7B 44 A7 28 B7 1F 74 B3
 EB 11 B5 7F 39 DB 24 77 65 7F CB 34 F2 2B 50 98
 27 0D 63 AD 65 8F 63 BE 8F C8 2C 32 99 58 FE 8F
 35 86 BE 4E 5C 73 AE FD 93 18 98 AB 18 56 B5 21
 92 7F B0 13 7A F4 E2 66 D2 9C 37 4B F7 BB 87 FF
 98 83 17 44 2F 2F DB EF 70 40 DD AA E6 0F C1 3D
 25 8D D0 FD BF 94 8D E2 71 71 58 04 2E 9D B2 8A
 A3 3E 31 93 0F E7 24 97 A4 D0 1C 72 35 44 7E C1
 80 06 57 C8 86 88 54 A8 7E 09 9C 31 C8 5B 49 E1
 8C 01 94 C1 D1 EC 31 75 B9 CD B2 C5 D5 71 72 75
 58 3C C1 F5 E5 8A 51 28 A0 E6 B8 CD A3 52 16 BF
 91 3F D2 15 89 8F E1 D8 3F 13 6E BF B4 E2 C2 8A
 2E 8D 40 CB D3 24 BE 13 08 49 AA FD 54 B2 B5 DA
 9E B9 54 A7 CD 4E DE 55 40 1D 77 CF 94 8B 16 F6
 32 27 4B 8C ED D1 C6 2D EF D9 A1 DF B0 59 35 D9
 C4 7A 4B 3E 43 36 87 BE DB F9 75 4D C9 B5 3D 79
 5B C3 69 61 78 02 94 5A 63 E8 85 09 2F 1A A3 90
 DF 63 51 14 1A 65 29 4F 38 88 11 71 1B 40 5E E5
 14 A8 E4 BE B5 03 E4 EF 35 72 7F 1D 5E 73 63 95
 0D 5F 66 3E 00 0C DE A6 A2 CD 01 84 BC E5 4E 09
 B0 82 7A A9 81 EB EC 8B 5A BD 4F FD 44 1B F7 6B
 C1 EF 2E 1B 62 FA 69 40 16 F9 EB D2 FB AB 7D F9
 1B 5B 88 67 5A DE 72 B5 97 E6 08 AD 4B 5B D2 A9
 8C 47 26 6E 31 40 DA E0 31 A9 CD B1 B0 6D 41 15
 32 9E 7E 90 31 39 B9 38 5A E3 CA BD 16 C9 E0 FF
 1E 96 CF D2 BC E6 99 8C 52 FE D9 FE 19 9E B6 EA
 9F 84 D2 0A D3 C2 36 EA E7 5E 59 ED 77 40 9E D9
 BD 69 33 73 81 AA 19 73 D4 00 FC 2B 7A B7 F3 B8
 26 AE 94 D2 6D C2 9E A7 EF 22 66 EA 59 FC 1A B5
 4B 91 39 84 4B D3 7C A0 2F 96 DB 6D 2A FE CC 9D
 CA DC BF 97 4E 4A C2 0F 42 A4 EE 3D A2 4A 82 CD
 FB D2 6E A4 01 2A F6 68 B3 AA C7 A5 F5 C8 31 51
 98 29 28 4D 69 7F C8 CF FF CB 25 98 A7 9B 05 B5
 5C 1E 28 3A DB AC B7 E3 24 70 A6 13 40 6F D6 CB
 92 9E D9 36 3F 42 24 74 9B 3C A6 65 B1 24 18 D1
 79 EE B2 ED 2A FD 56 77 CF 03 A6 85 BD B4 90 1F
 CF 38 49 BE A4 25 C3 81 16 58 AE 12 B5 A1 96 95
 B2 35 71 75 25 4C 49 0E 93 5B 04 26 B9 FA 62 33
 CA 50 DC BE 14 CF 5D 81 95 65 9D E4 AE 47 EE 24
 D2 DF D7 82 6E C5 BB D3 15 0F 5C EF E6 EA 4F CE
 19 87 42 D0 B5 7D 99 1E AD 5E B4 39 3B 91 55 04
 8E 00 36 7A 27 63 83 A7 EA 92 1C BB FA 36 23 A5
 D0 AA CE 90 AB 6A CA 15 99 56 C5 71 67 E6 EB 34
 4C 33 E7 95 29 7B A4 D8 A1 F2 66 E7 CA C5 98 67
 98 27 35 DD EA E9 97 54 2B 0B 96 CF D0 84 C8 34
 D7 C1 E0 BA 29 FB 1F 1E 08 36 93 3B AA 7A D3 C0
 74 DE 3C DD 4C A3 62 31 38 9F D6 3C 66 4C 24 4E
 3C E0 06 E9 3E F6 83 CD 35 41 1E 55 54 70 9F B9
 FA A4 2D 77 8B 85 2E D1 C0 D1 BC E0 7A 90 20 FF
 BD 42 B3 3E 5F 62 E9 DE 1E 1F 65 1C 7B B8 43 D1
 75 B9 E5 45 94 84 07 95 14 29 BB 8F A3 68 B3 64
 2F A0 99 53 37 F0 E1 F3 48 03 35 AC 9E A2 4F F6
 7F 80 FF E7 96 51 E4 42 F3 EC FC 9A 99 0F C0 55
 DF 0F 41 5B EC E4 9C 7E 29 4C 27 A9 06 5B 79 84
 20 66 9A 8A 6A 01 82 83 85 0A 59 8F 48 E7 45 64
 71 43 9C 34 B9 B1 4B 05 CD 25 15 28 4F 66 8D 4B
 EA 91 BB ED 75 56 51 67 9C 3D 49 58 16 69 52 5E
 2A 51 19 5A 5C 43 03 5D 00 A6 1B E2 F9 9C 85 73
 36 2E A2 2E 1A FA EB 79 73 09 DA 2E C4 55 B5 30
 7A A1 E7 EA 23 8A 31 7C ED BE A5 FC 95 20 E8 D2
 5F EC A5 E3 AF A2 A2 6E 89 41 73 E6 B3 46 C5 34
 DE 45 EE 80 41 C8 09 27 DC FF 33 C3 03 AE 21 41
 AE 67 88 F6 6A E6 67 E5 9F CD 49 EB B9 94 06 BF
 10 E0 99 70 48 A6 69 17 22 B9 4E D1 8F 45 06 12
 0E 72 C2 90 F5 59 D4 8D E6 C3 D4 31 1D DF 4C 17
 79 60 87 64 DE 40 AF 5B 4C C7 F9 4D 73 0E F9 7E
 34 85 54 AC C8 DE 26 56 F6 5D 37 96 2A F3 52 EC
 8F 78 FC 8F 6C 46 9B C0 E5 17 71 AB 6C 43 D8 8D
 B5 7B A7 2E 2C 04 DD 14 64 C4 98 B6 CA C9 05 05
 A9 A8 22 F1 C2 3E AB DC 0B FE 2B EE DF 88 12 24
 59 27 8F E6 E5 F8 F0 E1 F9 D4 A1 36 A1 B6 38 32
 4C C9 49 0B B2 52 18 FE 38 A6 E9 CE 29 A3 4C 90
 11 36 75 DC 98 F4 DD 13 AC D0 8A 01 E7 5D 74 8B
 58 7F 33 53 8F 7A 4C 95 DC 03 9C 95 1D 59 D7 C3
 26 5F 32 58 CC BD 4E F2 3C 07 4D BD CA 38 0C E0
 B6 31 37 13 23 1D BB A2 67 6F E9 06 0F 20 61 1E
 30 73 1E 62 05 02 3C 8A 5A 20 3D EC 67 99 64 84
 14 43 52 08 74 69 48 B6 85 B2 3E F4 97 AA 46 60
 4D 3C FF A0 5F DB 3A AB 4E B1 A8 19 B8 8F 20 77
 CC B9 BE 21 DA FC 54 4C D9 11 CF C5 FE 9D 00 94
 E0 6A 00 C8 B9 DD C9 35 FF 8D 65 49 AB 37 3A 73
 13 F5 AA 4D B1 47 07 5C 77 8D C8 54 40 55 86 0F
 6F 5E 8C 5C 7C 44 34 F3 EE 8B C6 9C 31 15 0D 25
 E7 9D D9 3B 6C 25 F5 E8 34 F5 B1 1C DD 76 C8 90
 C6 97 19 A8 BC 95 B3 D7 F5 39 63 E6 FD 58 E6 9A
 36 57 A1 68 FE 30 21 5B F5 79 E5 2A 53 65 99 D4
 67 8B 8D D1 1F 29 3E 62 25 B8 84 31 56 1B 17 D6
 49 55 5C EE 41 1D 8A 7F BF B6 95 46 41 8C BB 1A
 3D 66 EE 2E B4 13 27 5B 28 AA 46 FF 3A 7A 18 22
 8F D5 A1 78 FF DC D0 58 F3 65 A2 81 0E 03 F0 D3
 1F EE 2E 21 22 B0 E8 77 42 3C 03 38 6B 90 D4 26
 D6 1B AA 3D 4A 25 25 EF 22 F4 9A B3 9B E4 CC 2F
 57 42 0D A7 7A F0 3D 7C 43 B0 11 73 89 67 AA A3
 77 52 E4 3D 4C 3A 1A 34 40 EE 65 49 7A E8 62 12
 42 8F 5B 56 D2 18 37 D7 98 A0 A2 E6 7B 52 69 73
 5E 75 7F 24 3F C7 63 58 04 22 55 BC F3 82 4D A9
 02 C9 DF EE FE 89 51 7B 51 BD 05 62 3D B4 04 88
 EA FA 86 B4 0A 09 97 67 32 FC 69 40 C7 B4 9B 8F
 E9 55 B5 B4 F0 17 CE 9D 08 CA 1E 15 75 9D 47 5D
 75 78 B3 D2 EA 5B ED C9 68 7F 11 4F 71 17 D9 82
 8F B8 C4 47 43 63 A4 A8 C6 19 D6 EB AF 91 03 6D
 81 07 3D 28 33 29 DD 51 82 28 0C AB 74 C4 5B 74
 09 B3 6D E4 6D DD CF 9B AB 6F 5F 3A 2A EF 87 6E
 8E 69 46 38 A7 D7 79 CE FF D3 B5 97 64 2E 4D 06
 67 5E A3 39 96 E4 6A F4 58 D5 A7 29 01 F6 09 0B
 84 D9 31 CD C0 9E D9 DE EC F3 EE 21 6D B0 F1 CA
 CE 63 24 3D 39 D1 5C 2A 51 EA 08 F6 9E 90 65 D9
 D2 5B 4A 87 84 70 4D B0 72 C1 9D A8 4E D1 93 39
 21 37 3A BD 4F 80 0C 2A 10 9A C1 90 2B D3 2F AC
 DA E2 82 7F 57 E7 64 CC 4B 63 7B D8 81 6E 4E 2C
 86 84 68 13 C3 69 9A B4 CA D7 FF 0E F8 ED 79 D7
 DD 72 E6 DC 2A FE 7F A4 09 7B DA FB 24 F8 06 43
 F8 F7 D9 D3 68 C3 72 D5 B8 4A 36 E8 F9 41 22 0D
 25 44 56 A9 07 43 CE 0F FB F2 93 4F 9F 0C 42 DA
 18 A6 6C 12 0D 6C 02 4C DE 9D 72 5B 64 30 72 FF
 49 E3 F5 60 CF F6 8F BA 6C E9 4B F0 E6 A1 12 E1
 92 52 54 75 DC EE 0B 7B B4 F6 3F 48 FD EA 86 7E
 D0 8D C7 FF B9 CD 8F 8E B0 D3 84 9E C2 67 74 A0
 69 52 9C 59 41 8B 56 69 40 F5 55 49 A8 FA BD F1
 93 0E 34 E5 A0 CF 99 38 F7 79 CF C9 4D 96 C4 33
 5B E5 02 AB 43 C3 C4 AF B5 F0 E7 BB D3 B1 6C 70
 3D 37 18 49 72 DD CC 40 93 D7 82 49 2D 80 9A 66
 2C 9D 1E 09 AD 45 0C FA 79 E4 95 11 37 DD E3 E8
 23 9C 54 46 0D AC 78 10 A5 03 B6 54 5E 7C E4 83
 AE 7B 36 D3 D2 2A A2 F1 67 6C B6 50 A0 5A 87 9D
 D8 1F 6F 30 D9 3B D1 64 87 50 FA 34 02 5A 29 3F
 92 31 81 40 5A 84 25 95 64 E9 03 32 E5 3B 6E F1
 D5 42 43 46 10 F1 29 6A 6E 99 11 48 61 26 45 AD
 0C 3E 54 2C 7C 33 CB 45 00 42 1D 22 9F 1A D6 46
 BD AC BD BB 82 83 8B 7D 19 3D D3 8A 65 22 4C 9E
 E1 EC BE 8C 8F 1C DD 3D 70 56 AF AF AD 5A ED 9A
 D0 28 8C 21 A4 AB F2 3B 3E 9F 06 C6 B6 A2 2D 15
 92 3A 17 88 05 B4 32 6A 24 D6 F4 69 67 8A 65 CD
 B3 11 53 88 C1 AC 3F D8 83 CB 54 A9 F0 84 64 CF
 DA BC 5E 9F 19 B3 5D 87 29 EF 8A 42 7D 12 6D 8F
 F4 CC 2B 17 54 A7 6B A3 F7 F2 66 04 8B F5 3C 42
 C5 D4 EF 8D 10 0B 3C 23 DE 7B FA 4D B3 2F 32 DE
 4F FE 03 88 46 35 F3 E3 BB 65 E0 81 05 3A 57 C2
 DB EE 95 FD 29 E5 F2 00 85 58 AB 26 CE AF 6D 07
 FA 30 83 1C 9C 7F F9 C2 4A 90 FC 31 2B FD B1 D4
 EF 1B CD 50 7B 51 D5 78 21 BF FB A9 1F 72 22 A0
 2A 85 5D BF F7 DF 45 57 C7 DF 46 2B 93 9A 78 F2
 DA D3 56 A6 3A 7E 15 42 AC 6E 6C 01 DC 8D 17 D7
 D4 BD 04 CF E4 23 04 33 89 79 43 CA 72 0B 9A 71
 A3 BF 31 AF 4C 60 7D 2E 20 F3 81 4D F5 6C D6 41
 52 9E 8D 4B E7 FE BB 2D CE F2 98 5E E9 C8 79 DE
 27 94 BD 60 AC B6 FD 26 BF 6B A5 F2 89 32 D2 3A
 6D CF DB DA 00 F7 1C BA FA EA B3 DA 08 65 FE 6C
 BC 88 29 8D 04 04 EF 56 74 1E CA 76 A4 78 AE 07
 FB 5E 59 0A 57 88 29 F9 4B 14 50 2F 66 D5 CC 85
 30 D1 49 B2 BD 81 C3 1E BA 55 14 2C F3 B6 AF 34
 AB A7 18 F7 29 81 E2 DE 13 B0 BD 32 72 34 9D AE
 02 7F A9 FB B6 2F C7 E1 22 15 78 68 35 6A 7B 2A
 23 C8 D5 7E D4 52 E1 0D AD C2 80 4B 12 E7 C6 11
 46 98 8C 01 9F 2A 93 CF DB 95 90 77 CF C6 E3 E4
 D7 D8 D8 22 D6 F6 1D 74 4F E8 D4 5C DC 70 5D 40
 4E 92 E4 DC 17 C3 6C 0A 3F 80 B9 F0 2D AE 16 42
 F4 99 30 F4 AD 7C 9E 86 21 49 C6 E7 06 ED D1 CF
 30 8D B4 8E 1A 88 7C 75 C1 16 AE E7 77 CA 3C 1E
 CC 5A 66 59 F1 D0 64 E9 C5 18 7C 1C 2A F2 C2 6C
 20 7A 87 DC 80 76 F7 06 DE BE 4E 14 88 84 12 8D
 F3 1B 8B 2E 55 29 F6 7A 2F 19 28 98 74 AA 35 CA
 53 F7 9F B8 36 1E 55 ED 2D DC F0 2F FC D0 13 F0
 08 5F D9 94 B7 F6 E4 79 00 1B BA 43 45 FB 39 A3
 95 86 26 1D D0 D0 3F AA 5A 93 EB 50 62 7A 51 06
 06 47 F8 8C 08 59 2A E6 08 54 C5 68 B2 EF 21 F5
 BA BD 19 A9 17 45 C2 38 CF 5D BF AE 06 51 50 DD
 D3 32 72 2C BD A2 E4 7F DC 81 DD 41 08 CB ED 07
 1C 6B 8D 7D B6 C0 F4 86 F8 6F D9 35 C3 AD 59 CC
 C0 C9 FF 88 08 A6 CC B6 7B FF BA C3 10 C3 A4 5F
 C9 D8 80 D0 0C 7F 90 8A CD 92 D4 EC 14 62 34 07
 C4 CF 44 34 E3 FF 72 0E F2 4D FF D6 1A 1C E8 BA
 EC 62 D6 B7 DA A0 6C 53 A4 F0 87 01 EC 4E E7 70
 3D AA 46 B9 20 C4 EC 4D 12 26 11 14 B2 D0 5F B4
 1F 77 71 DE D5 64 65 B5 72 0D B2 99 B7 46 2C CE
 76 92 D0 D2 87 3C AC B5 2D 65 D3 C7 91 9B 55 4F
 3B FA 3F 1E D7 64 F9 BF FD F6 E2 58 D6 45 0D 67
 55 C4 B3 01 8F DE DC E8 0C A7 96 71 3A FA 98 7D
 E1 FD EE FB 46 D3 21 53 B6 1A 31 D1 61 5A 4C 2F
 5D 80 67 E4 D1 ED 85 B7 A5 AA 25 AC 61 2E BE CB
 5D EC 43 13 A5 4B DA 8B 77 0A 3F EF 06 2A AE 67
 10 B7 B4 20 53 55 0A EC 04 D7 87 7C 6D A7 15 C8
 1F 0A 77 52 3D 49 C4 9D 0E B3 E5 0D 1C B5 7D F9
 D8 0F 18 9E 7C 32 75 5C 8A FB 3E F8 4D 6A 18 AC
 EB AB 1E 35 E9 17 88 4A 32 2F 06 E1 57 BD 94 F6
 73 63 F7 A5 3D 3E 85 67 66 7F E9 1A B8 37 C6 9D
 B8 1F EA 07 1D D5 AD B4 77 D2 82 3B 1E 8F 78 66
 9F 1F 71 4F EE 9A 66 FF 84 AE 87 EB 16 8B 63 49
 3E AB 9E B8 55 89 C2 F6 8B A3 CC 29 AB 30 6F 4A
 67 8D 0F FC E8 B6 60 95 84 4A 5C FA 8F 28 C6 99
 48 52 41 7D 2C BD F8 1D 35 4D 4F 32 F4 6C 72 10
 ED D8 8A C3 8F 45 BC 01 55 BA DB F7 27 75 00 E3
 69 74 72 5B FD E0 98 D7 A4 EA 9D EE 2A 9F B4 4B
 C6 B8 93 49 01 4B 3F 8B 3A D3 EB 5C BA 11 C2 FC
 5E CC 6A C0 64 C8 13 64 9B 1E 12 9E BE FB A8 63
 8B 23 C2 5A 11 86 04 F5 28 FC 9C 9F 81 13 40 A0
 F0 BE C0 B6 87 C3 E4 EB 93 37 48 2E 3A CE C8 5C
 3F FD 99 34 BC 15 B7 9F 6B FB D0 16 1B B1 1E 95
 7F 3D 20 FF 29 3C 90 16 BE CF 1D 76 C8 BD 89 3E
 8E 51 CB 6E 41 F7 C9 41 4E C7 9B A0 78 FD B2 9D
 89 3B 06 9A 1A EA 0E D1 C6 C5 BC 16 5A 03 C0 75
 3B 9A 70 E4 68 00 16 FC 6C AE 0D DF E5 F3 E9 70
 85 AC C2 C5 FC 6B 90 45 E9 04 FE 9F 5A 16 61 3C
 04 D6 C1 1C 40 B5 AA 35 35 9E 8E 1B C7 A4 A8 E2
 3B 4A 29 1D 3B FF 8F 68 FC 06 92 00 AF E2 78 74
 CE 74 BD 13 FC 03 73 E3 99 FB FA 0C 37 1B 0C 05
 5A FD 19 43 79 E5 9B 2D E4 42 B2 DF A8 A7 2E DA
 38 D8 DC 74 A4 6B D7 1B D9 24 CA 31 27 2F 94 FF
 6D 59 F1 D4 33 F4 05 87 28 78 17 A2 D9 21 32 09
 4E FB 80 5C 79 38 D4 BF DA A8 BD 53 83 15 0F 9F
 F6 30 8D 68 7F A5 1D E3 E7 88 1E 1B 12 97 4D 6B
 48 67 8B 34 99 72 63 C8 AD 71 AF 49 45 5B BF AF
 FD 09 64 DD A4 32 E1 DD 64 70 CE 9A C4 96 37 3B
 64 42 1F 53 78 B1 EC 68 BC BF DC 82 06 FC 0B A8
 B3 1D 5A C2 08 8E 8A E5 2A AB FE 6F FE 5E 2D 3A
 D5 53 79 87 E1 49 C5 5B FA 65 AA 03 6C 82 15 30
 4B C5 47 7B B6 DE 7F 7B C9 3B 7B 90 A6 50 9A 1E
 12 0A 0D 9D EE 34 39 85 25 6A 6C DA 67 00 A7 00
 12 27 AE 4E 38 08 2B 37 BA 2F 3F A9 6D 76 49 21
 5E A3 2C C2 EF 85 C8 46 38 66 78 DB EB B1 C6 66
 B2 9B ED 8B 21 4D 98 13 01 49 C6 A7 46 CB 0F 67
 DC 44 39 D8 5A BD 6F 5F C4 22 03 D3 55 E4 DD 17
 91 FE 45 A9 38 5D 6B 9D 80 91 0B E8 CF FB 61 ED
 8E CB 31 22 7B 46 EB AA E6 17 B7 D3 74 BF 89 7B
 FA DC 50 26 97 64 7C B8 8B BC 78 AB 59 70 BA 4C
 AB 4F 7C 14 5A 3A B9 F3 F0 DD 11 58 6B BD EC 2A
 51 B4 97 32 E2 63 FB 6B 56 F9 70 78 5D 9B 1C 88
 6D 25 6B A4 1A 9C 8B B2 90 5E 56 D8 F1 09 4B B7
 5F D4 53 26 C4 4A 4D 35 57 D2 03 8E 1B AB 91 6A
 8D CA 64 12 94 18 79 7B 70 37 84 E0 F0 45 6E 67
 D4 25 5A 07 E0 A5 F3 D6 94 0F 1E B9 28 A8 15 0E
 81 36 B8 AB 69 6B AC B7 24 1E ED 6D 1F 09 A0 DC
 DE 05 10 64 F6 35 83 F8 89 AB B6 54 FC 7C C3 E9
 27 0D 27 1F 16 6F 7D 76 90 8C 46 F5 5B 40 3B E0
 32 9B 74 45 48 65 C6 CD FF 20 3D 41 91 19 73 C0
 57 75 CB 80 44 8B 2F 13 65 17 E0 EE 78 5D 83 BC
 1F 18 EC 9C 99 B3 D8 4F D3 4B A3 AB BA C8 69 8D
 00 3E 1A 2C 23 FC 02 2C 5C C8 D4 35 7A 84 1C 6E
 00 0E 59 31 46 ED 76 DC 79 18 9D D4 A0 32 C3 1E
 69 B0 2F BA B2 ED 26 1F A7 C4 F1 B1 CA BC 8A 46
 CC 14 BA C4 2B 46 96 90 0C 46 A9 B4 46 B9 6F E1
 37 2F 4F F4 F3 E6 74 59 DB EC 78 26 47 64 D3 FE
 1B 88 B6 88 F4 F0 A5 21 7D EE 0E 34 C2 00 7A D6
 94 8E 5E 26 73 5F CC 85 4A CF 42 17 0F 8F 69 96
 C9 BF 31 2F 86 D9 F1 DA EB 75 0B AD 60 3E 89 66
 16 06 F6 F7 9C 44 4C 35 2C F4 80 29 F0 34 26 B9
 16 17 1E B9 05 CD E8 DB 33 1E E1 A7 36 1B 58 D1
 F3 B0 E2 72 C2 32 19 6E CF 84 08 E5 86 7C 54 F8
 35 A0 D6 E5 96 D0 3F F2 09 F7 1D FE 51 C2 0E 14
 65 90 0F 6A F6 E9 1E 61 28 14 C7 23 D4 5B EB E8
 3E 06 54 2A FE 2B D5 6F 90 DA 95 7E 97 64 E9 C6
 47 A2 24 B8 5A 0C 10 65 CE 58 1F 1C EA 8A DC F2
 60 9D 6A 2A 25 E3 66 AE 5B DE 18 C7 01 35 87 FC
 53 C5 12 45 CF 3B D1 62 49 DC 7A FD 80 42 C3 CE
 F9 CE 98 E2 1C 4A 80 1C EC 11 F3 32 48 FB 11 A7
 4A FC 13 CD CF AA C9 8B BB 29 D9 55 40 91 99 AE
 DF 0A D2 28 48 D1 D3 85 ED FE 16 19 41 63 50 5E
 39 1B 26 BD F9 2B BC BE 04 28 19 1E 50 2B 5E AC
 27 E7 E4 7A FB 65 54 9E 10 8D 0F 69 03 C3 9F 34
 2B 31 2B 35 70 BF BB 6C 12 EE E9 81 E7 4C 98 D8
 78 C1 55 98 19 30 CB 67 AD 10 33 46 01 7F 78 4E
 1A 40 CA 7A 09 8F 3B 71 7C B1 0F 50 4F 85 2B BD
 F2 3A BD 0A D6 8F 83 34 6D A2 2C 1B EB 00 66 9D
 D2 05 FE 45 1D C4 B9 AF 41 92 75 80 3B 1F 41 A3
 E6 70 33 B3 07 FA 58 72 E6 BE 8B 10 AF A5 98 38
 A8 01 A4 0C 0B 18 45 7A 7D C8 40 A7 51 82 9F A5
 5D 3A BF 9F 17 BA CA 5E BB 4E C5 47 C5 75 46 FE
 3E 5D A2 28 DA 39 F3 DD 09 59 F9 97 2F 64 C2 0D
 65 47 14 D2 34 FF 71 B5 9C 25 F4 E3 56 36 1B E9
 E4 3E 04 6E 2F 8A E0 14 19 71 ED 23 8F 7C DA 42
 E6 52 B9 BB 17 EC BB 71 B9 DD 73 74 D6 31 ED 2E
 3C E6 9B F6 94 8F FD 27 15 A0 BD 1E A3 6B 9A 8D
 10 5C 76 AB BB CC 4D C9 AA 99 91 AC 32 57 83 D0
 9D AA 85 3B 42 2F FE AA 35 C5 B1 13 E4 E6 8D A0
 DE 65 C1 81 9D 27 EE 6B 12 6F 95 F7 A2 8C 2A C2
 8C A9 C0 25 BC 52 14 75 77 91 C4 E9 5D 25 AF 96
 53 1F CF 9A 08 EB 48 16 FF 11 19 10 F1 2D 7B 48
 16 4A 94 B7 F3 47 15 5C A6 43 41 A0 36 12 78 1B
 55 4E C1 0C F5 25 37 87 FB A5 AA E0 60 9C 2C 59
 23 E1 6B 1C FA 7D 6F BA 2F D4 0D 3F 3A 78 AA F3
 8B A0 DC AC AD 3E 90 AD 0F 79 46 89 CB D0 BF 98
 7F CC D3 14 08 7B 24 24 9E 57 67 31 59 1A 90 61
 EA A7 9E AD 67 E5 A9 FF 5B B0 89 7D 61 D9 EF 3D
 8D 24 BA 52 33 83 FC 57 60 63 07 FD 93 8D 8F EE
 EB 44 61 FC 93 0B FD C0 8C A0 07 06 CC 54 33 CD
 BE A4 9F 4E F6 65 6F CB 29 47 8F 9C F7 4D B1 6F
 2A AD 61 E9 C3 6E 19 83 95 B6 D4 E0 1B 9B 6D 44
 DA 9E 78 C0 0A A1 1E AD EE 99 13 54 C5 7D F9 22
 DC F3 08 35 67 21 76 41 FC 4B 70 B6 FC EC E1 D8
 56 8C F9 C1 C0 A3 41 E8 BB 26 B9 C5 0B D5 8B 81
 99 B2 56 E8 74 04 75 CF 7F E5 82 2C FB 7B E5 C6
 D5 46 9C 71 0F 7F B8 9F CA 70 15 B9 8D 57 00 33
 26 EA 91 28 B6 6F B2 31 63 41 8A A9 82 C8 58 6F
 29 41 F8 DE 30 86 E7 6F 0A BC BD E4 D8 9D 0E ED
 CC 70 C7 DB 5E E7 86 20 27 66 C6 E3 F3 1C 25 A9
 FD 1F 8C 65 79 17 7F A3 A9 99 19 52 FD 86 70 1C
 F1 48 50 F1 AB 39 42 BA 9C 9A 23 C1 33 27 9E 1E
 35 CA A1 17 55 F4 0C 7B 82 F2 7F C3 A5 48 53 98
 61 69 0E E8 3D 80 0F 28 63 7A DA 76 2B 2A D6 69
 01 97 DE 02 2F 84 73 AD 79 FF 21 F4 FC 23 34 62
 16 B1 F5 CA 85 B3 90 5D 58 99 83 6D 2E 56 33 B6
 7C 03 20 0B E5 78 3F 44 16 D3 ED 46 65 EC 68 A3
 48 D6 C3 AC BA D5 7B 8B F1 03 06 0E 95 B9 CD 7B
 E5 DA A1 6D 86 ED B3 52 16 9F 54 3C 2B C9 5F 6D
 67 80 86 3A 43 44 4A 04 5F AB 15 2C 33 A2 B7 92
 D2 2D 5F 39 E7 BA 80 A8 B9 B9 CD D3 1B 14 5E C3
 D3 B8 F4 CA 79 2C A0 C7 D2 28 4E 66 FE 24 50 8C
 16 59 36 4C 65 C2 D0 41 FC 38 6C CE 7F 51 4B 80
 09 2A 5F 21 35 5A 73 1D EC 09 63 A6 63 51 F2 1E
 05 F4 A4 4E E4 DE 8D DD DD 1C F7 CF A7 D1 CC B4
 A0 3B A4 69 76 D8 9F 98 2D EF 25 92 95 F7 93 02
 90 80 7D C5 04 86 16 E8 91 15 5D D5 D0 60 35 11
 4E E0 3D 7F DE 0B EC 33 C5 82 56 C8 B2 98 44 81
 C3 33 B6 E6 1A CB 04 2C 0D CE CB 79 79 CF 03 92
 9B 6D 74 9A A4 A3 22 01 F1 1A 38 B7 75 B2 D9 10
 B4 FC CF 35 DC 42 DA C0 97 DB A0 31 C7 20 2F F7
 4E 47 A7 28 42 26 38 44 06 90 5C 41 A5 13 C9 5A
 FF 93 07 E4 C2 3B B8 D7 DE 1F 4B 26 C8 59 61 36
 76 39 75 8E E5 C9 97 44 D5 97 7A 98 8A F3 83 F1
 B3 DC 9A 5D F3 8D 93 9E 5F 30 DF 20 86 DD 55 6C
 AB 8E BA 18 BF 76 98 17 7A 27 1F 0F 81 14 88 C6
 16 0C C1 FA 9C 53 8B 8E A8 A1 2F 47 0A 71 8E 2E
 2D 6A 6F 5D F7 CC 9B 50 AF FE 20 41 F6 16 5D 92
 D1 03 B7 3A 20 62 E6 09 79 24 77 ED 86 7E 1B 5D
 66 36 F0 FC A5 0E 82 A6 DA 6C DD CB 94 FF D2 C8
 12 CF C2 AC E0 ED 5D 17 5B 13 EA CA 89 6D B7 46
 B7 C3 73 8E DD E9 4C DA D5 F8 4B 5D 1F B8 7E 88
 4D 52 94 DE 79 50 0E 2A 71 84 4A F3 CB ED 08 B7
 32 3F DA 34 E3 84 FC FE EB 95 94 2E 32 67 E1 81
 36 40 6B 7E 27 E7 D3 E3 8E B3 81 9C 16 7A C0 5F
 57 7B 7C B5 F6 4D 98 60 B5 B0 5E E8 48 D2 49 C4
 CE E1 40 5F CA 4A 05 C9 C3 7C BC 79 15 62 D1 F4
 5F 95 9D EA A5 9E 07 A4 81 66 25 B4 FF 41 8E D2
 63 84 5E 4C C0 93 3A 31 EA B2 60 CB 48 EF 4C 1C
 6C 46 F5 CC 55 26 AE 53 98 86 A3 FF 2D 45 70 86
 35 E3 C8 7D AB B5 DF F6 96 7D 17 11 5C F8 EF CB
 6B FC DB 99 65 D2 F6 58 78 E5 77 58 D9 89 AA 2C
 65 B2 01 FE 45 17 51 DA 7B 30 FB 82 77 D3 36 0E
 C8 49 DD 33 2C 5D F3 84 9F 25 A9 78 DB 5F 37 DC
 B3 D3 2B A2 F5 09 D6 72 58 A2 53 FA 95 5D D7 9F
 0E DC 4A 98 F5 B0 92 67 CD 3C 82 25 EC C9 4E 9E
 C2 6E 53 CC 00 02 FE 94 F8 43 10 FD 2A 6B 2C 93
 C7 83 BD 31 2D 66 5C DB D3 41 35 04 7E 5E B6 8D
 7F 56 2B F1 D6 B0 BF 7D 71 84 DB DA 24 53 DD D8
 72 DD 74 6F E0 96 65 66 36 B7 85 53 B4 72 94 19
 B7 67 47 8A 5F 63 D3 96 59 5C C3 EC 9B 68 F5 F3
 4F DA 52 47 A3 A6 BF C4 78 ED C1 B0 FB 06 4A B2
 F1 ED 9A BF 05 80 49 2D 0F 49 DC 72 72 1B D2 11
 80 A0 70 B6 08 DF 78 CD 06 3C 20 67 33 AC 76 96
 13 B7 62 DB 0D 1F 23 89 FD 41 0A 1E 46 47 79 21
 DA AC 60 61 D1 35 C8 90 49 53 4F 73 78 60 9C 45
 E6 4C 13 58 19 8F D9 E3 B3 D9 11 87 A9 BA 06 AA
 BA 73 F2 76 C0 00 FF 7F AD AC 6B DF CE 36 4B B4
 4D 62 54 8E 59 BC 63 19 70 45 D0 74 3E 5D 9E 04
 23 AB D9 F8 55 B6 55 57 8A 78 0C CE 7F C9 51 FD
 B8 34 AC F1 4D 19 C0 DA A7 24 DA 75 A9 EE D3 E1
 CB 13 AA 38 C9 FF 02 E9 38 69 99 A1 27 B9 12 EE
 C9 0D 6F EE 41 96 C0 FD 73 7B E3 F1 0B 18 CD 2F
 6C C3 35 CC 5A 72 B1 B7 C5 F8 53 4F 49 E3 AF 75
 47 F8 4E 55 CD 28 05 50 F9 80 5C 42 9F 63 76 99
 3D CA D8 E8 A3 8E 78 D7 D1 10 58 4D 2C 38 81 4F
 22 00 E1 84 2D B8 47 BB 3A B5 65 FF 27 94 40 CC
 38 63 24 42 69 E1 AD 0C 76 A6 9A 41 BD B5 CD C5
 06 FE 09 08 99 E1 C7 28 04 73 DA 66 74 8E 72 44
 9A DC AC 30 A6 A5 14 93 C9 AB D1 7F CD DB 4D BB
 20 34 3F 5A 9E 38 EF E7 BF E2 AB 7A 69 CA E8 9C
 DD C6 CE 20 D9 11 D3 65 C5 0C E9 23 E2 26 F3 6B
 3E FD FB 5E 80 71 FA 59 49 79 4A 65 6B B6 3A E3
 66 1F AC 28 5A 57 C4 32 54 6A A3 A9 26 A5 79 E6
 24 D6 40 32 77 61 C2 56 E4 C4 CE 5C 06 04 FF 10
 FF D3 38 43 BA F2 6B 23 F5 1D 81 34 94 83 8E EF
 FF 3B 48 8C E2 1B 7A 0E FB 36 F2 78 61 12 10 53
 D6 92 95 AE 24 C7 17 85 81 19 26 13 54 FB AD 3C
 C3 83 7E 04 67 C9 DE 82 7D 8A 67 22 79 E7 C1 E7
 67 B0 AA 05 10 51 BF D2 56 53 5F 5A 30 54 D7 9E
 1B 62 DA 76 6A 1C 82 9B 75 20 FA 5E 71 D2 49 D7
 CF C5 F6 50 B6 F0 29 AA DB 38 E4 D9 6C CB 58 14
 18 DE 68 45 E6 94 8F F1 17 FD D3 49 83 B6 96 84
 F3 6D F9 BF 4F B7 C8 9F CB 07 9B F6 D3 AD 18 11
 8E 9D 65 F3 28 63 F0 01 96 5E 9B E2 6B 64 FD 50
 7B B8 1F F9 03 38 52 0E 59 B7 F4 08 3F 57 C7 E4
 91 34 B3 2E 75 2D 36 AC C7 EB 59 BE 14 F3 CC 13
 D0 08 F0 F2 65 6F D6 8E B6 30 0F 33 8E 27 2F D8
 89 A4 AD 1D 24 BF 37 CD 1D 17 59 51 8B 47 AA 45
 56 3E 86 46 CE D4 9D 98 9F 5E E7 A1 0A 47 48 13
 B4 DA 27 44 C4 C8 38 35 98 10 34 3E B0 52 D9 7F
 83 E8 BC E5 CB 9A 1D 61 FD 35 4C A2 AA 0C 1E 7C
 22 75 E8 6A C4 14 CC 3D 58 40 34 76 D0 3D 3A DC
 BF C6 AD 00 12 A5 F5 74 75 BC D2 93 FB 5C D3 F4
 5F E1 E4 62 80 9F 22 E8 1D 29 B6 8B D0 A2 1D 06
 F1 AB EA D4 BF A1 F8 7A 2C E4 1A A2 3B B6 FC B4
 67 7B 47 FF 84 03 2D CA 4C 79 7E 08 9C 55 D3 5E
 AA 1D 28 3C 17 7A AE A6 43 39 D6 15 01 31 E3 18
 17 A0 64 B9 0B 01 A9 5A 36 A8 5C 6F 87 1E 36 9E
 99 4F ED 09 89 E5 75 07 CE 41 64 2C 6F 8A 0C D4
 4D 0F 44 46 8E 73 16 19 F1 D3 3F D2 2A A5 62 8D
 7F 68 43 07 C9 54 24 0A 93 BF 69 C8 64 3A 8C 55
 6A A4 EF CB 52 EE 03 0D 26 E1 40 36 26 E9 28 E7
 8D 74 B0 8D 09 AC 7D 03 A2 E2 1D C1 23 CF 3E 50
 E6 66 BC 64 24 FE 50 D6 D7 F8 48 04 56 F6 9C C4
 70 6E 95 AD 84 BD 19 BF 4D 40 CF 72 C0 0B BF B7
 50 FA 89 4F D1 C4 AC F5 C0 FC DD 26 C3 9B BA B3
 F8 59 DD AC 69 E0 CA B3 0A 71 B5 2F 44 B7 17 A5
 7D FB 9E EB 84 6B 09 84 D1 37 95 85 1E B1 E6 52
 92 6C F8 04 E5 C8 D5 9B 08 D2 C7 36 A4 48 4E FD
 8B DC ED A5 5C 0D 56 E8 D4 1C 00 CF C7 2F DD E7
 32 E1 3F F4 55 F7 4F 3E 0B 67 6B E2 DB FC 68 B4
 0A 6B AB 7E B1 E8 8A 1C 5E 2B F3 DB 29 13 21 14
 88 4F BE 4A 76 22 47 9A 2F FA B0 DC 1F 61 E5 8D
 7A 60 FC 5B C3 7F 93 23 EF 30 90 6F BF 6F CA CD
 32 73 61 A7 12 E4 38 BD 5F 6C 6C 5F 0E DB 1D 34
 FE FC 2D C3 20 C6 85 47 02 1B B7 F8 E5 F4 85 F3
 1B D9 0E E1 28 B7 61 92 B5 85 95 3C ED 14 22 9C
 78 E2 7B 6A 89 CB 18 98 B5 94 27 D2 36 5C 25 8D
 45 52 11 DC E1 39 91 B3 4A 8E 05 79 84 12 07 67
 27 C2 EB E3 03 91 E5 F0 45 01 9E 56 80 A7 C0 5F
 4B 1B C4 06 33 66 55 A6 1D 77 1E 59 3D 3B BE 06
 A7 7E 19 81 CD 21 C2 8B CC 14 78 8F 6A 23 9A 56
 BC EC 26 28 D4 83 A3 63 16 01 2B F5 E7 BD FB E1
 C4 D4 94 A2 EE 73 39 EE C0 2B 29 FD EC BD BF B2
 4A 5F 00 97 09 E3 47 2B D1 58 AE A1 E7 41 DC CF
 51 20 6C 33 A4 00 A6 BB C7 36 42 B8 09 E6 55 18
 AB 95 E3 50 1A AA F4 2F 7E 4D 48 16 8F 14 34 ED
 2A 43 C2 AA 01 C7 AC CA C9 4E FA 05 88 B4 1B 40
 FE 71 AB FC 72 81 03 DB F6 9A 19 3B 0D AD 45 6C
 C6 3F 8A 52 DC CD 5D 6F 6A 26 36 15 9C 1D D4 56
 5E 24 81 BB CE A2 25 BC BD 3F 18 FE A1 4E AF B2
 10 EC D5 FC C2 F8 FA E9 9C 7E B6 04 AA 6F 63 64
 28 66 90 EE F9 08 83 1E EB 2F 23 50 6C 07 43 79
 2C 06 57 33 EC 81 7D F8 5C E3 EB A1 8B 0B 2E 4E
 30 B6 BD BB 41 AB 71 AB D8 F2 2C 71 24 6E 60 77
 4C 43 82 05 20 66 FD 50 C7 E4 97 E4 66 D8 C5 E9
 5C 5D 4F 33 D2 C1 43 45 29 13 11 D8 7B C6 7C 8E
 CE 9D 17 88 66 D0 A8 D2 7E 99 F7 87 C8 9B A9 BF
 BA 40 D9 17 58 61 F7 92 0F 4A 99 4D 1F 1F DA 51
 34 7D B2 B9 69 90 25 37 9C 91 A5 C4 D9 DC EC 59
 9A 9A 9A 1C 23 10 70 4B 98 D5 48 6A 9A 75 A0 76
 2B 19 FF 43 9C A3 7E 14 2B D2 4F 12 FD 49 20 E2
 6E 19 17 B4 AA 24 7F F3 55 AF 04 47 3E 09 37 4F
 32 E0 F2 D0 BE 09 FE B7 BB 70 4D 3B 13 76 D3 8A
 8A 2C 52 01 A8 ED C4 83 CA 7B B3 34 B9 CB 3B A2
 6E 46 63 9D 54 A2 3B E0 28 4E 72 1F 63 ED A2 3B
 6D CD 8C D3 B4 62 D0 5A 5B 01 0C D2 09 54 70 67
 E2 FB 9C C0 F1 62 F9 3B 80 AC 2E 1F 88 54 B4 FE
 7D 10 19 DC 87 7C C8 08 A7 F4 E8 27 85 52 87 76
 3F 3A 1B 10 6B 3F 22 E8 2F 3C F2 F5 43 F5 03 FE
 EC CF 7A EF 80 A6 F8 D9 CD 5B E9 FE 8F 39 0D EB
 97 0D 13 97 02 94 75 A1 22 AB 29 10 DA C5 BC CF
 7C CE 3A D6 22 52 58 83 13 6A 53 06 13 AB 25 E4
 47 0B 56 A2 53 4B E5 F4 69 D6 5E 15 0E 57 43 8E
 38 91 D8 E3 B3 1B 84 3F F7 DF 59 E4 45 2F 90 C6
 6F 4B F3 10 F9 AD 35 B7 58 06 24 69 32 20 68 46
 15 8C E1 A4 A9 E8 AB 08 5B 7F 0A C2 B0 D6 78 8F
 75 BD 48 BC 43 EE 49 9E 02 57 43 A4 B4 E6 30 A8
 C2 88 7E 58 EE 1D 2C 5D D6 F2 78 BE 5D D0 C1 C0
 51 7B E3 6B 43 F9 A5 35 65 A8 99 70 B1 24 BD 70
 EB CE 2F 78 36 B2 96 2F DC 2F 70 D5 62 8C E6 B5
 9C 17 7F 05 1C 75 D3 36 11 0A C1 9C D9 FC 36 29
 FE 77 E0 26 08 48 6F C9 25 95 16 98 3D 20 72 DC
 D1 72 9B CC 04 4F BD 5A 74 D7 5F C4 D2 74 A8 EC
 41 B1 C8 6C 25 31 89 AC 58 0E 54 7D 5A 4E C1 A1
 38 3F 5C DE 3A 42 32 E0 BA 31 A3 E8 1E 40 6A 41
 D5 E4 44 B0 0B DA C7 ED 12 BC 82 15 4D 46 29 92
 CE 36 AE 56 D3 C8 16 32 A2 8D 6C DA DC C6 FB 76
 11 99 96 ED 17 B8 96 16 F9 67 CB C9 32 B6 66 C6
 7F 64 71 8C F5 04 4C 8E 03 3E 54 FA 75 F0 27 E1
 99 FA 97 FD A6 A9 5B F6 D0 BD 73 53 97 C6 5B 8C
 A3 CA C3 A2 FB A3 B6 A0 E5 15 53 DE 2F E7 6D E9
 78 D3 32 85 5C 2A 82 69 3B F6 E4 72 06 AF F5 9E
 71 32 17 3A 0C 63 18 07 FD C0 7D 44 01 02 92 13
 6F 94 E1 FD 30 7B E0 D4 88 21 67 7B CC 0A A5 8B
 5A 61 12 CF BA 32 5C 76 96 8B 7C C2 15 F7 68 B0
 BF 28 66 F3 DC FA 05 3B FC 24 91 C8 20 48 D8 A7
 A1 CD 9E 6A CC D9 5E CF A1 AE 5B 1F AE CD 2E 96
 B5 96 87 15 62 25 7A 6A 0E 65 28 CD CC 65 B5 31
 C7 F7 A1 6F 03 18 90 BC CE 10 15 37 53 76 D2 DC
 A3 51 68 DB D0 6F E7 52 A3 8E A6 51 F5 4B 96 CA
 DD A9 60 A6 6E 3B BB 0E 96 F2 52 78 93 18 8F 03
 C1 15 B2 96 15 42 19 FB 9B 26 E8 5A 11 DA 67 E0
 C8 42 47 00 22 8B 3C A8 5F EE 68 0C CD 8F C3 65
 7F 07 CE 21 9C CA 3A B8 F7 42 11 CA 5A 39 6D 72
 77 3C 37 8B 97 C4 A5 0B D9 5C 88 B8 FF 71 B7 8A
 84 9B C3 3E A9 24 31 C5 90 2B 35 48 1B A9 1D 14
 38 EE E7 88 F9 CE 46 39 61 D2 57 59 A5 E9 3E CD
 61 ED 8E F1 50 E7 A3 0E 0A F4 12 A6 4A 96 0D 3E
 9E 57 DC F0 DD AC BF 32 E9 ED BB F8 FF 4E E2 82
 2B 35 FB 36 7F 54 5E BB 96 4E 24 60 88 B7 6F DC
 24 57 E1 AF 15 0C 65 33 F0 18 1F 9C AC D6 84 AA
 44 F8 DC DC 82 1C 0C 13 7A 9F E5 BB 21 58 BD 3D
 E4 C0 4D 97 03 77 FA 32 E5 38 D3 54 08 CA 44 7A
 D0 6E 9E 6D F1 0C BC 8D 33 56 BF 53 21 67 30 1A
 8D 3A 18 EF CE 79 FF 1E BE 45 2E F4 8A D4 9D 0B
 73 AB 5A C3 F1 65 CD 9B BB A1 C5 FF DF 49 E0 CB
 CE ED 4C AA 3D 49 15 51 5C 44 3C DE 46 36 C4 6C
 80 42 FD E7 F8 7B 56 84 A0 F4 6B 46 06 29 94 79
 0A 9B D7 80 C1 B0 4C 4D 69 44 36 FF 70 4C 4A 84
 8E 30 6D 3C 33 02 87 68 8A 86 C5 2B A3 BE 2D 2F
 29 8B EA 39 2E 03 D3 68 32 D7 8A 35 BD C8 79 FE
 7B 4F 4C 67 92 F3 62 67 14 F0 16 70 90 22 C4 DC
 36 84 4B 27 9C C6 6D 0C 33 D2 B5 8E 58 BC 4C 5E
 A0 A9 C6 01 E6 3A 37 D2 A0 26 5F BD 95 CD D8 53
 3A 72 1B 7F 46 54 21 C3 AF 7A 67 CF 8B D7 A7 3E
 9D 57 EB 63 E2 3D B4 8C EE 34 D7 4E D7 34 A4 04
 17 1A F0 D2 9E F5 00 05 9D 6B 6C B1 FC B6 65 4E
 2E 53 05 32 5E A8 EC 63 CF B6 BE 4D FA 4F 1B 6C
 11 AA A7 5E FB EA AE 0F EF CA 30 7D 4D C7 5A A2
 93 C8 60 65 4E 6E AB B3 53 B2 DB 26 13 76 84 07
 8B 69 DC B1 9E 73 95 19 B6 11 C2 3A 52 A9 86 87
 3A EB 49 DB 24 93 41 40 09 10 B7 4C 90 CB 7C 19
 24 02 49 32 1C 10 26 2C 64 8E B0 F9 48 16 9C 59
 D5 DE 22 85 5D FB D6 0B 9A F7 04 60 C8 7E F7 86
 B9 27 39 9F 24 5D E1 5C 70 E1 B6 C4 28 E5 61 14
 29 D3 E6 DB 8E A8 FB AC 33 25 C0 65 CA 7D 61 20
 B5 C0 AE 02 69 41 24 91 05 FC 9D DC C3 CF D4 9F
 52 29 99 7D 5B B3 78 80 5F 5E 41 FB 8A DA 16 24
 C0 32 1B 20 30 1F 07 1F 12 40 EC D6 8C EE 09 AB
 BF 3A 52 BF F0 10 5E 4B 5A B1 FA 41 8E 8D 73 20
 63 99 67 0B E0 99 B2 92 9B DE CF 24 FB 50 71 60
 E9 9F 8A 87 1E 7C C4 5E 38 38 19 14 39 1E CF 60
 C6 09 82 E1 16 8B AE 3F 87 89 18 59 69 1E 91 DC
 62 7A 20 66 7F 41 15 18 06 A6 73 03 8C 61 9D F7
 59 89 D3 02 39 EC BF 31 75 9C 38 28 6A C8 6F 0D
 14 29 BB 16 98 E4 12 34 BE 38 D2 D1 AD D9 9C 26
 A4 80 61 95 78 49 48 09 B5 EC 48 C8 8B D7 7C A8
 5F 28 F0 7B 23 A2 2F 53 3B EB FD 93 B1 AD 01 15
 8D A4 6A F9 37 B9 9F B4 CD 71 3F 3F AC 54 51 DB
 DF AC DF 3F 01 01 96 36 A5 38 BC 3D C4 4C BE 4B
 57 4D 8D F9 B3 3F BB 82 6C B6 5F DB E7 E3 67 5C
 1F 2A 1C 7F 74 CB EB B8 A3 90 FC A9 0D 49 12 41
 C6 63 77 9D 99 60 77 86 8A CF A9 C4 B1 F2 05 C7
 2D EA 2E F2 19 38 C7 E0 2C 51 E6 C7 C1 5B 0E 72
 2C 64 AB EB BA 68 CF 03 51 F6 64 18 29 37 A7 D0
 8E 8B FC 43 76 12 3F 0B E1 2E A7 0A CE 79 FB F2
 AB F2 DD 0B 1F 09 58 B5 97 22 E8 C6 CE 01 D8 2A
 93 DF F7 C6 E2 A1 65 B7 6C 58 C0 AC 99 8E 6A 70
 A6 71 26 89 E9 27 FB 47 71 56 30 6E 89 94 B6 97
 7B 48 28 C8 34 5F 52 A7 6C 63 94 87 34 17 CF 95
 C3 46 22 7B 73 78 B1 6A 6B 55 37 86 BC 16 6F C3
 02 D4 54 F8 A7 F7 62 47 82 5B AE AA 46 FA 28 C2
 F6 20 E4 8B 8E B4 ED D5 68 AC 0B AE AC 27 1D 1B
 5B 75 5C 6F 1C FE 0B B4 34 DB AA 79 62 3F 83 D4
 C8 ED 97 6B 5D 1A C3 2D F7 DB 3D 24 DB 18 B2 D5
 C6 BB 0C AC EE 02 B3 B6 46 D7 AC AA 81 CC 4F CB
 8E E3 43 A1 8B 59 9C 65 D6 F9 E5 65 D1 C0 21 E9
 94 3E 0D 66 36 EC 79 E5 6C F5 07 DC 28 07 F4 04
 6B 1B 94 D8 04 F9 77 73 94 5F CC D3 0F FA BB 71
 EB 2B 66 BB C2 28 0C CF C5 63 1B 07 81 C1 71 82
 0C 28 A8 55 08 1A 91 0A 27 C7 8A E9 D8 26 1A F9
 29 D4 98 DB 17 D5 E6 EB B1 52 78 14 25 41 5C A8
 2F 0B 42 C1 C7 FB 00 5B B7 96 A7 8E 76 98 D0 9A
 34 3B 52 25 B6 FF 4A DF 1C 1E 17 29 99 40 A9 BA
 5F 16 12 48 8D CA 7E E9 BF FE 2C 6F 4D 9A 48 F6
 CA 1A C0 4A A0 16 59 8D A2 3A E0 17 03 32 05 13
 92 98 CB 20 DF FA 65 53 83 15 21 D6 01 AD 57 A8
 BC 2D 7A C4 4E 59 BB F2 99 D6 25 38 BB 26 3E A6
 22 AB B6 CF 23 0D 39 A4 49 6D 28 50 C0 63 C7 77
 51 F8 E7 BD 56 D2 B5 51 15 BB D8 D6 18 0C 89 AC
 44 12 F5 D8 D9 D1 98 6C 54 4C 60 F7 D3 38 15 8B
 34 54 31 C8 43 25 5D 48 1B EA 9D CA 79 B0 DF 28
 58 A8 34 10 4F B6 E4 46 0D 4C C9 66 27 A8 44 F3
 01 C7 35 E1 3A 79 22 61 A5 E6 35 DE 27 D2 8C A5
 F0 4B 16 7E F4 54 E3 8C D9 68 1C 3C 2C 76 C3 84
 C6 EC B9 35 45 85 61 0F 52 73 97 83 C8 2A 68 88
 B9 50 73 88 87 40 3C 1D 86 40 76 41 DD CC 13 81
 AD DE 1F 44 A1 19 4B FF 6E B6 3C 93 61 DF FF A8
 D9 C1 11 5A 08 BC 7A B8 23 06 1A 10 EA 5B F1 EF
 99 DF FB DA 35 1B 22 1B B1 35 FD 99 11 3D 7B 0B
 D0 0D 59 2E 67 CC 47 40 23 E9 A6 D0 57 16 22 59
 9B A9 40 A6 05 CD 8E D7 5A 29 3E 2B 04 A9 4D 2C
 2C 06 62 FB 93 58 FE 92 10 0B 19 62 E9 76 C4 E4
 37 22 30 E6 A2 E9 97 D9 DC 05 D6 96 18 B0 BB 2A
 3F DF 60 A1 55 AC 1F 6C FA 45 D6 A6 3A 73 44 B8
 EC F3 52 93 2B 2D 37 23 15 40 C0 0A 95 A4 70 F5
 B7 CA 63 A0 E5 87 1A 99 16 CD 3E 24 70 13 0A 10
 A0 E2 84 91 7F 2D 34 B1 DA FE 78 3E 39 12 A4 40
 A5 0E 39 86 0B D3 D9 AE 0D 6C 98 DF 12 CE 6A 5F
 DE 85 D6 04 05 DB 01 79 83 E0 18 72 75 27 C8 42
 A8 3D 68 21 81 BD 81 61 07 FF 1C 08 47 0B 18 A7
 A5 AC CF 8F 39 F5 14 38 F6 4F 63 01 0B 59 C9 27
 85 BC 4D 52 1F 61 1D 2F F7 8F B1 8F 76 B1 D6 80
 E0 38 8D 71 34 F9 04 E4 B8 90 04 CC CD D4 F1 66
 9C FD 8F BA C0 90 21 E9 37 E1 6D 25 46 48 98 FB
 BA 44 65 FA D6 CE C0 23 62 9C 68 54 1E 2D 38 AA
 42 5A 67 8A AF E5 A7 DA 19 60 04 14 75 3F 96 8F
 83 4C 14 3F 84 84 6E 73 A4 C8 8D F7 29 FE A5 F2
 A5 96 AC 3B 88 4E 98 0F 93 56 CD B1 C3 F3 89 60
 66 0A 67 3C 4B AC 5D 3F 01 E0 0E AF EB 56 B1 0F
 A4 E0 2E 04 59 79 7D E1 EC 75 9B 7E 72 3A C3 6E
 3A 11 66 81 A4 4D 75 0C 80 01 A9 29 BD DD 88 E4
 0A DD 16 57 1E C8 22 22 D1 AC 51 25 99 84 94 9A
 F3 41 57 52 99 C1 F4 FB F4 28 E9 56 89 EE B6 2C
 19 99 64 0C C9 5C DD 48 01 B1 0B 56 A4 54 90 0B
 F6 4D E8 97 88 AA 82 00 44 2B 09 2C 43 C2 52 BF
 06 89 21 6E 2F 73 7C 61 8A 30 36 14 56 01 EA 10
 1F 29 C1 2B 11 3A E3 53 FC D2 9F FF E2 AE 4D DB
 EA 0B 86 1A E6 09 4C B6 2D 41 A2 7A E1 8C 8A FE
 07 3F 8E A8 87 99 63 1E C2 B9 9A 2D 68 83 64 40
 B5 0C E9 A9 69 26 C3 17 3D D1 05 C2 67 87 AF 6F
 FF 49 25 D1 59 39 93 D0 AC 62 57 DB 42 00 88 13
 00 E5 F4 9A 1C 20 47 5B E4 22 E7 65 A1 B3 83 BA
 0C 72 D0 37 C6 99 8F E4 4D ED FE 2F 86 B6 6B 37
 A2 54 5F C1 7C 3A 0B 32 B3 4B 9C CA 4F 49 77 41
 0F 19 26 1E 11 00 21 A0 2C 86 50 61 71 EA 80 71
 23 D4 D0 99 6B 72 3F 56 C9 3A 6D 91 4A C8 1F 4E
 38 4F F9 01 D7 90 89 4B 89 23 8D 49 D2 3A 07 ED
 60 6F 74 CA 75 49 AC DD 97 F8 38 71 68 D6 10 8C
 16 06 B5 97 6C 4E 27 26 D3 CA CC 39 13 46 0C BF
 C6 44 A0 DE 13 58 39 C0 90 43 17 C7 E4 1F 89 02
 61 5C 5E 40 33 EF 27 B8 1C 0D 14 2C CD 8C 95 4E
 C7 A9 A0 FB D2 12 1B 66 12 EE E5 A7 21 AA BF 62
 72 7E 24 43 BB 37 EA A9 E3 5E CE 61 F8 0D 1F 9C
 88 F6 C6 B7 B6 DC 3F F8 73 A9 86 AC 6E 7F 32 0A
 B6 74 27 C7 8D 1A 86 51 6A 39 3B D9 86 82 DC B3
 94 9F 3C 9B 4C F0 5A 0E C0 15 A3 27 9D 78 2A 22
 EA 0B 9D F3 29 8A 12 17 9F 08 C3 64 6C B1 49 FC
 DA 29 98 36 EF 54 6B 54 5D 10 15 24 EF 1C ED 1B
 A4 01 61 7B 93 A0 87 11 26 55 77 1C 2F DF BC 33
 54 09 38 C8 2C CF BD 78 A7 57 77 AF 8D D6 84 A9
 9A 39 45 60 24 28 46 2C 61 A9 FB 85 D7 51 BC F2
 E0 CA 24 3D 91 03 D1 FB 08 8E 53 9C 97 4D B8 1C
 0E 37 B9 47 A3 26 53 C6 1F 3C 90 0E E0 95 0A DA
 D1 A8 92 85 AE 1B 04 11 6C 53 1A BA 36 8C EA 19
 78 79 02 45 29 06 F4 CC 8E B0 62 6F 0B 60 45 9A
 61 CE A6 91 42 BF 17 4A 86 03 CC 18 47 81 45 B5
 08 E6 0D 16 F5 C0 61 26 8E AD A1 32 5F 87 31 59
 C2 BB 85 9B 49 46 40 0B 3D 2D BC F9 66 D6 D1 94
 52 3B 63 92 FA 12 ED 7E 1D C7 CB 24 F8 7D 77 F3
 A1 92 12 C1 D2 7F CF 0D 90 75 90 EA 06 4A F9 3F
 27 D0 A1 C1 46 81 25 45 4D A9 48 7B 89 90 08 21
 6D F6 6E 5B F9 A6 91 A7 72 F7 0E C0 1E 83 04 5E
 DE 4E 4B F3 FB 75 A1 8A 92 A8 42 E3 D9 AD 2B 9D
 CB 82 2D 20 3C E5 C6 ED FD 56 00 9B A6 6F 90 72
 C8 16 8B F0 42 85 88 9E C6 E3 B1 28 6B 67 53 D4
 54 3C 2B 54 42 33 55 6E 45 6B E7 0A 91 7F 16 B1
 C8 FF 36 12 5A 7E F9 AD 68 53 9E 52 3E 28 61 9B
 43 3B DE 69 6E BC 23 0F 18 59 F9 40 C4 34 90 0A
 D2 9F 14 39 E0 E9 2D DF 42 42 72 73 62 77 E5 4D
 BE 05 CB FD DA B2 89 DB 00 24 8C 99 3C E5 D8 71
 A8 3B 64 13 02 F8 61 45 53 5B 49 6F A9 36 25 DA
 B6 DF 26 CC 44 52 99 BC 28 F5 D1 C0 D1 0E 90 42
 85 E3 C8 B1 9F 2F C1 1C 02 59 B3 16 24 B6 11 73
 8D 38 52 98 4D A7 E2 EA 5D 4D 12 B3 CA 5A CC E4
 33 33 45 4D 21 DB 0E D2 27 76 9A 7C F3 F9 8F C1
 C5 03 4E EF 6F 54 2E EE 1F F0 DA 6F 85 BC 62 7A
 08 9B 22 15 FF 5A AE 53 27 04 1C D8 C8 B7 65 E5
 00 9A 6A 7D AD 0E 4E F5 70 CF 35 E7 A9 6F 73 CD
 B7 6D CC AB A5 23 28 8E EE 2B 7A 4E 6C B0 BD E7
 70 D0 34 DC 24 4D 15 7F 66 BB 33 60 FF 19 EA C3
 CB C2 97 2D BF 1F B1 28 1D 22 9E D3 66 1C F5 64
 A0 CF 99 9B 4E F2 6C 8B E2 DB DF A3 83 9A AD 54
 5B 20 BE DB 0F 9D E5 B9 B8 AA 11 46 C6 87 DD 3C
 BB E1 36 C1 58 1F 6A 46 DE 30 F3 6E F6 90 00 EA
 2F 71 FD D2 03 2A 4B 28 9B 9D 77 18 8A CD 9E 3A
 19 E1 5D 0D FA 30 01 0D 83 90 52 BB 2B 86 72 AE
 B8 35 B0 B7 B9 D8 C5 43 56 05 9C 14 AD 4D 84 0A
 F3 5B AB 94 9C 74 C1 F4 98 1A F8 C2 B7 2E 75 71
 70 45 EF EE 02 62 71 3F B4 64 55 62 01 4A 61 AF
 9C 37 8D DA BD 4D 52 2D 3A 32 3B 38 9E 49 5F 14
 1F 80 2C 29 AB 15 C8 14 50 A6 B2 1E D6 A7 16 F9
 60 82 3C 07 9E E9 DB 5B 30 AD 32 0D 8D 47 23 AC
 6A 19 02 7B C8 07 66 4B C9 19 BB 32 F2 C4 FE E8
 3B 8A 66 0A F1 07 82 8E 46 94 90 56 67 EE 06 FE
 D9 9B 78 0C 25 43 C9 00 F1 0E 9C 1D F2 EB BA 94
 A1 F3 35 B6 6B 85 D8 3C 5C 3B F0 53 A4 1B 0B 42
 14 23 62 89 DE 68 3C 22 6C BA F6 B2 59 1E F1 0C
 AA C9 67 D3 33 35 CD CB A4 5A 65 C1 AD F3 0A 3F
 48 3E 94 FC D7 9B B6 29 5B 03 67 73 DD F7 56 0E
 3C A9 51 D0 F1 77 26 0F 07 D8 EA FA A2 1C B2 47
 76 06 DC 2A A9 1E E4 A6 FC 73 51 E7 6B 93 4C F9
 F7 C6 9D FE 00 7F 9E 94 63 33 11 EC A1 43 28 B0
 FC 6F 21 73 15 FA C5 27 FE 0E 75 31 C2 4D E9 64
 5C 47 1A CD B0 58 A5 3C 02 78 1B AC 1C AC 79 3F
 03 FE 18 7B E7 15 8F 05 0A A1 AE 92 31 BC 0C C0
 04 26 6C 10 F6 0E F0 98 96 5C 7F A2 8F BC 75 26
 5F F4 0E F5 5A D1 24 4D 8E 82 3D 3B D8 AB 23 EF
 91 C8 57 BF 10 30 C3 F6 0A 54 7C 4E 27 4D 0E D1
 88 E6 A2 CD 24 95 BB 73 0B 43 47 05 F7 F7 BD DF
 D9 DA 81 40 37 36 89 10 8F D0 13 99 FA D7 1F 1B
 07 34 5A 3D 82 2C 15 75 18 62 30 E0 FF ED DC BD
 FB D3 6E F1 3D E0 03 D4 99 3D 09 34 10 2B 16 67
 F9 DA FD C2 94 A8 F8 51 80 0B 86 F6 C7 AA 8B C4
 9F 17 FF CD 41 F7 F7 7D 25 97 A8 F3 30 E9 CB 20
 23 8E D4 49 E6 79 2B 07 4F CF AF 8D AD C2 48 D9
 B8 D4 D7 49 27 BC F1 F4 52 E2 5B 25 FF 40 A2 AB
 12 BE 0C 96 01 9A 77 34 39 51 A4 26 58 E7 CA 9D
 FD 57 CE 4F 66 22 3A 98 C5 52 AC 04 81 ED 7A 0B
 CD F7 28 89 50 05 A6 DB 7A 28 DC C5 7F D3 E8 93
 73 85 0F F0 91 E1 C7 21 A4 D8 C0 13 88 4C 1A E8
 D8 2B 4F DA 1F 3B 20 42 D7 13 DC 28 1B 26 CD BF
 CA B5 D1 A3 B6 F8 39 E9 4D F7 2A C3 54 95 16 4E
 CE DE C4 70 BF 32 BC 79 85 07 B1 47 34 8D 6C C7
 BB 47 40 38 00 21 51 7F 9A 95 4E 14 CE D2 41 82
 26 B5 B2 B8 DD 35 6C 68 6C 3E 22 F3 A9 11 3F 14
 EF 36 85 1D 7C 8C E2 94 0D 38 DB 13 74 C2 C3 AA
 02 E6 14 A2 DC EE F6 00 5A 61 E5 B6 A1 5A 8A 5E
 F7 BA 8B 0A 6E D5 08 8F 46 2E F7 58 76 CF 19 3C
 75 4D 50 63 E8 3D CE EC A1 CC 71 12 31 F4 13 90
 33 7B CB 38 6D 95 70 38 E1 02 70 2B 6D 56 82 77
 AB 89 58 15 83 2D C5 B2 96 F1 1F 54 8B 0F AF 37
 32 E4 98 3B C7 04 3A 1B 70 01 6D 6F 7F 45 68 E7
 80 E8 A0 1D 1B 1D 15 19 1E 9D 58 BE 67 CA 4C BE
 6C A8 B4 12 68 A7 3B 83 99 26 D7 FA D6 8F 96 E1
 8A 33 46 43 05 C7 CA 24 9F B2 A4 0F EC DB 50 B2
 19 BC 07 C9 A1 2B 6C 58 7B D5 3F 2E FD B7 A6 9D
 2D AC 24 13 6A 29 28 DA 3C 78 50 CC FD 2C 4B 96
 89 83 DA B3 1B D0 95 CE F8 DC E7 B0 CC A9 11 CD
 95 B7 C0 52 D1 2A 02 DF A7 9A EE C1 58 B6 6C CE
 C2 55 DD C0 5B 10 B9 7C 1B 35 8C D5 99 CD EC 45
 EE FF AB 75 8A E2 B9 8E 96 31 66 5D 7E 2F DD F4
 2F E2 CE EB 7E ED F5 AF 81 1F B0 D4 E7 C3 0A E9
 67 0A E7 3A 6D A8 D6 8D 79 D7 23 26 6F 45 69 36
 D0 B3 DF 00 29 CE BD 18 71 60 79 A5 24 5C 4C 54
 4A D0 74 FF 22 2D 9F 4A 73 69 FB 42 1F F3 77 03
 EC AE E3 D7 F0 85 15 21 AE 81 5D A3 0D F9 DD EC
 F2 8B 79 05 AD A1 78 84 43 6A 22 1A 89 D4 3A DD
 9C D5 13 F3 C2 9E E1 60 DB 82 58 DC D8 96 49 9B
 F4 9E FE DF 68 A7 FB C3 2C F1 A5 6B 3D C0 E0 6C
 F5 B2 96 E6 58 E6 E0 F5 49 21 EF A0 71 F9 CD 67
 24 7A 03 95 05 81 54 15 E4 8C C8 F9 16 25 B5 DC
 0F 12 F0 20 01 C6 04 2A 21 17 5E 03 8A B3 AA BE
 CF AB C7 57 E1 74 BE EC 05 DD 97 AE F3 34 9A F9
 39 E5 2E 02 A3 6C 53 E2 9B 30 38 8E 82 A2 7F 12
 AF C2 BF 98 99 0B 8C DE 1B 6D B4 12 6B BF 4E 97
 7C 25 44 38 F8 52 48 B3 EA 70 E1 04 36 AE 8B 3E
 B9 EE F4 8B F3 EC 57 56 61 AA A5 3E 7E FB 13 A3
 79 EF 72 25 94 C5 41 FD A3 F5 FD 67 4F 2F 7B 50
 77 09 EE 2E E8 7C D5 ED F4 F5 6E 61 6E 4B C1 C5
 B1 9F D5 C8 07 72 B3 DA F0 2F 69 43 E7 2C 04 39
 20 D2 FF F2 C4 02 8A 22 3C 3A 71 2A F9 6E FC 6A
 D4 AF 8B 05 36 8B FB 5B 8F 38 2C EE DB 50 47 02
 73 AF 17 4C C5 16 98 50 19 17 15 A6 82 70 8C 5C
 F3 64 66 4B 7D F5 FD 25 CA E5 4E 93 49 C5 4D 17
 DB A2 F0 3C C5 7C B6 BF 75 5B A8 1A 41 62 1F 14
 55 B5 9C 1D 93 64 8F 65 41 4C 9C 63 F1 23 B9 9F
 DC 6E BB 6B 9F A4 E5 39 D2 4A C6 85 60 5C C1 40
 0D C8 24 4D 56 7C B5 74 D4 CC 2C BA 49 0A F4 91
 27 3E 62 93 CE 11 71 CF 05 C1 3B 12 89 6D 58 40
 F5 F9 76 7D A6 CD A7 94 2D F8 9F AE 31 A5 C8 22
 2C 65 C1 5F 86 C0 E9 4E C8 D1 1B DC 17 7B 2C F2
 2B D6 13 AB E8 8E 11 2F 2E C9 B5 4C F2 4C 92 18
 53 51 EE 37 FF 27 D3 B1 7B F8 4C EF BE F3 6E 33
 19 65 1E A1 49 D9 CF 4A EF BF 2A 8D F9 8D 5B 69
 20 C3 25 69 57 C2 D3 25 8D EF 9C 3D 6D 38 75 BA
 A7 FE 62 03 D9 F3 0A D6 37 E3 BC BA 69 6F ED 03
 DA 29 3C 1A 61 7D E2 24 E3 34 07 31 03 97 6E E1
 6A EC 5F 9B 48 74 9F 07 DE 26 0D 99 9D 20 FD 68
 D7 10 AC A6 F6 7D 5B BF FB AA 6F 6E E4 91 35 45
 DA 3A B1 73 BF E5 3A 6B 85 15 2D 77 C8 A6 7C BB
 76 2C 74 5F 35 EF C4 46 6A B6 F0 AD E7 9B F9 6A
 B8 56 38 34 71 A1 B8 B8 CB DC 21 C2 E7 6D CA DB
 A7 99 21 02 C5 7E A8 8C D7 6D 0E 58 85 63 D5 ED
 55 B5 92 E2 96 A7 C2 A3 59 D0 BD 60 B2 F4 F3 0F
 C3 CA 53 7E 78 24 30 A4 A0 3C 9E B8 B7 33 D6 B6
 A4 CF 9D ED 10 01 48 4E 03 C1 6A 7C 8E 10 5E F8
 E5 21 96 AA C6 95 79 C6 69 BE 1F B1 1B 82 F7 1C
 56 24 E4 A6 0E 32 AB 53 BE C7 A1 17 3F 36 7C 78
 5B B2 21 B2 E4 8E 71 74 98 15 01 76 DD 2F FA 7F
 EF FC 34 25 86 E2 DC 5C E3 70 18 11 8F EC D0 AC
 32 E6 89 C5 06 EC 23 C7 10 76 89 4A 0C EA 9F 78
 8C 9B 5C B6 B5 69 9E 65 21 8D 7C B6 9F D6 5D 98
 33 C7 5B 90 AD 46 12 05 35 5A 18 36 64 F8 5A 7E
 92 B3 3D FF 9D 60 3B D7 4A 5A 90 7B 1B 8B 91 CE
 75 6A E5 E3 F9 A2 06 13 06 0F 3D A3 AC 17 2D 26
 4B D8 84 CD DD 72 7C 36 2F DC 38 A4 A3 98 7D 5F
 E8 E8 11 02 A7 0A D4 D1 5D 96 FC 8F 8F 9E 13 5C
 5E 76 33 1D 5B 7C 73 00 14 D3 6A 76 71 33 9B D0
 D7 39 41 06 45 80 03 B7 98 3E 51 40 5D B0 FF F6
 2D 8A E5 55 34 A8 3D 66 E0 95 93 2A 32 E7 A1 88
 D2 D8 C0 94 8C 80 55 2D A2 97 58 81 2D 6A 5F 45
 6C E9 CA 6C B4 CA 89 78 41 91 F7 30 39 84 42 F6
 8F B6 1E 24 1E 5D F1 45 D1 99 85 D8 15 69 8F 29
 93 EA 3F F8 2D 6D D9 4F 34 DF F5 44 7D 12 0F D9
 3D 8A 12 C7 94 27 61 5B 38 17 72 78 A0 97 04 65
 5F 48 96 8B 39 FB FE 11 6B 23 83 9D D4 0D 03 27
 D4 14 81 CD 3B A6 D5 C3 EF F8 E0 09 FB 4D B3 F0
 DC 43 E1 A8 14 C2 31 1D A4 C6 CC 51 D0 DE 6D 12
 CC 31 47 94 7A 66 32 B6 C5 DC 9E 47 A6 C6 B8 F8
 67 DE C0 EA F1 2E E3 94 A7 71 36 16 FF 19 CF 52
 8C A1 15 78 E4 54 EB A0 F7 66 A1 18 81 9C F9 05
 09 80 CB 98 26 6A 77 FF 87 6F A4 83 3B 74 EC F6
 A8 99 F6 A6 7A 91 E4 95 B1 73 7D 15 9A 32 56 1B
 86 D9 27 27 0A AB EC AF 8D 03 74 23 DA A4 CD 84
 0C 66 FD D9 2B 77 00 3E 1F BF E3 D3 F6 08 F7 79
 5C 01 A9 A5 FA 55 60 71 53 5D 8A 71 D1 CE BB 5A
 3C 2D 87 E4 98 DA EE EB B1 EF 23 04 FA 97 22 D5
 93 EC CD 78 C9 93 E4 0E 64 56 C9 B4 7E 06 6D AD
 1F 13 34 42 99 03 73 24 FB CD B2 ED E1 DA AB C4
 B8 91 10 38 88 5A 56 1C 7A DD 8A 61 E7 D7 0A 05
 62 98 A7 2B 0A C3 A9 C6 33 0C D9 8F 64 16 DE 8E
 ED 94 02 7A DC F0 CF 36 CD FF F8 7D 44 1F 13 6E
 88 DA 92 05 C9 8A FB DF C1 77 CC 1C F4 F8 74 3B
 32 8A 19 7C 6E AE A2 B0 57 4A 33 70 21 08 E1 9A
 82 C9 6D BB 50 5F DF 19 B7 49 E9 46 C9 26 20 29
 38 DF ED 8D 5D BC 0E 0E 10 26 B6 80 2B 79 EC 8B
 35 62 DB CE AE 34 0C 8F 71 54 5E 81 8B 7E DC 19
 FD 1A 53 F6 BB CA A1 45 BF B9 9A 24 96 60 8F 72
 27 35 E4 3E 6C 6F D8 02 B7 BC 19 1F 24 8C DF E3
 2D A7 3B 44 E8 15 91 D1 E7 2A D8 59 8A AD 43 DD
 7A 2A C1 4C C8 5E 5D 21 2F 2E 5E F0 9D 58 75 7D
 B6 8F AB 05 83 BC B4 12 6A 00 3E F1 8E A7 5F 7D
 EE C5 AB CF CC D3 DE 8C EF 47 0E 3F 99 A2 12 49
 F7 96 21 36 27 C5 B4 B7 24 DA 9B E4 92 8C 8D 50
 EA 08 31 A4 6D E2 02 68 C2 1B 40 1C 9A B0 6B 20
 BF 27 49 46 08 92 51 1E 65 48 75 1B 41 F8 7A 44
 AD 9A 85 7F 15 E3 1F 24 F3 7C 06 B5 5F AE 55 3D
 E0 52 1A 84 E7 EA 0A 00 6D 3C 1E 26 56 AF 4F 4B
 0B 0C AF 67 19 A6 B8 80 37 4B A8 37 C8 94 4C D9
 8E 8E E1 37 D6 1C E1 69 E4 82 72 FD 22 A5 F5 F2
 BE 06 2E 4F 47 B9 E7 52 90 C6 FB 99 3F 2D 67 76
 C2 60 36 69 BB 08 5A 7D B8 BF E8 CF A5 B8 CC D0
 CD AC D4 16 9B 30 A9 FC C7 43 63 2E 1B 6C D9 C4
 82 73 D6 59 86 59 0A 1F 05 2C 59 56 A6 A1 1A B0
 59 69 85 E1 54 7D 55 09 2A DF AA CE 98 D3 86 27
 90 8C 32 46 64 7B 01 00 0D 5D 72 E4 1F 66 B4 D8
 DE 2D 77 12 E2 54 CA B3 2F 3B 0C F1 FF D7 22 1B
 BA CE F6 88 AF 61 9B 54 54 C6 D7 72 41 C1 FF EB
 C7 02 98 2F 2B 2F E5 FD 4B AC 87 58 31 99 2E 25
 A9 D8 33 42 5D 62 D9 5A 48 3C 1F FD E2 81 5B 0D
 CD B9 91 95 D3 7E 98 5F 5A 76 AF AB EE F3 B8 16
 BE 08 F9 59 0D 38 DD F1 AC 10 3D 83 D4 DD 0A B2
 0B 01 C7 ED 97 4C 88 21 F0 D8 D4 3B 3B FD 95 BC
 26 69 C4 F7 CE 88 2A F9 35 0C 5D 0E 4D 50 C2 06
 37 CF 93 15 59 0B BA 6B A1 D2 D4 9B EF 8C 70 A6
 8A C0 57 B8 B7 64 44 3B 7C A4 E1 8D 7D 1D 5E 9D
 8E 2B 5B EA 7B 13 F2 00 3C 1D EC 3C 93 BA 77 B8
 75 9D 02 C1 67 AC 89 3A 18 02 4B EE 17 C5 F2 E5
 B9 4F AA 2E 56 B8 29 D6 1A 04 98 44 17 69 48 FE
 F7 7F 31 E9 42 00 5C 6F 30 54 F7 7A 1F C3 0B 31
 A7 99 BC 26 AD 66 D0 CF DB 0D AC 52 81 C5 D5 0A
 EB F5 68 D2 C4 D4 6B 0A 22 33 A1 67 2A 8F DA 2A
 E5 1A A1 EE 5E CF 03 62 80 79 2E CC 17 AB 16 16
 C2 50 F3 64 95 EF 39 24 C6 1D 78 92 DE 21 C3 F4
 BC 40 7E 92 20 62 1A 73 3C B4 55 C5 6D 67 C9 E7
 EC B9 26 08 E2 B6 6A 8B 99 2D BB FC 41 BB 9C 56
 21 AC 73 0A 2F 2E 1B E5 6C BB A9 99 85 6F 27 AB
 AD A1 C1 3A 09 52 B1 CB B4 84 8E 03 90 59 D3 B6
 41 A5 45 0E 3E 42 C4 C5 D0 95 99 76 7B 1B D8 01
 84 59 03 19 F0 B1 65 70 97 63 EF B5 BC 73 E6 EF
 F0 68 45 C4 57 20 01 91 50 54 51 DE 08 C5 48 C1
 02 74 5E AF 9D D0 10 81 65 20 48 93 44 E8 C5 F4
 9C DA E0 BF 03 57 A9 7E 30 5E 92 B2 D2 94 17 25
 47 33 D6 87 67 74 C6 60 66 BC F6 01 C3 4A 1A F5
 5F 0B 21 2C B6 B3 B9 2A 57 8B E3 53 92 2A 08 BA
 35 AB C7 9D 9A D0 50 58 B1 12 D7 7C FF 16 8E 94
 C8 13 2D 33 99 94 4B 24 E2 7C 53 18 C5 AF 57 5F
 49 2D A4 D5 21 77 7D 95 A2 A7 95 50 FB 42 10 A6
 FE 55 B8 64 CF 7C 36 60 AF 4F 2B 23 9A 2A 8D C8
 E8 98 31 BA ED F2 93 1B 22 7F 23 5F 50 42 88 45
 91 89 65 D2 71 99 22 84 26 0E 83 7F AA C1 43 8A
 24 0F E7 61 AF BD B0 05 D0 47 B4 8E EB D1 3C DD
 14 12 32 24 8E 05 F8 30 EF 7D CB 41 69 CB D8 A9
 B1 94 52 72 C1 35 B3 F6 6C 5E 40 90 EC 84 73 E6
 DC 9C 78 C1 46 1F B4 6C E4 C6 12 EF 48 5D B5 51
 63 3F 5D A7 96 E3 A0 8E D9 FE FA F8 23 FB F0 1A
 E9 5A 07 88 73 6C D9 68 53 17 95 53 CD 96 BC 0D
 AF B6 0A A6 C7 F1 7F E9 95 82 DE C8 F6 B6 C5 DC
 A5 86 0A F8 14 6F D5 A4 52 70 C7 B6 15 F3 5E 7F
 43 45 D5 2B 31 70 E0 0A 2C 17 F6 B6 B5 4B 10 AA
 9C BA 37 CD 44 21 31 C3 73 A1 5F 04 C0 86 CB 8E
 54 A6 AD 18 D8 12 EB 90 F5 70 62 3F 6D F8 E1 7A
 1B 54 71 03 63 D5 FB 40 58 16 64 AA BC 5A 9E 4A
 D7 A3 15 F1 11 E7 F9 74 E3 19 27 22 0D 9E 39 7C
 AE BB 9F D6 F2 AB B1 9B 41 A5 1B 88 1D 6A EC 71
 18 8B 5E A6 0C 23 6F B8 15 1E 32 A8 C7 56 88 3E
 22 BB FE 87 08 74 6E 9D 27 54 73 27 96 B6 80 4A
 AD 5C AC EA 89 BD 2B 1C 10 73 86 BF 3D C3 98 EA
 43 16 2E 8B C5 1F 79 BF B1 C4 43 D6 AF 74 4E F3
 4E 51 07 74 1A 8F 3F A4 2C 53 FC 56 5E AC 7E 5F
 0A E7 1A FE F0 7B 40 1F 99 2F A5 45 08 60 3A 5B
 81 BE EE 21 E0 C8 FC 7F D1 E2 C8 9C 2F 98 43 5E
 C5 43 28 AB 1F 57 C3 50 A3 E0 DD 9B D4 6F BF 48
 EE 6D A7 0D EA 2D DA 43 47 66 E1 F2 92 0C 0F 74
 86 0B 05 FE F6 63 36 2C 40 23 40 6C 28 92 A9 49
 34 9A 80 C4 78 75 DD AD F1 25 E8 34 08 C5 CC 95
 D0 C6 4B 46 8D 2B 7C 6C 88 A4 33 16 E9 66 28 5E
 D4 FB 66 40 88 92 72 0A AC DF A1 74 66 B2 F2 CA
 AB 5A 62 83 D6 26 5D 3B 9A AF 33 42 87 18 97 33
 99 40 3B 1F F2 E7 BC F9 63 86 AF A3 06 E4 70 74
 E1 C0 8F C8 04 4A 2A C9 D8 45 30 33 C1 F8 E5 DF
 1F B2 C9 2B 9B CB 2A AC 1A E0 2E 73 6A 47 19 9E
 79 BC D0 0D A8 BF 6E FD E9 B4 8A 98 EE 84 8C 41
 A3 B3 52 FA E7 D1 29 EC 35 2F 75 58 88 12 DE 58
 C8 71 B8 48 B4 B3 50 BD FE D3 A5 56 0E F1 DA 5F
 57 00 BC 0A 87 94 DB D8 5F 9B B8 B0 F1 69 3D 20
 9E 0C 01 89 DD D2 EB A5 C4 1E 41 D0 4E 3D 6F 2B
 7F B6 2D D0 69 A8 0D F6 F7 E8 9B 29 B1 3C B6 BA
 BD CF 88 4C 70 D1 0A 88 D1 5E 5F 39 BA A1 B4 B0
 CD 43 17 B6 47 51 51 64 DF 82 BB BD 15 1F 7A 3C
 A5 C8 7E D5 B6 E3 C0 03 E3 B8 D3 FC 74 CC 67 13
 85 D1 DD 0A E1 B0 26 4B 2F 1B 58 C0 C2 5A 9C E2
 BE 65 E0 97 4B 66 5F DF 1B 01 74 5A EC 3E AC 23
 AA F4 DD BA C4 11 AB 17 8D 84 78 6C 3A 51 15 0A
 04 C7 44 BA 02 5D 32 15 30 00 D0 EA E9 5C D0 66
 6D 56 19 C3 A4 9D 65 6A 87 72 CC A5 19 17 04 9F
 31 5A 01 52 3E 74 A8 88 A1 75 34 0F 58 5D D1 31
 9A 14 3E F7 CA 1C B3 BE 55 45 93 9D 58 73 33 8F
 EB 32 08 CA EC CA B9 E1 6A A2 97 85 2E B6 D9 3A
 C1 D4 6A 49 66 DB DC 07 23 91 B1 66 F7 06 B0 F9
 F1 16 68 F8 BE 68 8B 1B DC 14 BA DF D4 38 AD C8
 23 02 EB 85 2C A6 E4 A6 BD 5A 07 4F 2D 56 32 F0
 7A 28 B1 40 48 81 FC D9 88 91 FB A8 7B F6 DC BE
 54 42 A3 67 F7 13 BC AB EE E9 9B B1 BD A8 51 A5
 5E 96 51 FA B8 E3 DD 20 C6 0E 88 86 13 8F D8 69
 EF 1D F4 17 9D 63 50 31 33 BF 75 77 61 57 94 D9
 C9 37 1A 26 29 08 D5 4C C2 16 B0 71 CB AB A3 88
 46 03 8C 23 10 26 02 5A 10 D9 78 88 9F CA FD 70
 FE 69 C1 A0 5F 61 58 52 09 38 0E 2B 11 48 BF 8F
 97 F8 FE EF F8 49 28 4A 46 58 80 0D A8 FC E6 80
 AE 46 9A 8B 74 A9 AE 3A F6 B8 09 24 B1 AC 6F 0F
 20 78 70 13 15 96 4B E5 8F D1 D0 1B C8 BE 65 AF
 0A AE C8 D4 F1 D9 A6 9E 01 01 C9 95 4F 16 08 37
 43 92 33 7C 04 BD 27 26 F9 85 A9 45 2F AA 7C C6
 1B C9 D8 08 D7 79 FE 43 1C 98 EF EF BD 6C 05 2C
 9A 64 AF FA E9 31 D6 9E 5D DC 73 E8 23 0E 6D B1
 9D 9E A3 30 A1 86 98 65 BC 33 29 FF 3C 80 84 4F
 37 55 10 CF D4 3B 54 82 C9 6B 6F 4D E1 91 B0 E7
 6F 4E 68 EA 9C 6E 17 A7 DE F4 2A BD 61 CA 17 85
 0D 3C 12 FA B3 89 68 2E 71 DE 28 BC DE 45 3A A4
 55 03 8C 6C CC 21 0E 22 F2 7D 49 26 64 50 18 8A
 03 BD 7F D4 77 C7 8A 72 39 6F CF 84 1B 4A 40 CF
 CC D1 E6 C6 0E 14 85 9B 64 10 C1 AB F0 22 FC 42
 A8 43 09 9F 25 B1 1C 81 08 5C AE C0 6E 3A AC 77
 13 E5 68 59 9A 07 6A 29 E7 19 F9 04 DD D5 BE DF
 FC C4 76 A4 C3 ED 7B A8 11 98 5B 7E 3E D4 82 3E
 F2 33 7B 7B 40 A1 3A 31 FD 42 EE 9D D1 4A FB A8
 E5 BE EB 02 3F 2D 48 43 FA 64 18 FB 4B 62 DE 01
 4D 7F 38 BB F6 83 BB B9 64 1E D5 C9 13 2B 01 33
 D0 D8 C9 CE A0 0D 7D 0A 9A A8 79 DC 32 B3 21 F4
 A8 DB B4 29 DE B0 D6 34 A6 1B 45 FA 32 87 00 F1
 78 FF 9E 1B 86 18 2E 32 7C C4 A9 2E B7 6A BC 0D
 FA 08 E8 AA 09 FE 96 33 0E EC 32 F2 07 E3 A1 05
 BC 8A 1A EE C9 BC 7D 35 CB 1E 16 85 78 97 63 50
 05 69 83 C8 77 B2 E9 3E 8A A5 EE BD CF 09 08 94
 05 BD 33 BF ED B1 5C 14 97 73 91 54 40 9D 44 A0
 0E EE 45 DE C4 6B 48 26 2D 89 72 F2 E3 3C 43 1A
 AF E9 FF 2E BF 2A 2E 82 C5 27 27 A0 96 C3 18 AA
 10 72 02 11 EF 14 DE 1A 43 56 05 4B 32 13 A8 09
 DB 09 4F B3 9C EB 2D 7B DF 0B DB EC BE 77 41 B0
 99 16 87 8C BE CD BE 32 56 7C 2B 6B 75 44 67 04
 AF EF 16 86 F7 FB 01 C9 AD D3 46 F6 D6 19 BC 38
 80 DE 88 90 54 32 3B EE 4B AA 51 07 6D 6F 48 6D
 A9 25 0D 5C BF 9E ED BD 29 62 D0 12 C1 9B 0A 3C
 76 80 CE 1A 1F 17 9B 2E FD 2A F8 CE 66 5D 02 86
 46 4D D1 E0 06 EC AA 24 89 4B E2 AA CC 63 D1 BB
 30 EF 02 99 7A A2 98 6C 8C DA 36 6C 4F 8B 1E 43
 7A A4 2C D3 E7 66 79 E1 B5 74 98 74 9A 9C 35 32
 FD F5 44 57 C3 3F D5 D8 76 EA AE 79 D9 1D FD D7
 6E 0B 5E 11 F7 A8 14 C8 7A 28 55 63 B7 EA B8 99
 58 74 D8 83 7F 55 F1 C5 50 17 83 1D 82 B7 39 A9
 50 5B DA 9E A3 0C 96 A5 F2 96 E8 39 8F 38 5C A0
 A9 E6 2E D6 F9 02 36 41 1A 17 15 C1 88 CE D2 17
 0E 4A E1 98 DE 93 D3 36 CB 18 36 4B D5 7A B6 28
 6E 52 76 CF CE 66 BD CD 59 3C 38 E9 7C 46 A6 31
 F9 73 43 4D 1B CF F3 93 9F C1 B2 58 2B C2 0F 1A
 DB 77 7D 39 FA A9 BE B2 C2 CC 24 29 B8 03 1A F6
 11 21 50 4B DE 9A 34 8D 09 7D A2 26 91 18 4C F3
 F7 F4 8F DB E2 8B 72 62 78 1C EC 1A FD E5 67 A5
 CB F2 1D BD 27 6A 56 17 EA 6B 49 AE 53 8D C7 33
 74 C0 6C 11 48 36 7A 89 B8 BB DF 89 95 FD 3E 78
 A8 47 DD 52 D1 85 17 EE 29 A6 92 08 F5 5A AA 78
 DE B7 07 45 A4 7A 3B 6B 6A D7 4E B6 C0 1F 96 97
 F3 09 E3 52 29 F3 02 2A 5A 26 9E 13 29 B0 59 44
 A0 BB E5 04 02 63 09 FA 33 D7 98 17 4A DA 37 57
 0D 97 44 C7 BD 22 60 1E B9 3F 3D 16 82 B9 52 1B
 DA 31 BB 8B 7B 38 1B AD 4C 8D 3E 40 2A A7 B2 0E
 8A 00 CA 46 5C 7D 15 7C 58 0D EE 2D 4C AF C1 0F
 3C ED 87 DD F4 DD 34 A6 4E F9 89 2F D3 62 60 26
 D4 30 68 B8 82 31 5B EA 88 E5 53 80 3A AE 9A 75
 6C 01 1C 21 74 E9 80 C7 F5 5E 5A A8 69 F5 E3 55
 A3 67 0E AD 02 F9 A8 5D B7 71 FC 09 61 DD 96 B5
 34 44 77 AA E2 B9 DF 77 05 F1 EE C8 E6 55 AA E6
 91 9F F1 59 BB 44 FE 76 F1 19 C0 45 BC F5 B4 62
 FA FA 63 36 5A D7 06 FE A3 BF 59 57 46 30 65 FB
 46 15 A4 F7 05 09 24 CE 28 D7 5C 5E 77 8B 36 DF
 2F B5 63 9C 91 41 93 23 CB D3 F2 F8 73 B4 B7 F6
 4B BF BB 7F 9A E2 59 39 AD 01 AD 1F 09 4A FD 27
 02 48 43 14 77 59 19 5F A4 D7 D2 E9 B2 15 82 00
 A5 FB C4 1E 94 83 69 1F 61 3F 92 C0 B9 2E 2F 8B
 76 EF 21 E9 AB F6 EA 3B D1 15 BB BA 7D D4 3E 56
 49 29 44 4A 97 00 85 36 3E 33 63 F7 FD 73 73 87
 E2 69 29 1C E3 34 12 2F 87 B0 2B C0 BD 66 76 B1
 50 51 60 DE F7 C5 8D 1D C5 92 69 75 11 88 64 01
 B4 8B 2D 5F 26 EF 8E 97 5F CB C2 0E 00 E4 7E 4C
 B9 FB C7 49 B9 21 D6 4C 67 FD C2 5F 96 D6 66 B5
 53 CE CF E1 2B E9 17 FE 30 60 71 44 F7 04 48 98
 82 EB 2E D9 51 9F 8E 19 EF 45 87 B7 DF 51 6D 55
 6C ED 68 D7 82 FB 10 E1 15 8C E2 88 3B 42 16 B7
 91 CC A2 49 15 51 0E FA 8E FF 1A 84 65 54 9E 78
 FB 37 88 07 7F 0A 13 73 76 E0 B6 D5 5B E7 43 7E
 2D 35 62 06 43 29 7E 62 76 80 77 FA C5 A2 09 21
 2E 72 7F 1F 87 10 08 4F 79 BF F9 A9 65 64 B0 8E
 50 6C 45 9F F7 40 39 46 9E 8A BF BB 67 CA 20 FF
 5E E3 3E 8B 34 0A 44 AF 96 B3 BB 5B 99 78 72 0E
 9C C4 2C D0 CD 82 B1 26 18 AE 59 62 57 08 24 09
 5E 2E 87 A2 D0 BE E1 C7 AE DF A3 08 1C 06 82 C7
 BE 5B EC 4D F6 F7 DF 1A 26 F2 FB 2E 54 46 96 07
 44 5B 3E 73 E3 3E 34 00 54 14 9B 49 58 92 BB 0F
 D3 7A AF 8A 84 EF 0A 5E 27 42 80 A0 FA FB 22 45
 77 95 FE 77 DF 4F 42 E7 17 3F 6A 62 A9 00 CE 55
 39 A8 ED 5F D2 3A 89 4A 10 D0 25 7B C1 31 8E D2
 EF BD BF FF 21 4C 8D 3E 18 9E 70 1E F4 25 09 23
 7D 6A EF 09 1D C7 B2 87 0D 34 76 C8 86 CD C3 0B
 8B 88 CF 39 61 09 FD A0 D8 67 E0 25 DD 48 06 40
 B8 E7 FE A3 A4 7E 29 0B 7F 42 7E 1C BE 7A 80 F5
 CF 0A 72 82 18 A6 64 B1 0A 4F E4 3D BC F5 E3 15
 55 9D B6 FC E1 AD CB CB E4 2A 8B 96 E5 B1 B0 0B
 03 93 CA 19 51 7C AE 32 C6 8A 25 64 66 59 E7 28
 00 34 44 A7 36 7A 80 07 67 D3 25 CF C8 F8 A5 39
 CF EB 61 9E 35 8F 7D 1B 98 00 A2 65 8A 0F 2C FF
 72 1F FA 18 68 26 19 E0 3E 7D 87 7C 4A 08 F5 C4
 34 10 AB 91 BC D8 B5 51 CA AC 4F E3 1D 2F 76 16
 64 E6 79 33 87 F9 4C 07 23 63 F9 11 CD 15 4B BA
 17 67 8B EC B2 AA 59 F2 EB 79 0F 6F EF 88 90 4F
 3C 1B 86 D0 0E A3 5E D0 74 E2 38 92 13 36 FB 9D
 11 D3 5B 32 0C 5E 98 77 1B AF 23 CB 77 7D D7 CF
 26 26 17 2D F7 09 C6 81 A1 0D 54 0F 18 50 FA 1D
 E1 25 C1 D4 71 39 31 95 50 98 C0 48 38 E3 67 F1
 3C 26 6B 44 52 B2 08 38 B6 90 27 EC AE C5 97 B1
 F4 84 3C EF 19 1D C9 C1 51 D0 55 55 11 F1 58 21
 8C F7 26 A2 9B D2 60 5F 38 04 C6 75 2A 30 38 EB
 55 48 C1 EC 0D 00 D2 76 51 0F 4D C8 51 DF D9 D9
 B2 96 1C FD 68 F9 66 DF D2 A6 D8 30 21 C1 AB 45
 E3 5A 34 42 BE 63 F1 12 E3 DF 84 E4 BB 9D FE A5
 7B 4A F0 67 B3 AE CF 4E B6 23 1C A9 51 9F E0 84
 DA B7 74 A7 CD F8 3F 9F 21 6C 48 A9 07 BD CE 0D
 CD B8 C1 D7 99 3A 88 6C FD 97 37 9F 3E DD 0D AE
 CA D6 EA 4B 51 AF 36 4E EE 6F 6F F4 00 D0 CA 73
 D9 B2 85 1E BD 44 3A D5 C2 01 FF 84 92 6C 67 E4
 F2 E3 D3 25 9E AC FD 2D A2 47 6D C0 AC C3 A5 C1
 F7 ED 29 CD 91 D5 D5 29 D1 E0 F7 21 71 3B B9 EE
 4D F5 0A D4 7A CF B7 1C 66 B1 53 25 9A 35 4C E7
 E6 8A 99 87 EC E6 E2 11 BC 26 35 CD 37 FF 33 E7
 FF 5D C3 F5 94 64 38 BA F4 D3 C1 73 DE 55 BC 18
 2E 36 34 07 E3 62 C8 5F 0D D3 92 BE 1D 01 F4 4A
 42 04 90 E2 2B 53 A5 75 0E FC 30 EA B9 FD 8B 58
 6B 55 D5 73 86 1F 88 7A 89 47 E5 CC 6A 1A 58 9B
 31 A3 D2 9A E8 A1 DA 85 91 6E D7 44 BA 74 08 6D
 27 0B DA 0F 58 3D 2A AD 9D 7B 95 FF D6 E0 76 7B
 51 C1 0A 04 88 F1 E3 C7 20 A9 28 62 36 70 33 A6
 A8 09 AF 82 E3 20 07 EB 3A 94 B5 A9 18 4B 21 E8
 FA CA CF CA 0D 39 DA EA 83 C5 B9 98 DC 7A CD 6C
 58 B3 6B AA 73 02 2E 02 4A C4 8D 5D 3F 81 02 3D
 08 F4 10 98 24 07 65 3D 17 7B E8 1A CE 05 A5 E9
 AB 73 FF 6D F6 EC 44 CC D8 79 AC 56 E8 CB 1E EF
 D3 94 AE 92 66 40 09 8F E4 6D 20 1B 4A 62 10 D5
 12 55 29 3F 37 A0 D8 BE 74 AA C9 F2 B7 A8 08 A9
 38 18 C0 E1 E0 66 F2 33 95 A7 BE 7B 8B 5A F6 F8
 B8 78 14 C6 62 B5 63 32 A3 EC B7 F0 20 E7 6F BC
 22 BE 75 EF AA 51 33 57 66 BB 1D EA CC 9C 32 08
 3A 52 33 E0 C6 B6 DD D5 E6 E2 ED F6 EA B1 95 6D
 E9 88 82 F7 1D 2E 1A 87 E7 5E 6A 21 BF 7C D1 AF
 0E 83 DA 12 57 60 9C C5 9E 11 53 8F 95 E6 D9 E7
 9C 4A 82 42 C5 C9 7B 2C B0 12 74 06 BC E2 83 C5
 75 2D 81 09 E2 8D C6 1C A7 1B 62 FE B6 35 38 F5
 A4 8E 2B 95 65 0E 2A 37 E2 1A 8D 7B CA 0A 33 97
 1E 7F 7B BF B5 53 16 92 0D 84 70 F0 F8 9E B8 8A
 28 8A 40 55 B9 E3 C0 75 61 04 8D DA F7 54 E6 F2
 B6 50 BB FC DA 33 35 21 36 78 6F 47 01 78 C8 D8
 A4 2F 60 AA 5E 30 7D AB 49 19 52 F8 8F 12 D4 BE
 66 4A 4B 1B DD C8 8E 4C 8B 80 98 6C 60 27 CB 97
 2A B5 CA 93 DC 35 4E 13 F4 7D 4F 6B 4B A0 79 2B
 E5 E6 E2 72 74 FE 88 FA DE FF C1 47 7C DD A0 37
 B5 BC 93 C5 89 D6 8A 25 C8 AD 58 3B 6D EB DC E2
 D2 8D 12 E1 AA 24 46 B0 48 9E 5A 6B DE 58 6F C4
 3D 7C 21 9D BB B2 22 76 61 0E 70 47 9E DE 34 3A
 3D 2F 8A 34 66 4E 51 77 92 7C 25 40 6C 4E 6A 35
 32 65 8E 3E E8 12 1C 94 63 91 DF 4F 76 34 ED 38
 7F 64 6A C2 53 F8 61 C4 F4 BF 11 56 CD 6F 0B 1F
 EF FF 02 06 71 6B B7 B6 78 31 31 8A CF B0 80 25
 90 E2 45 42 80 0F E1 34 DE 8C 86 A3 72 29 2B BD
 C7 72 DE 30 F7 06 E3 A6 6F F4 7E 29 F0 A5 AC A5
 0A 21 19 0F 27 58 EA 8C B5 D8 CB 28 DD 02 9C 80
 1B A5 4A 0B AB 10 B5 0C 53 2E F6 02 D7 99 04 BF
 9D DF 3A 05 9A 31 FD 7F 09 17 44 5D 7D FD E1 90
 AD 09 9C 93 76 11 21 B2 CC 14 A6 83 A5 23 5E 56
 95 7F 4E F2 FB D2 F5 C3 F3 72 C0 AF 10 80 D9 68
 DF 3A BE 40 5C E7 30 00 D8 D0 CE D0 3D F5 88 3C
 75 1C 5A 56 85 C3 69 37 E0 33 CD 3C E5 7F CA ED
 B2 67 37 2B 60 82 49 AB 24 85 96 22 03 14 EB 77
 7C E5 DF DD A2 7D 99 16 30 DD 79 1C 6A 6F 90 7A
 58 5C 81 0B 52 9A 77 31 B6 DE B3 9E 21 BE E3 15
 89 71 0D FB 4B 81 07 BC 72 2A 60 6D 64 B2 C7 53
 DB E1 82 E9 49 6C 43 65 B8 D3 38 21 BE B2 67 D5
 37 35 C5 B3 68 A7 E6 B5 32 0E B1 C0 8D 75 C9 E6
 EA 8F 9A 18 0F CC 7F 21 8E 0C 9A 91 DB 45 E1 F3
 B4 C6 7B 84 7F 5E C9 A8 6C 6D EF 16 A5 AB EA 68
 2A EA FA 3B E3 7F EB A6 93 40 E7 4F C7 D1 D1 44
 35 AF D8 D2 C8 08 E5 04 27 FE 97 05 7E AF 29 C5
 25 17 81 76 9D C0 D5 99 04 A4 64 0B 57 34 C2 1D
 BE 5D B8 70 A7 18 AD F3 F9 40 35 C6 55 0B 2F 45
 86 2D 81 BC 34 59 D0 3C FB 01 8A 35 3A 87 A5 5A
 45 F0 EF DD DB A9 C6 F3 B0 E9 97 F5 8F 48 65 5A
 C6 55 20 DB 8F 39 74 16 FD 9E 2D 25 59 EA 5C A6
 3F 3E DE AA 80 49 C1 A4 81 83 4F 26 54 81 ED F1
 FD AE 3F CE F6 7F AF B6 A0 FE 68 86 8F 68 D5 70
 C4 69 9D 8E 20 0A 81 0B 6A C0 2F 40 54 32 24 AA
 9C C6 F7 4C 37 19 27 79 5D E5 1D 5F E8 67 4F DF
 46 63 8C 06 F6 59 C7 5D 6C B8 5B D1 6B 1B 65 F3
 64 04 4D 97 58 52 EF DD 5A 1D 87 4C C5 4E FA 5A
 B6 30 27 95 7C E3 62 2D CA 2D FC 69 C5 44 0F 1E
 7F 51 A9 77 65 65 C6 A2 3C 7A 97 82 6E 30 E8 F1
 6A C3 43 B3 74 BD 10 96 B2 C0 BD 16 86 68 17 09
 2D BD 76 F6 FD E8 24 CF 9D 34 93 27 27 D0 FE 02
 0C F4 BE 03 42 35 99 5F 4E A6 2E A8 4B 2A 4A 1F
 0E 3E 6C CF 07 94 68 9B 69 FC AB C6 EF C3 03 16
 9C 15 BA A2 4C 29 AC B0 BD 39 F7 39 86 E5 59 BD
 0D 0F 34 5D F3 CD 71 FE CD 09 DD F1 6B E5 2B 16
 26 41 E7 43 7B 8D FF 65 EE 32 96 4C A0 F9 A6 1C
 D8 A4 26 65 34 87 81 0D C6 DD CD C5 22 A0 3B 3E
 DC EF C0 C3 30 34 03 AF A2 2B 2D C2 F9 3E B8 CA
 41 92 76 77 59 2A 7E AF CD A8 56 76 4B 57 6E 68
 B9 1B F7 73 A5 C4 AF 78 94 14 80 99 69 D0 68 62
 B6 C3 B7 18 C6 15 E1 EC BC 44 70 4D 80 4B A0 BF
 82 0C 84 3F AF C1 83 1C 82 2B EC B1 9B 99 5D E5
 E0 DA D5 B1 33 40 E8 D5 A3 C8 7F CC AA 8F 7B 51
 D5 6A 8D E8 07 FF E1 65 19 2E CD 7A 4E 6A 8E D0
 62 BE 6A E5 3C 56 5A 18 80 0A 97 81 0D E4 D0 C3
 08 88 1B 9C 53 6C 35 67 D5 C0 0D 3C E3 2E B4 5C
 A7 34 41 7B 18 20 EF 38 0A 1F 7A 14 CD 20 61 4B
 A4 67 2D 1C 10 84 1F 5C AF 4C 2C E5 64 5B 8F 36
 A9 FA AE 06 C2 14 C6 B1 8F DA 86 46 6A ED 0B 09
 AD 8B EA 9B 91 7A 01 E4 96 34 6D A6 B4 70 C6 02
 04 22 5F 96 6E B3 C3 BC 38 39 11 E4 C9 71 DF DC
 36 94 EC 03 B0 6D 37 8A 1D 02 98 20 EE B7 FE B0
 4E 6D 7A 6E CD 73 25 76 7D B9 F1 4C 1B C7 24 B5
 CB 7C 8F C4 90 F9 43 05 D1 B6 B6 C1 46 C5 02 00
 62 97 52 A3 72 60 42 F6 85 A2 31 1F 32 DC 6C E7
 A4 14 34 B8 D1 81 0D 64 F1 80 13 77 D5 07 BC 83
 85 6B 74 72 AE 24 92 E8 A0 3E 90 C3 C2 B2 71 EA
 F6 5F F2 E0 13 E6 6E E0 41 E7 94 CF 0D 71 64 13
 63 57 65 F6 BA 8C 40 B5 A0 D8 B6 98 C8 95 2C E1
 60 03 00 8C 8F AC D6 AC 41 9B 08 F2 D1 D2 57 22
 32 BD 76 62 44 D7 07 D2 02 B4 90 08 CB 06 B1 FA
 F6 6F 92 CE DE 67 00 17 D8 24 B1 35 04 25 E1 A3
 CC B4 0E 3D D4 64 69 38 51 FF 50 D0 B0 C3 B3 B4
 1D 86 FC 2F 20 A3 E7 72 93 C6 DD A7 8E 1E 6F EE
 0B 18 9C F6 BE D3 19 D6 87 90 91 28 FB 4E FA C4
 E5 16 00 52 98 46 5A 1A 8B 9E 62 6E 5E 88 5F DB
 49 36 E6 D7 A7 B0 5A C6 7C D1 D7 18 52 B4 66 67
 63 EF A5 21 05 84 EF 0A A7 CB 33 14 3C 52 09 E0
 C9 D2 54 55 A1 2F 02 AF FD 3B A7 77 2F 8A 9A 21
 90 C5 82 EE 3D 60 A0 DD 31 4C F9 77 20 DE F4 06
 7A 31 43 89 6C BC 50 DA A7 4D 26 D0 C5 32 01 59
 B7 82 F7 1A CF 6E B8 43 20 39 89 79 FD 06 E9 1E
 2C D1 59 E4 2E 66 92 CD 11 F6 92 DD 1B A4 3E 88
 B3 77 D4 6C 93 32 B9 BF 8D E4 AC 15 94 0D D2 72
 40 25 05 35 A9 91 89 DA 70 56 E3 A8 AA 05 0D 80
 91 F1 D9 AA 8C A1 A8 AD D1 EC D3 A5 A1 8C F9 C5
 0F 7A 6C 8D 0C C3 04 A5 89 75 C7 BF B1 ED D4 E0
 56 73 8D 2A 88 C9 AA 09 5A C4 EA 88 E8 B5 EA 44
 97 E0 73 FE 73 CD 79 ED 87 9B C2 92 92 43 FE 0B
 12 EF BF C0 71 41 31 3B FB E0 DE 55 E8 B6 A8 1B
 CC 53 B8 1B 08 8C 26 C2 47 45 8F 7E DF F3 25 8D
 1C 5D 34 57 2D 6A 20 54 24 53 D2 DA B5 41 53 97
 13 5A D0 E3 A2 2C E1 FC 9A 3B 04 0A 59 F4 0B 42
 4A 18 7E 43 8C FD CB 6B D0 3D BC 0B 59 C9 98 40
 F2 64 78 C5 46 AC 54 39 35 BD 45 B1 2A 27 4D 7B
 8B 81 C6 9E D4 C3 C6 67 2A C7 4A C9 DF 03 18 01
 AB AE 13 A8 37 B0 FE 03 9E FA B3 C5 E4 AD FB 42
 80 F5 53 34 4D 4D 33 ED 03 05 1A EA 07 EB 75 29
 D8 85 C2 A0 56 A7 F5 C8 5C D1 F0 FC 1C 7C AA 3D
 4E F8 E3 15 6E 4F D0 41 64 CF 08 92 EA C0 F7 C9
 F0 3C 38 90 D8 6A A6 7D D2 5A 0E F4 88 C4 33 70
 B3 A0 14 56 0C 79 C1 32 DB A0 6A 95 61 FB A3 64
 04 11 B0 19 F1 BD 8B 41 7F 92 B3 09 A4 77 5C B7
 4B 55 A5 32 E4 F6 94 99 A0 62 18 EF 06 AD 57 55
 56 42 F2 CB A3 94 62 54 45 F4 42 91 94 E4 14 0D
 36 8E F9 D8 E9 A2 78 06 BB E5 96 E1 CC AF 57 EE
 F3 01 36 E9 64 02 D7 E6 44 77 29 70 2C A9 D6 60
 45 E2 A8 92 12 89 F3 C4 71 3F 35 EA 82 AD 77 CA
 05 F0 E2 4F B5 F7 46 C3 E5 FB 47 A4 F3 1D 20 B8
 AA 36 3A 00 8D 4F 50 AA DB 0F D2 BF EE 4A 95 AC
 C0 A1 26 6F B7 7F BC 35 60 54 0A 7B 54 C6 C3 CC
 2E A5 9D 3B 62 34 FC CA 35 F6 C2 03 9F F9 1F 2D
 0E DD 34 E6 C9 8A D6 E1 8F 16 F8 4F BB 24 9B 74
 97 B1 52 B1 F9 3C E4 91 6F FD C1 0E E3 F3 E0 F8
 0B 1C D0 AE 87 71 DF 5D 98 65 1F 97 20 42 AA AC
 25 F0 FE AB 0F DC 4C E7 F7 E5 B6 79 2B 6B B4 56
 30 43 9E 18 E0 E8 B4 35 17 79 88 E2 EF 27 67 B0
 7D 55 47 BD F3 A2 5B 9C 82 E0 EE 4D 94 9F 2E 81
 06 61 4B 53 9B 64 AD 60 24 4D 9A F6 B3 21 F8 E6
 29 23 30 F6 6F BB ED 08 B0 F4 58 81 3E DD 49 19
 64 FB C2 89 A6 89 7F E4 0A 8F A5 1B 5F BB 48 81
 4A 57 9C 9E CF 76 CD 43 57 1D 05 86 E8 BA 39 6A
 E9 7D 7A A1 D2 16 89 1A 10 3B BE E3 A3 B1 95 FA
 3D E7 A8 12 F0 9A 60 39 EE 3B A1 A4 CA 10 95 99
 4C DC 88 34 61 6E CD 88 0C 2A 74 C9 F9 49 27 06
 89 2B FB 9A 63 B0 D1 7C 5B 16 12 E6 05 A6 45 C1
 95 A1 55 73 E5 1C 37 5F 33 BD B2 A7 2B EF E9 A3
 18 E4 F8 97 02 48 69 D0 3D 44 09 90 B9 4A AD 67
 67 C6 2A 12 8E 1A 2A B0 37 36 56 F9 65 7A 83 51
 06 23 F9 0A 02 F1 9E B3 DB 6B 07 5E 46 4E 64 E5
 D1 F7 99 2D 7A 3D D8 B8 3C 95 FC 3A 76 CB 27 51
 95 EE D3 F4 1E 7D 1C 25 3B 80 43 61 76 93 9F D2
 49 64 A9 0F 95 88 1C 6B B5 00 9B A7 47 20 CE 3F
 64 36 5B 8C 9A FD 45 64 9E BF FF C7 F7 16 E1 31
 6A 53 D3 8F 8A CF 68 88 C2 24 E0 FB 8B F8 C3 F6
 3D F9 58 C5 7E A6 09 89 F5 10 C3 4C 53 94 30 93
 BF 17 B7 7D 1A B6 AF 74 DD 3B A6 7C 72 78 91 AD
 C3 19 02 10 61 03 C9 B1 0A 9E 01 68 EA 45 90 B7
 BB B9 0D 46 91 56 DE 55 13 5A A7 C9 F6 FF 03 42
 2F 58 0B C3 F5 08 32 C7 BD 1E D6 96 62 E3 CC E9
 5F A4 30 61 55 1E 57 5C AD 2A 2A 72 A4 24 D0 18
 00 D2 D7 3D 9B 46 8A 81 DF 10 E2 7B 66 27 76 5C
 43 9C 2D B2 33 6F 61 9C 40 BC 81 FA 25 A3 80 43
 66 F4 6D 78 4D 20 E3 10 F3 36 3F D1 9D C9 09 76
 11 52 50 C8 82 0E 6E 20 A3 29 C6 95 56 0A 76 39
 75 F8 E4 27 1E 94 D8 07 75 E7 19 26 57 21 D9 3F
 ED 06 DF 13 E0 C8 41 31 3C 44 7B 40 A5 5E 7B 5F
 B3 9D 38 0F 97 1C 28 7D B0 D1 4C 10 4A 65 20 EE
 E5 3A 70 66 6A EB 99 3A 2B 02 23 FA 0D EC 4F 43
 11 55 88 41 87 26 98 0E A4 37 FB 4C 24 0C C0 63
 7E 4D 00 43 0F CE 29 DB 2A AF C7 57 15 5B CC A0
 05 7B 2E 4C 39 E2 48 81 32 AF 4C F5 93 EE 6A 20
 A7 58 31 ED 9E D2 51 1F 0C AD EC 73 F5 30 92 E6
 7F CB A6 CC 73 0D 9D C2 81 C4 A4 AE F5 B5 3C 7C
 F1 31 24 15 56 CB E5 D7 6D DA 71 78 70 6B 1D B9
 19 E9 C2 E3 CB 24 6F 58 5D DC 17 70 B0 C9 12 CB
 75 5A A5 6B 2F 6D 97 86 D0 E3 DF 39 03 7A 6F 3F
 63 66 53 75 A6 98 97 B4 A6 ED 62 EA 0C B1 D6 9F
 7C 8F 03 DD A6 AB 77 FB 9C 92 FB 8E 8A 26 91 00
 BF 95 28 F1 56 83 73 79 3B 46 87 8E 94 98 DF DF
 1E 2C 9F 58 8D 54 D2 4D BE 2C 57 30 7A E7 58 2E
 90 63 8A 0A A9 19 A9 BF 80 DE 62 BF CA 16 16 93
 AB 5B 54 EB DF C4 D3 3F 8E D5 02 4D EF F5 FD 52
 7A C2 BB DA B1 96 E9 D1 AB E4 7C 21 B0 C4 B3 0C
 63 FA B0 6D EB 28 F3 37 03 54 F7 F8 DC D9 64 39
 90 68 48 56 3C 07 8B EA 58 CA 94 18 44 C4 CE 00
 34 FA 20 B5 A8 54 4B 0B F9 E5 4B 2D CC 2B 90 FB
 3B 32 89 CA 33 54 DC B7 0C 5A 28 C8 F1 8B 2C 57
 7B E2 5E B2 85 34 40 3A 74 15 97 DE B8 55 87 B2
 E9 8B 6D 88 BB 6F 31 F3 B1 3C DC 66 46 A1 D0 AE
 64 F5 E7 B5 4C A6 1C 38 55 8B 72 40 C2 33 AE E2
 24 9E E7 FD 38 30 07 71 99 72 02 48 2A 22 A7 03
 5A CA CE 13 EB 68 72 68 2A 99 D5 C0 3D F4 89 86
 68 95 05 CE 98 87 D0 53 46 4B 64 44 35 2A 6A 37
 34 6A 47 EC 8F D6 2E 60 1A E0 41 1F EA BC FD B1
 FD CE 3B 74 CD 67 67 0B 64 9F 1D 40 0B 0D 0E 51
 6D 4E C1 E3 AA 72 CE 2C 96 CE 46 F5 AA 9F 1B BA
 72 79 22 E1 EF 75 F2 42 6B D5 B6 C9 3F 4F 16 5F
 48 56 24 27 2E 4A EB B9 54 0A 48 15 01 66 10 E8
 65 69 AD 4E 0F EB 6D 94 B8 23 11 1A 24 10 FC 65
 48 F5 1D 30 E9 50 E9 9E 50 DD 13 04 D2 CB 85 0D
 C3 6E AB 95 80 24 4D 26 11 3F 22 DC C4 2C B3 C2
 8F A2 98 C9 51 4F 46 7C 6A 41 EE EB AB 50 96 B2
 90 6B F0 0E 6A F4 FC 20 59 9E A7 70 48 64 94 95
 E0 67 D4 6E DB 5F F4 FB 3C B9 56 E5 EC 94 B7 58
 9F 4E A4 0C CB BC F2 5B 90 89 3E 05 A5 6B 84 0C
 DE 81 4B D6 AE 35 6C 33 B9 DC 72 6E BD BB 94 56
 29 88 64 BD 4D 10 87 83 5F 16 33 84 D1 84 5F 9E
 86 29 80 2C CC B1 2A 42 38 70 0E D1 D2 8D 6B 11
 CD C3 BD 99 A1 94 EF 72 4E 49 93 21 BC E9 DA 54
 53 69 B7 A5 DF 72 B1 7E 65 DF 4F 56 DB 59 E8 0B
 61 7B 45 6E 17 8A DD 13 8A F7 FE 0C E8 0C 90 74
 E2 B2 95 AA 31 98 7B D3 1F DB AC A6 20 24 22 49
 B5 2D 54 C5 CE BC E9 D9 EB 8B 5B 77 B0 E8 60 E1
 1C C2 44 2D 7A DD 23 3E 5C 01 EC A8 63 26 54 78
 AE 09 98 F4 31 10 75 14 51 78 50 E8 D9 11 21 22
 F7 21 0B F8 B8 2A C4 2F E1 44 6A 7E BC 23 90 9D
 40 54 8A 20 4A D2 6C BB 34 3E CD C8 CC AA A8 AE
 B5 B8 20 41 17 24 E1 1F 94 31 94 4F AD A1 63 65
 73 F4 49 A4 54 DE 9E 53 EB A1 1F 6C C1 4A 3B 82
 5A 5C 3F EC E3 AB 78 71 3A 44 DC D4 B1 A6 45 BC
 D2 21 65 B3 74 BA A9 7D 2C F9 38 97 5E 6E 35 A3
 C8 0C 19 1D 0A B5 25 E5 88 A4 F3 EF FD F5 53 21
 8D EB 2B 50 AB 0B 46 B8 57 AB 45 4E 96 D5 D8 AE
 10 D2 1A B1 8B 16 CA 4E E6 31 F9 AC 84 4B 9D 30
 C2 72 1C 63 15 2A C1 30 FF 98 3B 44 4B FD 95 52
 7B C8 7C A9 29 00 3A BA 25 A1 A9 FE B3 D6 3B 03
 AF 11 A8 63 91 6F 28 AD CC 84 2F 4D 31 89 8C 76
 27 39 DB 33 C8 FB 6B 95 2C 3F 7C C3 24 08 52 64
 FA 5B D0 18 16 9E A8 03 3E FC 83 35 B3 B1 48 FB
 8F C5 8C EE FF D9 E6 26 7F 2C 7C A7 FD 97 9B AE
 8B 6E 94 3E 10 11 3C 39 F4 F3 16 16 61 98 51 8C
 E2 37 07 E2 9A FE F6 4A 3C C9 E7 86 93 B7 09 A5
 3D 6D BE ED DE 62 4A 5B F2 85 59 96 64 1C 5D 5C
 4D 5A EE 0B F6 08 0A C6 B2 58 DC 7C 74 52 4E 76
 83 5C A4 63 55 2D 7D 76 2F 6C 8E 43 9A E8 BA 1B
 A5 F6 3F F0 AA E6 50 6F 49 2E 9A 40 DB 0C D0 D3
 2C 15 E6 1B EF 64 09 B9 02 13 F5 7E E5 1A E5 9F
 1C 0F 8D 9B 6A 7E D5 DB 64 63 D6 42 DD 9F 30 FD
 81 52 A0 AE 2A FE 95 79 63 05 08 8F 7E F4 C7 22
 EE E3 2E 83 07 68 E9 BF CD D7 A4 3B 19 E2 4B 18
 27 65 26 25 3C F0 7F FA 9D A0 D9 50 4A 7A 7B F4
 87 58 8C F1 EA BE F2 1A E2 56 7E BF 5F FB 49 F1
 D6 BD FF 3D 2B A1 60 5C 1D 1D B8 DC FC 4A 0B 6D
 32 5B 2D CE 97 47 B4 21 A5 BE 97 A9 96 4A 86 9D
 3E 41 C2 B5 7B E1 6C 56 DE 0B 45 EF 7B 81 92 82
 5F 68 22 22 FE 41 51 1E A8 BC 90 2F 5A 04 D2 90
 ED A1 89 58 19 95 95 9C B3 BE AB 6E 82 9F 35 B9
 6F 26 37 77 3B 02 7D 38 AE 94 69 F4 9B DF CF 89
 2D F2 05 02 EB AE E9 78 24 CA 2B EE A2 91 A2 0E
 9C DA D8 7A 40 27 78 FB 79 83 34 93 AA C6 6A 62
 8E FB 07 F1 B5 78 1C 19 24 61 00 1B 84 97 69 C4
 A3 2A C7 5F FB BA 0A 0C AC 87 CF 05 6D 15 E7 F9
 B8 90 A8 65 FB D0 8B 30 1F 09 98 4F E2 C5 6E CB
 5C CF DE F8 CC A8 DF 03 DD 35 7B C9 36 F9 FC D5
 5C EF D6 5A CC D4 0C 0F 0C 60 9D 72 AE 3A E8 58
 66 90 C3 E1 60 3A 95 4C 79 CF 1A 4F AB 4F BF 3C
 CA 23 9C 66 C7 BE EC 47 26 4C 7E D0 DE 41 EC C6
 CF B8 25 F1 D1 CA C6 9A 09 B9 7C 95 BA 07 5F FB
 66 3E A5 05 19 0F A2 05 56 BB C0 3D 8E 5F 85 DC
 8E 3F 68 80 87 FE 40 CE 95 2A 3E 36 C4 AD BC A1
 F7 47 CF E4 A3 10 5B CF 8D D8 7D 19 0E B8 02 37
 E0 A6 CC FB 5C 60 A1 36 EF 9D D6 A8 8D EE 37 30
 C0 45 0E 67 B2 45 E4 C2 3D 4D 5F BE F3 E2 A8 8B
 95 FA 86 5D DF 7A 6B 69 DE 4E AB 02 61 A7 B4 DB
 7C 4A F9 60 E0 97 98 C2 89 23 AB AE FA F3 EE F2
 36 59 CF 38 16 92 B7 D2 17 73 4E 3B C9 95 90 22
 CA A0 5B F6 26 FA E0 F9 E0 18 2E 8C E7 F7 0C 99
 9D AA 16 22 3D A5 6B B3 F7 7E 5B 88 01 18 68 68
 EE 89 53 E6 78 A7 EE AD B5 1D EB 44 DF 55 15 AE
 FB 9B EE 03 58 7B C7 9E 15 D3 6E CD 30 0F 51 6A
 34 10 09 69 80 CA 1C AF 60 5D E1 8D 35 12 8B E1
 B4 3A 76 60 1C C8 48 C7 37 12 DE B2 58 63 6D DF
 13 8B 5D 58 DC 45 85 FE C5 A7 34 6D 2F 26 17 28
 D4 AA EF 83 CE CF 3A 6B B9 91 24 80 8B C0 28 FD
 CD 50 C1 04 48 5B 5C 65 EE BC 0F D1 F9 42 2F F0
 AA 1E F1 4D F9 36 91 93 17 2A 72 CF 32 F7 8C DC
 DA FF 08 A9 FE A1 72 E9 F4 B9 C1 BF 81 65 3D B8
 3E ED 6F 3A 33 10 92 23 59 BE 11 FE EA 1E 37 85
 18 5B F2 6D C2 78 0E 44 2F F1 FD E0 1D DC 90 6C
 03 41 00 5E 97 F8 82 FB 1B 86 A2 16 3E 82 C1 59
 DB BE 33 55 13 6E 21 01 42 07 B6 81 E5 41 E9 AD
 B7 FB 05 1E A4 A3 D8 07 0F A2 79 8D 61 A4 0C 4F
 6B A9 32 59 55 39 C8 3E 59 59 1D B3 BD A0 6F 2E
 7E B3 B1 F0 6A C8 66 2E 0E 5A B1 C2 07 2E AD 7C
 7C BB AC F6 17 14 E3 8D 7A F9 CF BB 65 1D 5C 72
 A3 B3 75 02 1F 95 B8 04 75 73 58 84 4E 17 8D 59
 17 8C 6B E2 41 61 F4 09 56 6E 37 A0 BF 8C B6 E6
 14 CB F6 72 71 0F 2D CB 5B 3C 31 4D 2A E9 BD A1
 06 28 92 75 DD 27 52 8D CD 71 F1 5C 96 35 12 B9
 38 0C 84 7D 44 4E 10 E0 35 5B 3B 9B 57 13 F7 28
 85 3D AE C8 B2 E9 B0 2E DA 12 F8 38 F6 6A 07 98
 2E 44 A2 3C FE 6D 35 ED C5 16 29 28 48 F4 8E 5B
 60 7E 1B C2 79 B9 4D 9E 0C 1A 80 4E 2E 15 27 49
 55 5E 42 F9 57 85 3B E8 9A D1 E9 E9 57 87 1B DD
 21 6F 4C 08 A5 45 8B 3E 95 D7 DB E5 DC 14 3D 88
 10 79 5E A5 F2 29 42 FF 35 9B F6 86 9A 0C 26 6E
 7D 8E 5D 8E 70 05 75 AA FB EB 27 21 2A 99 CB C1
 AA C8 67 CE A9 59 08 3E A8 2B EB 71 C3 21 92 55
 96 91 65 B1 00 E0 F7 15 27 F3 2B 85 42 83 73 CA
 F5 E0 0D 1F AF 40 78 ED 2B 88 80 4B 97 AB 01 D5
 90 88 F3 D6 DF 55 A4 8E 2C 58 DD 5D B1 67 AB C1
 83 E0 C2 DF C0 32 52 97 36 BF 3E C0 72 05 D5 D0
 D9 E4 DF 15 75 9C 2E 8F F6 96 D2 0A E8 1A 49 55
 DF BA FA 7C 86 45 00 6C 14 5B 7A 71 0D 28 7B DF
 09 6C 18 46 7C EA F4 85 40 AB 2B 08 71 C1 A3 78
 C2 EE 76 9A 8F DE D7 0F 94 A0 33 A2 52 55 03 8D
 57 EA B9 20 79 92 2A A4 7A 67 B8 BA F9 5F 50 86
 22 27 29 FB 48 28 9C 16 4F 8D 45 7F B0 FE 8A EF
 0F E5 89 FD 8B 53 88 30 11 67 CE 3D F4 B4 87 3A
 C0 55 6E BD CF 29 C6 C1 AE 56 B1 47 D5 DB 2F 80
 4B 07 CC 28 2B 65 DC E9 9E CC 0C 3F 85 28 4F 87
 E3 F6 35 9A 31 74 5C BD 80 02 FA 58 77 BF 77 80
 8F 7D 97 CD C2 E3 DB 0D 1D FA 32 9D 7A E5 50 F1
 28 13 44 C7 62 48 D4 13 21 75 BB 91 A6 58 F7 CD
 AD 8D CC 3D B1 77 4A 66 41 0A EF 92 40 F5 96 00
 1F 05 A0 7C 5F 97 69 72 C5 43 E4 67 8C DE F0 8F
 4C E3 88 D0 DF A6 C5 B9 D2 81 CD 25 5A 31 4C A1
 F7 23 3E FA 85 2B 71 60 70 95 C0 4B FA A4 62 C4
 8E 71 63 D9 5F FE 80 B6 F3 B0 FB 68 66 57 BD B9
 B2 71 44 DD EB 99 86 7F 1B FC FB 23 F8 07 1E F2
 B5 82 04 13 25 77 17 16 FB CC 46 0E 1F AE FA C1
 A5 36 6C 56 6D 49 73 E7 43 C1 24 17 DA 4F 63 6A
 A3 E5 E7 6C 90 1B 35 94 9F E2 4A 19 C7 A4 7F 8F
 CE 68 A1 3E FE AA 3B D3 AA FD BD 67 07 24 18 10
 B0 74 4A 2E 58 0D 03 71 97 E7 EA 20 B1 66 1C 6F
 28 04 8C 86 37 E4 FB 94 E7 01 F8 BD B6 3B 39 D8
 FB B7 ED 29 C0 9E 11 1D FF 02 FB 5B 37 2D A3 6F
 81 08 47 57 5C 40 52 34 31 1B 2E D6 8F FF D2 1A
 B5 37 49 03 9B 8D 52 71 81 04 50 C4 3A 34 3A A3
 6A CF FF F2 5E 01 62 BC D3 F2 0F EA 13 20 0F CF
 6C 91 8B 12 DA 11 74 73 83 CA 64 7F 42 84 1A CF
 56 7E 9B D6 D9 28 D1 7B 80 80 32 D6 67 7B E8 1B
 2C 0C F5 ED 2B 46 0B E5 63 BD 2A 01 94 5C 67 5B
 3D 75 BE 02 92 EA 2D E8 1B 00 64 FA 8B E1 EA EA
 D3 29 36 66 25 D7 A8 57 0E 7E 8C 31 FE 9C 8B 43
 6E 0B A1 D2 5D 6C 60 A0 ED 2D 52 28 1D 25 DC 1A
 16 48 4B A3 30 E9 C7 3C F1 34 A3 2E 9F 6A 11 64
 74 E8 EF 62 B8 48 0F 90 A2 D2 4F F3 99 CD 0C C7
 92 EC 18 62 7A 85 6A CE 15 44 AE EC B4 EF 28 D9
 B6 F3 4C 03 57 73 D8 33 F8 BE 7A 1C CD F6 21 CD
 8D 46 1D 79 E4 5E 31 89 48 09 64 83 EA 05 C6 BA
 67 D1 33 13 9F 2F 78 0F D4 82 80 96 6E 2A EF 95
 CD AF DA 84 21 B8 73 D1 A1 31 F1 92 26 C8 A2 15
 06 5D C0 81 06 8A 9C E1 29 B4 84 21 21 56 70 99
 BC 82 10 E3 2A 43 E6 E9 E1 34 54 C9 61 8F E4 FE
 46 D0 10 C7 56 D6 BB 2D 3C 7E 12 48 0C E7 26 77
 45 72 D6 F0 85 F6 8B 76 ED DA 25 3C 1E F7 ED 3B
 4E A6 53 55 EB 0C B2 EF 59 2E 68 54 A3 B4 B5 07
 3D 26 20 19 B4 72 F0 D6 3A 4C F6 67 05 06 DF C8
 D4 34 23 08 3B 90 DB B1 1F A2 01 67 69 90 65 4D
 CC 47 5E D6 91 E9 E5 1B 86 63 7B 99 A7 1F C5 32
 8D 2B 99 E5 97 FA B4 4F 81 37 97 97 4D 4F 33 B9
 26 2A 03 2B 7D DE 30 81 94 E7 29 33 1A 6C D0 78
 5C 8D C7 9C 59 EE 28 0A 1B ED B1 1B B3 E9 50 A1
 B0 6B 95 DC BE E0 3D 54 2C 77 3F C0 89 78 76 39
 CD 6F CE DF 6D 2F 03 BC 03 79 AD 81 6C 9C 1C 7B
 5A 86 88 DC A1 57 F0 41 A4 8B 46 9C 60 C5 F4 27
 1E 50 B1 61 9A 25 7E 90 F0 17 68 C5 63 E6 86 31
 02 AA 8A 1E 11 A8 62 92 DA 15 3C F0 99 18 30 45
 4E 2A 0D 9A EE 52 E4 5D 23 4B 7C B7 00 36 4E 53
 EA 44 9D 22 3D 3A C5 22 C8 F2 54 F1 F5 E7 BE 61
 96 F3 6B 01 FC 6C 9B 94 73 4C 21 FF 92 BB 79 F5
 18 6B CA 0B 10 FB FD C5 65 E2 FA 2A 22 BD 6B 33
 D2 87 86 FB A6 CB 4D 6C 1A 39 DD 4D 65 F4 BF DE
 FE 67 FE E1 05 E1 EF 14 D3 61 8E CC 97 F4 45 E8
 74 06 7B 1A 15 56 0B 89 49 1A 42 FF 4E D9 D0 47
 3D CE 45 3B 85 ED B7 01 65 3E 98 85 17 CE 19 91
 FE 85 1D EF 33 CA DD 3B 96 2B BB 3B 24 14 E3 68
 2A 54 53 35 DE F9 4D B3 AE 48 08 6F 93 67 46 3C
 A3 17 B6 4E 47 19 F0 F1 CB 30 40 5D CC 38 1E C0
 7A 9C 4B 26 3B 2E 70 74 BC 51 85 D9 B4 00 52 59
 45 CD FF 3A 52 0D AD 78 BF 9F 98 8F 41 93 EE EE
 14 5A 99 03 57 DF 9C D8 1E E4 8E B4 E9 EE 54 44
 37 27 19 06 44 86 AB 28 AF D2 14 CC 6E 1B 90 1A
 1A 4C A5 21 82 D8 05 50 47 CD 69 90 FE 46 29 71
 71 57 F5 37 BD 9C 44 D6 CE A2 5C 6B 00 C0 60 AC
 3C 0B 0E B6 4D 32 9D 50 4B 1F 2B 07 1F 4F 18 EE
 89 A4 18 0B C9 CD F3 63 49 AE 8B 7C 70 45 80 18
 D9 8F 64 C0 DB 88 8B E8 ED 4E DB 54 1A 2E 23 99
 77 69 16 B3 01 69 98 8A EF DC 77 DB 39 95 56 A4
 91 34 6B 8A CF CB D7 FB 52 F7 D5 85 8B A9 E9 45
 6B 8E 55 0C F6 A4 2F E6 7A 7C F3 7B 02 1F 61 49
 F3 B2 94 0D 4F A4 62 78 2C DE C5 6E E2 53 AB E4
 7F 79 91 1A C6 06 E7 DC 73 33 C0 3F 71 81 5A 68
 C5 E4 4E 1E 2B C8 E6 FF 95 D6 01 A9 E1 90 3E F9
 37 5F 2C 93 60 1B FB 1F 1D 45 7C 20 7E 20 B9 77
 54 66 FE 08 13 04 10 24 9C EB 87 40 E0 FA 2D A8
 F0 E3 E7 F9 00 4D 1A C9 B7 60 BA 3E 99 50 50 B9
 F6 72 5A 46 55 FD F6 12 4B A8 56 04 DE 3B 6D C3
 15 88 0C 02 E2 B5 48 99 2E 3A C0 90 1C B0 1A 1F
 40 73 16 2A C2 8A D2 45 BC E4 12 5C 59 35 0F A4
 58 FB 24 E7 AD 18 10 64 E2 EB FE FB 7D BD 6E 3C
 A8 A3 93 75 04 69 37 95 24 72 AC F5 4F 16 6C 6B
 44 8E F6 CF 1D 83 CB 40 3F 89 1A 55 8D B6 9B B9
 CF C6 62 8F 45 5C 43 0B C7 00 DC 0D F8 D6 74 54
 0A FF BE 5F BE 92 F0 57 C8 38 D0 6E 0E 46 F2 34
 88 CB 17 12 72 70 A3 50 1B C5 81 EC 56 2D A7 EF
 77 B5 9D 63 62 EF CC 91 10 D2 11 B1 CD 1B 33 CB
 4B 5A D4 35 B6 1A 19 DC D0 16 94 37 B1 78 B7 BA
 0C 63 89 7C 2E C2 9B F9 79 07 86 1E 1F 7C AB 57
 C1 CA 22 51 CF 7E EE D5 67 BC D5 00 A2 D2 1D 9F
 DD 1B 38 53 D3 FB 63 C7 BC B0 E7 CE CF C5 FD 8B
 E3 DC 84 EC E2 B5 FA 84 4C C5 32 B7 6D 4F AE 76
 F0 18 4B BA 88 E8 14 B5 08 B0 17 3A 37 19 4F BF
 D1 03 0D CC 42 B2 94 33 04 DD E8 F6 DB C4 BE C0
 A2 8E DC 62 10 9B 93 F7 DD 95 E9 46 DE B5 30 1F
 FC A1 D4 4B BA C5 29 BE 64 B9 3F BB 7A 4B 23 A2
 00 B2 9A 70 E6 9F 2A 21 ED 32 01 45 96 27 04 E7
 B0 FC 5E 96 CB 06 28 AC DA AE FD 30 4C 15 84 11
 CB 09 15 69 6F 35 99 9E 9F 30 1B 7B 46 3F 5D 50
 F1 C6 74 92 72 31 D5 F8 AA 7F 89 81 7F 8A 84 D7
 E2 75 F7 EB 12 54 99 E0 87 6C 19 3C 56 FF 39 10
 0B 4D 4E D6 7E 8B EC BE A3 19 61 C9 32 F0 1E B1
 E4 8C 18 24 8C 93 C4 AC D4 39 BB F8 F8 9A 0D C9
 E0 4D ED 12 32 AB 5E 6C DC AB B9 E7 C9 01 4E 61
 07 8E D5 F9 5E 62 9D 5D 50 BB 93 C3 EC 6C 3E E6
 34 C9 B9 00 B6 8A 26 C4 3A 9B 54 F9 79 EA BF 97
 B3 B0 9B EF 91 AA 27 7E 72 32 4D 02 32 A2 E3 CE
 8D EB 25 C1 DC E8 89 83 6A AC 92 7A 70 C7 EC 72
 0C B1 74 B7 BF 0C 7A E1 46 80 1B 28 87 9E F7 3A
 E7 F8 03 71 A5 65 FA 90 5B 02 2A 2D 7C 8B 23 05
 85 37 88 C6 17 8E 23 95 52 08 0F F4 75 9C 9B C0
 CD D5 68 2C 1B 7D B8 4F 54 EB 74 A4 17 4C 0A EE
 43 02 C4 4B 4B 95 04 BA E9 59 C9 09 0E 50 78 9F
 91 39 0B C9 08 A7 58 CF 6C 6F 84 16 0F F9 69 32
 B4 18 C0 12 D2 A4 1E 18 89 D2 EC 69 28 BF 8D DD
 54 D8 58 7F 89 5C CA 27 4D 98 82 F8 2B AF 2C 71
 96 A5 C2 AD 52 08 65 FB EE 2B 0C E6 D7 01 83 3F
 B0 3A 0A F2 1B 93 30 75 5E FD 83 EF 21 60 E7 4E
 03 E7 BA E4 42 25 91 71 88 48 92 EE 21 DD CF 1C
 3F 55 E1 C4 F1 6D 16 DA BF 3F 8E 30 28 EA A0 95
 6D 66 69 24 41 2A 82 17 20 82 21 8D 13 2E 4C C5
 58 9B E7 90 BA 7A 46 E7 D0 55 C9 8B 95 19 40 A2
 1B 1B 9A D4 EB 0E 83 DF A3 D5 A3 94 6F C4 2E FD
 57 4D D0 00 58 B6 73 4B 3C C9 E4 43 B7 3F 8A 72
 22 5C D1 F4 EF 1D 95 3C 20 9D 7E 7A F5 2F 04 CC
 0C 8E 42 FF 42 71 6B 7D CA 9D 57 25 22 3A 8D C6
 2B 25 D1 94 40 81 93 4F EB 3D 59 35 74 A1 F3 EE
 F3 EC 69 E5 B7 FD 3D 5B 08 AB B6 FC 91 DD 0D 03
 76 55 5A D0 CE CC 82 B3 2D 13 E5 E2 D2 F4 FF 63
 A2 82 B2 F4 7D 1C AA F1 A9 D9 FC 44 E0 70 FE 25
 BC EE 4D 4D 6C CC 06 2A EF AF B3 F5 89 8F 08 22
 24 08 51 ED BA 58 C2 60 49 24 84 CB D4 D2 0F 4B
 25 5C 52 30 03 CA 71 0D 25 15 31 C8 B2 A4 DD C3
 E2 53 0C BB 20 AA 18 C7 60 17 0C BB 01 7C 81 11
 F5 84 8C AB C7 CA 85 8B 7C DB 35 D8 55 4A 49 E3
 F3 44 6D 44 F1 DF 64 4C E6 2A 9A 61 86 A2 69 1A
 29 49 66 AD 05 37 29 3A C0 0F B1 F2 97 5B 6D E6
 B5 25 5E 43 AA AE 10 20 33 6F CC BD 64 A5 1B 87
 83 D5 5D 3D A3 C0 8C E9 10 CC F3 1A C9 85 31 17
 7A 32 90 BA 37 72 42 6A 8A 61 BE 84 CE 60 DF 15
 A2 AB 93 17 29 EC 63 E7 DF 90 9B 3B 52 18 0E 33
 CD 90 DE 2A 7A 77 A1 BB AB AB DA 71 5B D4 6C 63
 52 84 E4 A5 91 7A B9 BD D7 20 D4 7B 7D 03 A0 66
 72 38 F3 8D E4 25 8F 43 4E 59 CE 01 44 33 8B 12
 EF 7E D1 94 23 08 DE 1F 67 3C F6 17 05 C6 F4 39
 B6 BD D5 59 A4 A4 8E 1D 68 87 76 B5 D2 6F 8F 5E
 3F 62 9B D8 B5 75 91 96 3D 17 50 D5 69 8A B6 EB
 44 15 1F AA A7 65 B3 EB A4 0B 15 50 10 9D 54 BA
 61 1C 6C 53 CF B1 A6 82 CE F6 D7 61 8E AF F7 A7
 B6 A6 62 C1 0D 72 43 E1 52 E0 39 09 FF 76 3F 3D
 42 96 4B 0E 45 6B 85 D9 62 52 AB 52 D3 C1 17 57
 84 AC F0 4A 0C 4A E1 47 F2 76 D8 12 EB 11 91 75
 D4 97 77 D1 EC 98 5E AA 2D 5D E3 00 EE 43 DE 7B
 29 73 92 4E D6 1F D0 88 E5 5A 9D 37 F8 A9 DC 26
 AE 3B 7A DB 5B BB D8 F8 4C E4 06 9D 51 5D D7 9E
 F6 95 EF A7 E8 93 D4 6A 3A 05 6F B8 AC 37 4B 88
 89 CC 27 60 BC 55 24 40 4F 8C B9 AC 41 38 D0 21
 00 3A 17 CE 45 0F 0F C0 35 0E 83 DF 59 D6 20 42
 68 1C 80 8C 37 36 EA 31 70 44 17 A2 90 63 D3 51
 13 8E D2 7D 7F 53 26 D7 F6 5A 21 70 A7 10 A4 95
 96 8B 6A 43 A1 35 33 6B 02 26 83 D3 38 15 8D 3B
 D9 56 EC 70 D5 B1 FC 16 E3 7A 4B C8 F2 31 85 B7
 BB CB 20 64 19 D0 14 33 1C B2 0E 21 1C 29 AD 27
 B2 A6 9F 0B 66 41 B6 59 79 D1 D0 6A A5 A9 DB E8
 9B F5 AA 88 CF E1 4F 57 B8 C1 7D C2 AD E7 2B 02
 14 FF 0A BB 51 B5 E4 7A 6D 90 21 56 D1 63 D0 4E
 B5 D7 12 36 EB DF 47 AB 61 57 D2 B0 25 0F EF D4
 6B 99 C1 7E 43 9A D1 00 92 61 91 CE 0F B3 38 57
 E6 15 48 9A 19 76 E7 26 F6 76 97 E3 CA 0A C7 E0
 89 AD B5 D5 97 22 73 77 FD AD CB 11 8E 35 5F FA
 2A A0 62 3F E2 75 59 36 64 0C 34 D9 7D A5 34 5F
 21 68 8C C5 48 15 84 2E 46 41 C8 E2 2E 62 D2 72
 E2 DF 31 F3 5B B6 C5 42 80 2F 8B EC 53 57 BF B4
 58 0C CB DF 47 FA 85 BE C2 50 08 AB A7 29 0D B9
 C7 59 4C 06 17 FD 0E 7F 02 A7 57 83 B3 B3 D4 CE
 0F DD 29 C0 9A 64 9B E1 9C 08 08 C0 C9 A0 1F 06
 52 6E BE 3D 3F 0C 23 5D CD B8 8B C8 76 0A B0 E6
 BF 89 8A E2 85 ED 49 63 FA 15 BD 51 2A 50 39 A5
 48 D0 67 A0 32 BA 12 CE 63 21 BA AD B6 9D 53 4C
 F4 26 79 02 22 C2 BC B6 5C EE 4F 0A 17 24 67 09
 1B 5B A2 F1 B3 C9 B1 71 E9 29 B6 35 26 E4 4C 1F
 AB A5 0B 97 42 3C 74 E8 FC 9C 24 B9 94 68 FC AF
 F1 4C 75 E8 78 7D 80 30 24 08 DD D6 81 9D 69 98
 B2 2F D1 71 B0 DC E2 BC 44 7E CA E7 EA EF 36 F6
 D2 D9 58 26 B3 5F 87 18 30 71 0E A3 38 8C F8 45
 8D FD 0D 15 35 49 4A 12 2B 50 8E EF DE FC 7F C3
 D5 32 4E DD 92 11 24 1E A6 31 A8 B7 83 22 11 D8
 91 C8 8A 86 B2 01 AC 0A AB 45 38 EC 7F 75 99 27
 E9 E2 97 C4 71 BC 9D 5C E8 27 E0 41 E2 13 FB 6F
 B4 36 0E 5A 4D 4F 75 89 05 FC A7 DD 25 E7 F0 33
 13 1C AF CB 66 80 E3 94 69 90 D7 27 F5 AD AF DA
 06 F1 C3 5F A0 54 88 1E 6C 5B 80 72 1B AC F5 CD
 BA 5D F8 8E 4A BF 23 51 A5 BA 6C 85 B0 82 9E 49
 97 51 A3 67 F1 2D C4 51 AE EB 64 A6 E3 ED EB 69
 1B 15 9F F8 16 B7 A4 9D 93 07 6E 18 B1 D0 22 84
 67 60 E7 CE 98 ED 7F 95 D9 A7 5C 38 E2 97 5C F1
 C1 3F 24 87 27 2F CE 05 08 E0 7C BC 39 0A A7 53
 8F 45 14 F5 AE 9C EA 84 B3 FF 54 BA 31 0C 6F 44
 FB 3A CB D1 73 76 E9 EC C9 34 55 0B CA FA 5A 17
 D2 D5 BF BA D0 FE 3A 5D 2C 0D 6D 31 A3 3B 0D A9
 B6 FD 9D 54 20 27 12 0B 15 ED A7 30 A5 09 A0 D1
 32 4C B4 01 50 14 1F 1B 94 1E 3C BF EC 36 EF 73
 22 1B E0 2E 38 F3 90 81 17 E5 BF EF 6E 13 05 7B
 26 5E DA 0E 1B 43 94 C0 8A 84 4B DE E6 35 30 E0
 19 41 67 53 3E 14 27 07 5D 5B F3 47 57 ED 72 BF
 51 AD A4 71 31 97 12 9B E4 29 71 1F 71 61 39 8B
 FA 86 01 46 7B 43 B5 8C A4 35 10 5E 25 6F A5 F7
 80 85 DE C4 40 B7 2C 65 D7 AF 93 C4 D7 6A DC 37
 A7 3B E5 A9 4B 8C F5 D2 06 8B BC 60 FE 6F 18 81
 D2 8A B1 D1 3E 13 3B 43 48 1B 85 4B E5 4B 24 D1
 66 91 FC F9 44 85 2B 4E E9 2D 35 F9 8D 36 7E 88
 1F 59 EC EC 60 B7 52 3E 03 75 E0 38 76 07 14 A0
 A7 E2 03 53 4F B3 28 FF CC 03 98 4A 5B 19 49 EC
 10 0B 38 E2 4F A0 48 04 13 70 4D 5F AC 78 D8 A8
 3B C2 D4 94 77 5B BC 26 82 0B AA 64 C3 2D B2 F9
 E7 41 5B A6 06 AA 5E 32 79 0C 97 D9 9B 89 78 B5
 48 15 B0 4B 2D B1 C7 0B 4D 7B 0B 3B 5F A5 4F 4E
 39 02 1C 3D 50 A5 A1 E5 BA 5C 9B 28 1C 38 61 17
 A0 94 A4 EF EA FC 4A BE BD 79 18 E9 2F 39 B1 4F
 4D 51 64 18 32 EC 6F EB 3C AC CA D7 DE 66 F9 05
 FF 53 18 B3 2A 39 07 DB 60 8E 74 8F 07 B7 48 90
 18 1E B6 64 DF A1 51 8D BB 3C E2 88 2F BF 01 62
 18 F2 EA 15 57 1C FD 5B 8F 42 F6 24 34 AA D6 1A
 B9 8F 9D 18 AB 45 C3 34 66 F6 89 F1 E7 B8 B1 2B
 5C 1E 7B 7E 55 68 0E 59 9B 10 64 E6 FE E3 B1 94
 FD 19 CE 18 96 62 24 01 60 CC 3F DB CA 6C 2A F9
 D0 D5 37 59 A6 84 88 D7 53 B6 8B 33 E5 62 80 F5
 A9 EC E2 95 65 D3 D4 D7 7E D2 B4 3D BD A7 02 03
 C9 50 87 D0 5D AB DB E1 38 21 DD DE 2F D1 33 24
 3B 12 22 AC 4E 6D 06 0E C0 DB D2 D6 AD ED DD CE
 0C D6 5E 6D 4A 84 8B 8D C7 DC F4 E1 E7 33 C1 A6
 9C 06 83 66 0F E2 32 67 CF 12 04 8A 41 D7 2C 43
 A3 B5 18 95 79 77 C3 8F 10 3A B0 24 8D 92 E9 EE
 7C 3C 24 5D 58 65 9C 7A C9 C2 BA 99 DD 21 3E 6D
 1E F1 63 EA DC D4 1A 7F 87 B9 71 AF 05 5C F8 24
 47 AD 89 5B 56 A7 69 84 E1 5C C2 96 FB E3 11 8E
 C4 B5 B0 F5 81 E2 32 FB 97 7B 9A 9A 1A 2D 59 72
 96 9C 97 DC A6 66 48 CE F9 08 1F 65 69 15 C5 8F
 81 68 B1 20 24 F5 D4 7C 33 11 17 7F 87 79 E6 84
 BB EC 94 E8 4B 91 EB 69 A0 EA 0F 4A B4 FF 3C 99
 96 3B F1 E1 BD C1 F2 7D 1A 98 24 4A 0F BD 90 A5
 04 A3 4C DF EB C1 D9 5C 83 DB B9 11 18 25 FA 09
 23 CA A8 B1 3A 1B 33 19 B9 6F BB 8F B5 79 68 8F
 6C 4F 5D 34 2C 49 78 55 9C ED 82 F4 11 C0 D1 32
 CE 2B 93 FA 16 3B FF 65 F3 1C 0E 5B 5C 2E 0E 2C
 31 88 3C 03 5E 42 25 03 45 41 DA 12 E2 95 1E 76
 BF EB CD 09 7C BA FD A3 48 4A 2F 8A 3B 95 5B 41
 F0 7E CF 8F 05 B3 B9 45 52 74 75 73 DE C6 C5 45
 6B CE 57 CB 89 22 65 EA 3D 95 BB 77 09 FF EA 67
 59 45 87 84 A5 7C 71 F8 9B 12 89 4E 7A D4 3A 70
 B4 8B 2E 07 06 FE B6 B0 30 8B 48 A7 23 55 5F DB
 FC BE 56 45 F5 62 A0 3D D8 AF E2 E8 E8 47 DB 91
 AC A7 8D 99 E0 2E D5 2B 9A 53 31 CA 63 65 AD 9B
 99 86 F7 49 12 2C 7F 56 23 E1 B9 7E F3 C8 0D EA
 26 08 DF 2E 50 C6 E4 26 4D CC DD EF 9A 73 F7 35
 D8 8A B4 F9 24 CB C9 4E 62 C5 14 8C FE 77 71 4B
 C9 16 6F 43 4D 4A 8F 6C 29 BD 84 E5 46 90 F5 63
 42 1E 34 B6 CE CB 49 B2 AF 87 39 41 00 5A 6E 07
 FC 3E 44 AF D7 38 9A E5 8A A0 F0 34 7B F0 6A 2A
 BC F0 27 30 23 F0 82 62 F8 13 3E E4 BA 52 81 73
 4D D5 69 91 BC 62 2E 52 F7 4B E9 02 7F E4 A6 84
 12 FD 52 1A BC A4 DB 2E BD AE 64 D6 E8 75 07 D7
 ED 5D B3 3E 52 EB 78 9B 8B 32 3B D5 D2 D2 82 F1
 89 BB E6 2D 00 12 EA AD F1 AA 8A 5B 2F 18 8D 28
 5E 31 C8 E4 A5 B8 FA 38 9C F7 09 26 58 C3 36 4D
 D7 90 98 63 16 AD A7 62 DC B0 CA 28 40 32 7B 50
 34 FE 69 CA 6C DE 37 54 EC 9A 13 57 76 FF 89 62
 F6 39 02 C2 B0 EE 3B 7A B7 8C A7 C1 CA 4C B9 58
 27 04 ED 99 03 35 51 2D 2B 64 34 73 6E 39 62 AA
 8E 43 1B 58 C1 25 46 6A FC 0B 06 B8 71 33 2B 92
 C7 BA 18 40 86 7D E2 33 5A 17 75 72 D8 84 E5 80
 58 92 71 63 00 FE D4 93 90 70 E2 BE B3 51 45 27
 5D AB 5B 34 DC 9E DE 92 8C 07 C1 E4 8F D8 42 43
 33 D9 F7 21 1B BC 1E 95 F9 E9 3D A2 57 5F 50 B0
 1F F9 57 93 0D 41 91 0B 80 88 A3 F9 D5 13 52 B9
 36 4F 48 DE 6B 8A C9 A6 A2 51 07 9F D7 28 C1 B7
 03 CF A0 86 38 B2 C7 A5 08 DD EB 0A BD BC 0F E1
 E5 A0 51 06 46 F7 6C 67 29 BB 7C 61 0D 63 E4 ED
 45 22 EA 3E 9D 34 30 00 CA 0A 3A B0 EE 11 A7 F1
 C0 AB 95 C9 53 BD 61 4C D6 28 CA D7 F7 38 DF 7E
 48 BC B6 70 4E 82 F0 31 5C E6 DC 9A 9E A0 F3 9B
 1F DA DA 6D 4D 25 21 48 5F 1D 0E 5E A7 DA 06 20
 79 A7 2C 19 03 F0 40 DA 58 1D 16 1D CE 83 FD 29
 B5 78 9C DC 29 2B D4 B5 C7 41 67 25 15 AC F5 CC
 A8 4D B7 AE F0 DD 3A D5 1A 36 66 CE 8E 6A 9E 1E
 71 A8 D1 39 06 89 24 60 CF 7F 93 8E 43 36 98 95
 92 6A 05 C7 F6 D5 6E 78 8C 57 74 5C 4B CE 47 AE
 92 95 B4 6D A0 F0 E7 94 C9 18 59 B5 A2 8B 47 BE
 DF CD 9D 3B 1F F3 77 7B 99 C5 29 DD E0 38 F8 88
 6B 09 B2 FF 6A 4B 06 94 E8 2C A4 1C DF BA 88 5C
 7C 20 71 2D 13 D2 45 75 4C 47 72 25 83 84 EC 73
 D8 4C 95 5D 55 25 9D 0E 79 7F 47 E8 C9 E0 20 AC
 0D D6 2D 7B D1 0A FD 71 84 EB 3B F2 DD 3F 83 F2
 D3 92 86 A1 85 0A 75 FA 03 EA CF 0D BB 46 E2 CA
 09 30 AF D3 CB 85 2A 8C 75 75 87 03 8A B4 CB 2C
 A0 02 6B 25 53 19 1C 2C 2E 47 DF 74 BF 0B 25 06
 BC 81 CF 0F 54 F7 9F D7 87 C1 7F 3F DD 9E 45 D8
 D2 AE 8D 78 10 FB 87 C5 53 72 25 95 E9 AA 38 5C
 48 2A 95 BE D2 E9 84 B6 28 CF 16 8C F2 54 1C 4A
 83 BF FB 9A D5 DB 77 18 23 C1 2D 0C 01 2B 0F B5
 7F 03 BF D7 EE 0E EF 58 81 B5 69 48 95 60 97 EE
 9C 86 9A 17 FE D2 58 21 31 A3 EC DE 62 3D C1 3C
 1B 9F CB D7 2F BD 26 F7 C8 02 F7 A5 F4 51 FC 09
 C7 05 F1 E2 98 97 5B C4 87 3D 49 2D 97 9D 40 95
 AE 02 B1 33 0E FF 40 2C 6C F8 7B E2 90 ED E3 DF
 CE D3 DF D3 F9 AE CB 48 29 BA FE 98 F0 50 3F E6
 8A DF 14 6B 35 CD D8 C9 4B 39 55 1D D4 13 95 B6
 6B D5 4E C9 CA F5 F7 A5 7D C0 38 82 12 25 E9 61
 B8 DE 15 F7 CD 12 D4 7C 0C 08 B2 C9 49 97 19 97
 43 7C E7 1E 32 81 74 27 DB 57 8E 18 20 7C 4D 74
 25 46 89 AC 10 3B 74 FD 95 40 76 E7 61 0B 45 E3
 47 98 BE 05 28 37 A0 4E 73 50 85 6D D5 D6 25 E9
 1D 1C A8 71 69 09 5A EE 9F 5B 9D BE CD 08 25 87
 86 7E DC E6 86 02 E1 C6 05 65 9C AF 98 E0 65 D1
 17 57 11 62 6D FB DB 8A 1B 86 4E 85 5C B3 C0 67
 CB AF D0 5B 7F CE 9C 68 9C DD 48 52 0E AD 6B C6
 AB 67 08 6A 87 CA D9 E8 08 F5 32 16 AB 08 EC 0C
 66 6D FC 58 A0 25 D8 78 8B E8 D8 A6 DC D3 25 99
 A7 FA AC 22 B8 BB 9B 9E E3 40 88 FE B7 75 B8 E9
 E9 5A 64 80 19 E4 2B 62 A8 08 E9 2A 89 81 39 2C
 0D 86 E1 5B 6F A8 47 0C 26 78 E3 E5 37 C7 86 72
 66 84 F1 B5 E5 14 4B 7F F8 4E 5F B6 A7 98 18 50
 88 78 7F 7D AD 83 15 E6 09 40 3C 57 07 08 FB 8C
 8C 98 B2 19 CC 53 30 D3 D0 EA E8 8D 65 44 D5 4D
 B3 EC 00 BE 0A 4B 4A D7 77 F2 65 65 45 E8 AE 1C
 75 81 38 4C 83 B2 53 9C FC E5 9D 37 AA 15 6A C8
 E2 06 29 23 A6 DC D0 EA 15 BE B1 F1 3A 66 AE B7
 84 71 17 BA 89 68 25 C9 F1 86 B8 64 99 CE 57 05
 42 DA 50 7F BC D6 DD F5 55 8A CA 84 2E 88 91 49
 E5 5D FB 57 74 61 48 EE E0 F8 06 67 33 BF 8C F1
 F6 EF 0F 77 B0 57 F0 0D 97 42 A8 47 68 BD 12 B7
 92 76 DC F9 8E DE C0 2F 66 71 59 FB 6C 2F 22 46
 A7 13 B4 75 4E 05 16 DF 55 AD 17 31 A7 AF C6 E4
 5B E8 12 84 BF 52 A0 15 ED CC E9 4A 26 19 57 53
 B2 56 71 AF 4E 70 68 3A 16 00 FD 3F 55 2C D4 F1
 9E F0 3F 6E 3E A0 F8 E4 88 0F 3B 5E BF FF 2B 11
 D3 FB C9 DE F5 E7 3A 8A 98 FB C4 CD 70 4B ED 86
 F0 E9 4A 42 B5 F3 C7 05 84 69 EF 02 09 B7 53 DB
 0B F3 C5 07 8D AD 93 17 99 86 34 04 A5 DF A1 55
 AC AE 33 48 1E 20 57 CC B8 C6 C8 98 68 3C D1 E9
 50 75 87 92 6E E6 DC 41 EE 90 B0 9B D6 09 7A BB
 B8 2B B0 C8 F2 11 BF 16 37 2C 69 7D 34 94 8E 5B
 B7 97 9B 77 83 9C 39 45 A1 81 A5 AB F0 EA AB 45
 B6 C7 62 0C 10 18 C6 47 07 2F 42 1A AA 54 1A CD
 5D 2A 61 6B 37 23 A6 EE 28 87 8A C9 78 E2 60 4B
 4B 20 A7 EC 3E CE 4D B5 EB 7C AA 87 97 A2 40 FF
 08 15 9F 4D 8C 09 0A 9C 36 AB BC B7 B1 22 40 00
 BC 98 7F 62 97 B2 3E B3 E6 31 16 13 72 92 FD C7
 B2 73 49 42 8B 56 A5 1B 71 77 EA 77 8E 08 D4 4C
 C4 F5 6B 80 A4 8D D3 33 EF 64 85 61 B2 6A BE 69
 13 8B 79 EE 8A 23 ED 39 50 2C D6 62 E2 63 70 AD
 F4 ED E3 01 5D B0 64 C6 E5 3F 33 99 07 22 19 83
 45 2B C9 C4 96 84 82 44 DA 62 A8 3F 34 C5 3F 6A
 F4 9B B5 BB A1 5B F2 1A 35 EE F5 74 1A D9 E2 27
 75 7C 67 B9 5A 36 86 12 00 FD 80 C9 DD 95 15 6E
 B2 CC B1 11 68 36 B2 4F BC C6 36 8C 0A 58 64 5E
 B7 97 B4 EA FA 2F 81 3C 52 9C 32 EA 14 55 23 94
 4F C7 2A 5B 74 99 55 AC 7B 19 06 6B 5B 09 BF CD
 0C 28 79 06 28 90 25 DA D4 85 42 F1 8E 1C B3 E3
 15 48 92 CD 7F 93 37 85 8C B6 94 BE 3E F9 B4 8B
 B4 EB 12 24 43 46 C5 40 9C 78 37 33 90 F0 44 74
 FF 98 11 08 37 4E 15 EE B3 E0 BA 9B 9E 8B 64 F3
 A8 A3 D8 67 A9 27 FF 39 7A C7 C3 8C B9 65 18 A6
 6D 2B 2E 6E C3 BD 55 0A 48 0D 37 9F 42 68 CF 9B
 03 1C 0B 96 FD BF 90 82 1C D6 7C 4E F5 D0 AD 25
 65 AF 5F D2 BD 4B EE 64 EE 87 2A C5 A1 2F 52 EF
 E1 23 F9 E1 5C 96 3B 48 3B E6 D3 59 A2 F6 E8 72
 A6 E3 03 2B 5C C5 E0 33 84 6E D4 6A A8 1F DB 5B
 A5 ED 6B 2A 22 01 AC 64 31 32 8B 1F 38 37 C5 C3
 FE 6C 1D D3 9C 21 CE 27 FE A3 F9 78 06 A3 67 1E
 C3 7F 4E B4 83 A4 CC 71 AA 38 8B 3E C5 91 C0 CA
 99 D4 28 AF 02 CE E9 C8 41 A7 6E 37 AC AA 68 59
 08 5A C5 6D 6E 9A 81 5B 93 C9 11 3C CB 65 1F C7
 15 B5 B9 6F 56 DB BD 0C 2B 1C 07 7F D8 E8 3C 9F
 51 B7 70 5D 00 02 54 FE 3A 10 EC 9A A0 92 30 E3
 F2 92 79 55 84 29 56 E3 8C A6 55 B1 D2 12 EB 24
 45 68 2A 41 01 7D B7 7C 88 93 43 0D 9C EE F3 1D
 38 A1 09 AE 6C A0 D4 2C 8E 3C 63 FD 9D A4 A6 F9
 BA FE 0F 4A 6A 19 DB 8A 71 7D DC 66 67 2D 18 37
 93 A6 D5 20 74 B8 03 F9 87 94 79 4D 98 B0 67 D0
 17 04 4A 68 04 52 CF 2F 12 CC 8C 58 D3 04 73 0B
 97 19 0A D3 22 F6 99 21 D5 FD 29 EA 31 C5 B5 20
 31 D7 6E F4 89 03 28 23 82 95 47 40 74 90 56 61
 20 03 D9 80 60 3E 99 E2 64 73 64 83 4C C7 2A 7E
 CA 92 9E 90 3D 7C 50 81 EB 15 91 6D 2F 0B 76 3F
 78 EF 76 96 F6 14 27 4C 44 29 FA 5A ED 8C A5 B5
 21 09 57 22 C9 27 F3 02 83 CC 08 B1 06 15 96 00
 3F 07 39 3E 4F 8D A0 7E 62 08 F8 49 3E DD 4C C0
 86 5D D8 0D FA 07 D2 19 1F 37 F4 4E 76 26 63 B8
 58 CD 13 FD 96 C0 C4 DB A6 E1 D9 D8 F5 6A 07 D1
 9A 74 FD 33 84 95 6B BC B8 5D EB 74 6F 34 81 B3
 E7 D7 4C D7 3D 39 54 7E 96 22 C6 C6 54 0B 5A 58
 E4 91 DC 3E D0 C2 EC F4 FF E1 56 F8 66 C0 6E A6
 04 2C EC 5A C0 88 54 FD B3 DD AD 14 31 93 EE 15
 52 BC 70 26 74 49 D7 1C 6F FB B0 74 0C 8E 69 9E
 FF 3D 3B F6 BF 25 65 81 7C 1D 0A 4B B9 9C A8 24
 E8 F3 A3 78 DA 87 B9 B2 33 95 82 30 B7 03 BA 71
 8C 80 20 F8 5A 30 86 D9 1B EE F5 01 E1 60 6B 8F
 B5 3C 1E 52 09 0C 6E 86 45 E8 C2 A4 30 49 71 02
 4B 9F 12 31 AA BF 93 00 F8 5F BF ED F6 E8 4A AB
 70 C9 4B 30 2F D5 E8 4A 41 B0 E5 A1 37 06 B9 EB
 0A 40 D7 4F 95 53 CF 72 1B A4 45 A5 3A 46 0E AE
 F1 22 AA 9E A5 F4 29 AB E1 01 EB AA 58 AC AC C3
 58 51 10 6C B9 A2 D9 15 C8 13 DA D7 93 BD 07 F0
 56 75 F9 1D 5D 96 95 B8 95 F5 F1 36 A1 3D 23 78
 4E 73 22 F8 72 FD 56 84 AC 64 6F 88 4E 51 40 9C
 A0 8C 9D A7 05 68 47 16 3C F9 3B 20 0E CA 08 BB
 52 45 0C F2 F1 BE C4 0E 73 CB 2F 71 78 58 1E 47
 8C D5 08 DB 34 3B 0C 0B D3 CD 04 95 94 2D 25 54
 40 32 B9 E6 D3 9A 46 75 CB C0 5A 63 A6 E0 1F FD
 F0 40 1A B6 1D 61 29 12 F1 FB 2C 0F 44 B0 76 DC
 F4 55 1E 06 54 F9 E2 17 AC 89 3C 7D 7C 8C 55 ED
 7E 19 EE 6D AB 42 2E EB BF 8A 9B D5 3A 1F 00 76
 CA 0E 5B E0 F7 73 00 56 16 0F DA 61 E0 DD C8 6B
 73 CE 74 9B 96 18 0C F1 3D 00 3E 8C FC CC 5E E8
 8E A4 45 5F 70 5E CD 21 DB 10 30 EE 82 1B A8 21
 8C A9 55 85 59 D4 C4 80 F6 82 1D BE 2F 34 DB 88
 C4 80 1C D4 F2 FA 5F 03 4B DE B2 7A EC 13 61 95
 39 2E C9 DC 28 B1 8F 9A 66 42 4F 9E 9C 63 F3 24
 94 F9 80 1C 5D BA 6B C6 0E 51 EA FE 19 4F D0 7C
 29 33 4A 60 BB 8E 20 A8 F8 0D 85 7B 99 D2 F2 EE
 7B 18 F7 FE F7 1B 14 F3 86 8B C7 5E 46 73 44 FE
 F1 00 12 86 21 28 C7 BE 7A D4 4C 89 B3 91 DB 36
 66 F3 D1 B3 16 4E A9 B0 0F 8E B2 E7 F3 E3 C4 D8
 2F 3F 38 A3 DA 15 14 F6 7D DB BD F8 DE C3 65 88
 DB F7 13 E7 05 B9 53 DC 36 56 2D 0E F4 BC 62 3A
 D4 61 AD 3C CD 43 2F 05 33 BD E5 44 C0 9B C2 CD
 24 14 98 B4 A7 20 90 71 04 42 E6 47 EF B3 C0 69
 14 CA 82 08 78 CD C7 10 C1 E0 2E D3 71 2D 5A 0E
 D5 FB 1C 24 B1 FB 98 61 22 AC C1 CF 26 8A E6 A0
 EE A1 26 C3 71 E4 D8 C5 AB 9A 6D 1B 96 31 F6 DB
 35 F0 D5 3A DA 38 78 A2 A6 FC 3E D9 29 E1 5F B8
 F4 92 E3 5E 01 39 8E 91 1E A3 1B 65 6E D7 DE 4F
 9B 94 F7 52 FF C5 A0 D7 95 CF 50 D8 8C 47 EF D9
 E5 F2 4A 04 8B 09 2F A9 A2 01 55 0B 85 BC 6C 3B
 DD 8F D3 E1 5F D2 4E 2D 08 30 09 AC 21 AB F8 9A
 4D 7C 93 4C F9 FA 28 2E 55 C5 39 11 34 72 32 0A
 90 BE 15 36 3F D5 05 3D 90 8C 6F 58 A1 B7 C2 FF
 11 65 69 0F 6E 68 B4 AE B9 DD BD 16 AC BD 88 C9
 F8 F6 B9 BF 3F F7 0E 38 58 BB BD F8 C7 67 E6 01
 BA D5 21 C0 1E F8 4D F7 87 50 27 B9 47 D6 02 A5
 86 ED 97 2B 1A 8F D4 EF 15 82 48 84 C3 88 B0 CA
 99 1D 6E DE B3 F2 86 B5 69 7B 96 A2 7D 99 F1 15
 DC DF 52 68 B6 60 D1 7A 0F 9D 33 C4 8B F2 63 A7
 CD BD F0 E1 3A F7 D2 FA 28 BA 7C B9 76 63 47 7E
 16 7A 71 84 0B 46 18 15 B1 98 69 91 96 CF 34 1F
 47 89 EA 33 3B 27 B5 5D 0E 62 46 C3 BA 4C C4 DA
 79 F2 3D B7 18 B3 91 1F EE 23 97 27 9D 06 CC 78
 CA BD 42 BE 76 49 AA 0B 51 78 2D 73 64 D9 EA 86
 E8 A2 88 AC D8 04 70 14 2F BA 91 4A DC F3 FE E5
 27 9C 5F 7C 0B AC 33 72 6C 20 C2 D4 36 83 F2 FD
 31 D4 C3 0F 4D 4F B4 84 30 13 3B 23 A9 A6 C6 2C
 69 DB 95 CB E7 82 02 D8 73 68 2C F5 50 FD 75 33
 7C FC 5E DC 0C F0 5C 27 0C DB 1A 2A 6F 7E 4C F3
 9C D1 7E 28 3E 25 EB E7 DC 2B 5C 9F 76 56 E6 0A
 E1 16 26 22 C9 FD FE 27 AC 91 1A 03 36 2A F6 43
 4B E1 63 46 85 32 82 63 CE 13 6C AE 89 CC 1D 2D
 04 35 C0 9E 34 3B 1B 61 93 89 8E 34 8F FF BE 93
 EA AF 89 F3 04 16 90 63 39 0A E3 03 86 47 BD 04
 64 12 B2 F7 F9 F1 EB 23 A1 C5 B6 4D 61 35 75 54
 23 6B 58 D7 64 81 E9 F2 67 D9 1B BF 0E 53 B4 CA
 7D AE 10 14 87 FD 8D 10 E4 47 8B 7D 9E 22 71 FB
 0E 24 31 1E CA B8 83 A1 80 44 16 1F F3 F6 7D 14
 B9 4B 67 32 D7 49 A6 13 57 A7 00 F0 73 3C E7 F7
 27 33 19 04 4C 3C 5B 7C D4 38 93 28 DB ED 87 2B
 3C 82 41 C4 F1 17 B7 34 C3 B6 0B 74 8A 42 45 C8
 55 73 81 F5 60 37 26 9F 62 26 52 61 80 7D 71 D6
 69 FD 57 DF 56 64 4C 4F 37 9C D1 FA 6A 5D 7C CC
 08 DA D7 3E 50 53 EE 2B 78 5C 8B A2 75 7A AA B2
 B8 8E 9C 04 BF 49 98 2B CB C1 06 67 4B 54 EA 42
 A3 7F 97 5E 8A F6 6D FE 6F 91 9B 4C B7 C4 17 FA
 41 22 71 80 73 C7 29 D1 9D 77 AC 10 9D E4 4A ED
 56 13 3F 5A 26 41 F9 B2 AC BB 0B 95 AC 3A 3A 4D
 DA 28 B9 C2 7B 92 9D 58 A4 D0 97 DD 6F EC 3D C8
 36 06 F6 F9 81 0D 53 C4 53 0F 5B A4 1F 2A AA 3E
 65 06 39 08 C3 10 0D 4D 3E 7F FC 48 F0 07 54 6E
 A4 A6 A2 CD E1 F1 42 23 2A 81 FF 43 AD F4 A5 19
 32 AB 41 C6 26 3F 73 AB A4 29 4E 0F 9F 30 D0 9E
 F4 93 B4 58 C1 E7 DC CE 80 78 E5 B7 4E 1C 7C 41
 DE AE FE 4A F0 0E 57 C3 43 C7 95 00 0B 0E 51 1F
 92 56 E7 0C 71 01 D2 AD 30 0C 67 6C FC 4E 93 FC
 F0 E2 ED 7F 99 E0 F2 3E E4 3E C8 96 04 80 3D 3E
 D6 0A 10 83 47 26 2D C8 65 72 C0 2E E1 3D 39 EB
 DA 68 34 C7 22 89 2D 21 81 1B 55 5B 8B 38 CD 16
 20 97 22 12 5C 1C 93 92 B0 1A 6C CB 66 7C 58 34
 7F 08 3F B8 E1 AF 35 5C 24 5C 87 01 35 04 14 AB
 3D A7 4D D7 92 42 92 AF A0 68 2D 56 70 98 3C BC
 EC 92 D4 4E AC E7 F8 AE CD 08 85 0B 9D 29 4D EA
 28 06 E0 0E 46 ED 91 BA DE 4C 85 40 5E F9 F4 30
 A5 3C EC 54 C6 2A 68 DC C4 4D B6 2A 99 1B E6 DA
 C6 0B C6 DD BD 93 A2 77 E1 66 E9 8D C5 A0 F4 97
 00 F3 E4 0C 8B 49 57 3E 8F D9 23 A9 16 D9 0E 92
 01 3E DA 2A 26 0C AA 7F 6A C3 74 D3 BF 61 58 A5
 D1 0D 08 59 81 17 36 00 91 C1 CC 61 35 0D B0 E2
 A4 63 12 E4 A9 00 E5 24 B8 72 94 7B 4D CD 07 07
 B7 DA 88 4C 50 67 D3 C6 50 05 6B CE C3 BD A5 41
 34 71 26 35 EB 9C 84 BD 7A 49 57 DD AF C8 58 4E
 6E 54 B3 ED 2A 50 AB 60 24 A0 03 87 18 DC 13 F4
 AC BB 5C 3B 5F D7 99 A2 D7 B7 A2 96 FB B7 E2 40
 8E 5A 26 64 5D 6A 3A 0C 11 26 2E BB AA BE 74 D4
 BB EC B9 6E 6D E3 AF 1D 31 1D 1D 46 B1 EA EA 4B
 25 5F 0E DF 0D 33 EE 1D 08 05 D1 E5 B3 2D 81 EB
 15 BA 45 BA B1 A9 E4 A4 B0 99 73 21 A2 0C D1 34
 12 48 7E 95 20 0F 56 AF ED 11 82 28 D3 A7 73 EE
 2D AF 7E 51 ED AF 5F C4 23 B6 83 EB 32 1F 38 F7
 E1 F0 C3 B6 CA 70 E6 47 14 E6 DD E8 A5 CE E7 03
 C0 68 0A 90 05 50 85 BC 4C 30 86 C9 D9 52 55 F5
 F8 FB 09 EB 5F 8C 07 AB 7A 3B 85 E6 79 AE B8 27
 21 9E 90 B7 52 43 EA 21 7A 8D 3F E2 CA 09 7F AF
 74 41 98 72 C2 33 A6 8E 61 B3 6A AE 53 FB 56 D3
 84 0D E0 40 FB 8B 59 B6 06 26 E5 B5 39 ED 55 33
 6C CD C5 46 EB 1B 35 CC 3D 38 1A 8C 73 DB AF 49
 1F 97 25 BC 1E AB A0 9B 9B ED B8 55 E4 4C 4F 6F
 02 85 12 8E BA 24 B0 3C 00 DE 50 23 0D C6 F7 A7
 2E 23 D1 35 FB BE C7 24 F3 65 E9 C3 95 4D 49 88
 05 9C 2E 87 A2 C9 6C 1E 68 70 08 F2 6D 4B E0 B6
 87 B1 95 5A 37 30 EB D0 C3 26 C7 48 0D 0D 2C C2
 6F 38 17 2F 9C D3 DD AB 1E 29 4D C0 8B 7B 72 F1
 ED C8 EB D1 B3 59 83 EA B8 41 DC 24 E7 68 12 07
 31 18 A9 31 B7 A4 54 1E CD 6E 06 3D 42 6A 68 FE
 54 2D 69 2F 8C 87 46 6D D9 5C 56 DC 9A A1 8C 96
 C3 85 A9 B3 F5 B0 9F D3 90 85 88 2F 3A 29 EA 91
 22 DA 2B 95 E9 C8 92 55 53 66 80 22 F0 7E 26 30
 9E 7F 02 E8 03 B9 D5 F0 86 98 80 7B 0D 2D 92 DF
 2A D5 9A 36 AC B4 BC AB 8A 67 26 BD AA A1 2D EA
 BC 04 81 35 28 E5 1D B1 A3 E3 6C 81 61 33 01 87
 5E 88 3E 6B 1A 1C 4E 52 17 DC 53 5F 1E 54 24 8E
 C1 6A E8 A9 06 C5 81 29 BC AA 9C 61 6B 8B D3 97
 67 D5 75 4D DC 41 2D 52 C8 A2 54 AB D4 B4 8A 19
 6A 69 94 22 11 A2 F0 34 6C 91 F5 3E 6C 9F D0 A8
 26 E0 27 34 23 6A F8 29 7A 12 D5 80 2A 4E A0 76
 C7 3F 0D F9 EF 24 B1 71 24 04 A7 E3 E0 C6 AE 02
 17 77 FB 8B 21 B8 78 B8 5C 05 B6 98 05 19 DC 28
 3D FD B3 91 FF 43 26 A1 10 B4 D4 37 25 64 FD B1
 D8 F3 63 D9 2C 1E ED DA EA F8 A8 FF 88 9B 7B 30
 1A EC FE EE 01 DC 5E 74 68 5E E2 9B 30 C6 B1 BB
 BD 40 C1 30 CF C8 1E 14 58 AC 9E 81 C3 C8 A2 83
 76 55 87 20 C5 48 35 A6 BA 7C 45 FE A3 38 DF B5
 FA 15 E0 5F 62 F7 78 2E F4 ED 48 9B B0 83 D4 2C
 83 85 6F 52 65 3E 19 95 38 48 6C C8 66 6D 57 FB
 DC C2 94 5C 86 12 EF A8 A7 E8 24 26 59 AE 12 BB
 25 42 BE A1 56 97 16 6C 11 D0 F3 74 15 78 99 D5
 1B B1 B8 AE 73 6C E5 20 28 E3 01 47 73 20 5E 46
 D8 21 A0 03 A6 95 87 00 E2 1F A3 B4 C3 A3 8A 53
 43 FE 21 30 EA C2 EB 2C 40 C7 7F BE 8A BD 07 A5
 19 47 78 73 07 1B 27 47 1E EF B4 00 86 B3 DE 24
 7C 2C 5B 30 A7 46 7A 29 65 1B 00 B3 DA 42 3F 9E
 04 9C 83 39 FB 68 08 FF B5 C7 F4 FA FD 5B 22 D5
 5E 9F 8F BE EE DA 71 E2 E3 C6 DA AA 6B 53 A6 67
 94 45 F9 02 09 74 8F C3 C5 31 11 68 5F 5D 3D 5C
 C6 0C C6 F2 9C 81 B4 F3 DE 62 36 FA 6A B7 9E E7
 BC 45 DC E0 D7 BC B6 CA 51 76 49 23 BF 67 1D 15
 AA 50 B0 33 0E FE DF EE FB 37 A3 82 1F B3 5E 70
 B2 DC CF 3F 12 30 46 64 DD 04 D7 D4 F2 A0 FD DD
 E8 39 6C 28 14 71 7E B2 12 C2 0B B8 13 56 4D 1F
 FF F6 05 BB AB 51 03 2D 63 3B 16 54 C4 BA BD 09
 95 21 4B 9F 79 5B F2 B0 96 72 79 03 F1 E0 48 B1
 6B BF CC 20 70 73 94 FB EE E7 C6 9C E3 FE D3 52
 7D B4 A3 1B BD 0D C9 E6 96 CB C9 E0 FF 27 01 32
 98 41 CD 76 12 F1 5F BB 9B BC 44 26 84 C0 68 E4
 A4 EA 77 0F FA 5F EC 77 25 BD 83 34 6B EC 71 7C
 A2 7E B6 8B 44 5B 53 88 87 DE 8A B4 B8 D6 D5 C4
 35 DB DE DD 4D E7 91 11 69 F8 75 73 BB B5 FF 79
 95 BF 27 F5 40 A8 07 4E F4 8F 14 CE 99 FE 2A 78
 CC BC 3A 74 E1 18 66 C4 D3 48 19 5C 60 F2 2A 0A
 D8 05 CE 85 7C DD 71 B6 11 D9 EF 7A D9 32 9C 61
 B7 48 BC 32 39 FA DE 6D 89 E1 C5 D7 E8 4A 2D 8C
 5C 04 DF 7D EB F6 90 08 DF 7F B4 F5 71 03 F9 CD
 18 C4 43 56 15 BE 42 A9 2F DA 7E 4D 24 C8 7F C9
 24 83 91 6B E8 94 C4 96 54 8A 1E FE C7 8C 54 46
 AB B7 9D F9 DC 77 2D 72 2E 10 3E D6 4B 62 0F 68
 A7 76 B7 E3 A5 01 43 9B 06 03 8D 9D E9 2D 44 A3
 F9 0F 69 DB 1C BA 6D E7 F1 F8 E2 5B 8B 6D 4F D8
 C3 41 C7 F3 87 6D 22 DB 39 80 27 2E 5E EA 4B 52
 92 B4 A2 E3 DE 42 51 06 5C DC FA 98 E2 91 C1 4A
 3B B7 A9 A0 7D 0A 1F 59 BD 4D C2 3D C0 08 E1 EE
 09 E6 2B 1D 86 4E 43 7A EB B7 F9 AC 1F D5 D1 D1
 27 95 22 3A C5 E6 35 CA AE 30 32 E4 A1 30 EC BA
 78 AB B6 99 04 36 CE 4D 9E 4A B4 46 F7 63 7E 5E
 D3 EC 86 24 CE 8E D6 70 3E BC AF F5 BA D1 8C 2E
 C1 4C 19 D2 AD 5E 01 0B 20 DB C9 95 C4 1B 43 A3
 A1 0A 55 E3 C9 7D EF D7 9C BA E3 5E 86 FD 93 B3
 F2 8A 4E A7 FD F8 25 9F 10 A7 4F 94 E4 22 12 4A
 6D 39 01 AF 9B E0 D9 07 06 A1 59 45 03 3B 61 FA
 21 54 30 E4 D3 FE 1F 78 86 C0 A3 EC D0 EF 9F 75
 4A CD 5C EC DD C3 75 6B 76 3C DB CB C0 90 8E DD
 8C F5 C5 E4 25 33 74 CC 65 3F 8F 0A FC 85 4A 9A
 BE 35 DD 38 D5 29 77 F1 07 BD A0 F1 D8 AF B3 57
 43 1E 22 19 99 82 6C A6 98 37 DB DE 32 56 FF C1
 02 5F B7 A7 9C 05 8B 1E F7 51 0C 7B 1E F3 99 34
 18 65 4F 61 AE 00 5A AD 8C 12 8B FD 13 01 5B 3B
 9F C3 55 AE 1A 4E E9 51 BF B1 CD 10 FA 10 68 EF
 B5 01 7E 47 EB A7 60 B7 6C 3B FE 18 F6 5F B9 04
 9F AC F3 5D 6D 3A 3D E0 D9 EE A1 98 4C 8C 32 C0
 0F 12 CB 6F 7E A1 FD BB 7E AF 3D EA F2 5C 70 59
 E6 E2 1D 19 8B A0 7E 30 AD 8D 2D 78 E9 FC 15 69
 99 F9 93 5A 75 CF 25 7F 11 46 1B 32 59 08 A1 41
 FB B8 DF 69 75 B2 39 E5 68 AE BD 4D C5 9D A8 EE
 D5 02 EB 06 5F 71 FC 0F FB 3C 14 FC F6 92 27 F0
 C6 46 25 71 C4 4B 20 16 87 D2 B2 7C 82 28 39 3A
 A6 C1 A8 4E FF 0C FF 3B 76 D0 37 44 F3 0C C0 89
 62 0F BA 31 F6 2B 40 8D 7C 28 2F C2 13 FB 86 2D
 6A 93 D0 D8 20 BE 4E 79 7C 5A 52 74 11 8E A3 61
 1E CB E4 5E C0 F3 52 94 F4 57 2D CE AB 53 66 A8
 7C 8E 71 2A 02 81 0E 80 6A 79 51 11 81 57 4A 86
 CF B6 4D B7 88 F1 4A 2A C0 32 64 5C F3 FA 12 3D
 26 02 39 B6 40 14 36 13 24 92 52 15 E4 A1 7B 9C
 54 BD 74 89 13 3E D1 14 CC 0D EC 9F 82 B2 F3 56
 E1 9E A8 99 BE AD 33 6C 19 A9 54 AE 38 93 B6 5D
 FB D5 F9 D4 ED 00 AE 9D E2 E7 F1 8B 7F 34 15 57
 7E 7A DD 37 7C 50 C8 89 52 CC 69 EA A9 2D 3B 73
 5C FD 89 47 3E 17 95 D3 9D 9D 7A B5 A9 AA B0 5A
 8B 98 B0 2B A9 9B 08 87 3F 19 2C F8 08 C1 3A B2
 B4 CA BF 41 85 5C 28 F4 CB 77 5C 4F 50 F5 8D 12
 A2 C9 D4 E4 05 4E 86 AA 86 85 3C 6E F5 78 EB 3D
 25 40 B9 04 5E 8E D6 9B 62 30 0D C8 C3 0D B9 46
 A3 CF 59 49 33 F2 B0 3C 60 26 5F C4 1A 9D 1F 10
 F0 00 F8 D5 DC 78 B5 A9 BC 82 59 B6 A9 73 4B CA
 33 51 4B DC 79 33 FB 2A ED AE AC 05 4B D7 B9 EB
 10 0C 3E 77 7E 10 07 46 AA 75 4C 87 95 B0 12 14
 4E 94 C5 AB E7 19 56 D9 64 18 30 32 3A F7 64 42
 1E 22 7E 47 7B 30 B7 B0 B8 B2 4B 01 7F 15 84 47
 69 8A 84 29 94 33 1C B9 57 75 9B C2 50 74 3A A3
 D4 9F 1D 5D E9 94 B7 58 A7 8F DB 85 A7 69 C5 91
 BA 69 08 3B FB 63 E3 9D 34 39 4E B3 82 2D 45 0E
 E5 9F 7B 96 4C 23 7A 7D 86 E9 DB 89 5C 80 A3 7E
 3C FD 39 F2 37 AF 1E 5F 7A 36 DC B8 56 FE 51 F8
 D2 AF A8 1F 76 62 1B 64 38 F9 E1 3D 53 DE B6 38
 7D 9E 10 8A C3 7A BF 46 05 F6 DD 9C 8E BA 5E 81
 C6 17 9E 3A 5A 12 E3 E2 DA A3 B4 30 6E 15 6C F8
 B8 6A BE C8 7F 73 65 9C 9E 9F 9D B5 6C DF 7D C3
 71 4E BE E2 79 B8 6E 56 4E 6C 17 7C 4E D7 87 DF
 AE F1 A5 AD EC 70 81 A5 E5 57 2B CE 9D 0A 42 C5
 F7 4A A7 28 1B C0 71 4B 7E 67 2B CC 1D 14 2D 40
 68 5B B9 7A 25 EE 74 3A 49 5E 14 A0 F3 3D 94 6E
 2A C4 E1 CF 91 24 9F 07 8E 81 8E 13 D9 2B 78 CC
 66 A5 67 27 70 08 2B 32 AA A5 BB 01 03 7E 09 5C
 13 13 22 6C BD CD 05 1C 00 6A A8 36 A9 09 13 F8
 6C C9 95 15 35 12 AE 18 9C 94 64 C1 F9 5F 00 6C
 00 AE 63 7E DC 23 CF E3 1D B1 C3 CC 9E DE E6 94
 FA 1B 37 2C 66 73 C2 2C 85 48 9F 45 09 29 06 28
 2D E2 F4 04 3A 47 1A EC 33 EC 70 9F 95 2A 17 94
 1C 2D A3 F6 87 7B B4 94 DF 88 49 F3 52 73 40 BC
 BD FE 72 79 0B 13 2B 4F 9C 2D EB 6A E3 8B AA 4D
 D0 7F C2 E7 0C 49 17 A5 46 4B 50 CE 65 37 DE 0F
 01 6C F3 78 9F 45 83 EE 54 C2 62 FE 5B 77 6E 5B
 A3 48 B1 F1 30 31 D7 88 BB 3D 92 83 E5 B2 D4 1B
 CB 64 38 09 CA 47 CC AA 42 D4 D5 65 94 F4 FF B7
 C0 5D 9E 0F 6C E1 F5 A3 A4 B8 0C F9 64 41 6D 55
 0E 99 57 17 6B 14 79 13 7A 54 99 DA 36 A8 18 64
 D5 4E 1B 39 BC 7F B2 ED A3 E7 5B C3 01 4E 1D 21
 5A DC 6A 2D E6 4C FF BB CA 57 D9 D1 D1 52 0B 3E
 5D 5D A3 9A 1D 96 E6 0F 39 C5 79 08 38 BC 59 00
 07 E5 33 23 E8 E7 CA A1 5C EF A7 2F D0 EF 5F AD
 06 BB F1 C1 20 73 72 60 C5 BA CF F3 46 07 09 63
 80 03 06 96 57 61 96 91 4F 02 13 79 F9 4E EE C9
 87 AD 59 F6 61 52 06 FE 34 54 9E B1 05 CA 72 7D
 C3 BC 08 B6 C7 99 36 E2 82 5D CC E7 08 27 C4 F8
 1E 59 4F 09 33 DA 7D 58 57 D9 1C 36 34 CE C0 8D
 02 1F EF E1 1E B0 43 3C 33 17 A6 B1 3B 0B 74 A1
 D1 B7 AF 29 96 B0 38 01 BA B5 4B 9A 12 9A 55 02
 B0 26 5C 3D EA 64 0C E0 D0 C9 3C 68 86 A2 7E 30
 D3 12 54 6D FE AF EB 10 32 30 D6 57 BD 9E 16 B2
 E5 52 65 68 16 A8 0D E9 76 5D 5C ED B4 29 B8 73
 28 7F 00 7D 1F 72 73 8C 5A 28 82 A0 4E 40 05 D6
 49 AA 54 98 26 42 C9 B6 C0 10 DC 87 EC 23 89 18
 8F E3 15 6D 35 F1 F3 1D B4 96 E9 87 A1 60 C5 E9
 53 11 BC 72 F5 06 70 09 0E CD A1 10 A3 BE 02 1D
 EF 0F B0 30 06 45 E6 01 DC E1 9D 7C CF B2 52 1F
 96 15 5C 97 7D 00 CE 9E 1F 36 6A DE BC AD 56 9F
 BA 2B 94 95 98 81 D9 21 7F FF BB A0 CD 9D 6E 1C
 56 11 D7 69 78 C6 BA 2A 46 28 76 8D C5 41 78 A5
 10 8E 09 9E 50 D4 2B 4C 64 18 E4 43 75 1B FF 49
 E1 65 64 09 52 98 D5 28 07 79 38 13 63 9D 99 9A
 09 EF AC 7B A1 3A 84 07 D5 F2 5A E1 26 81 11 72
 8E CE 6C 03 53 44 5A 16 D8 CF 25 A3 6F 37 35 89
 A0 36 72 74 C0 0A 46 E6 B3 1C 5A 75 2E 4C C7 26
 8A 6E A8 F4 83 18 B0 54 DB 19 40 5B BD 36 8F 6C
 C2 E4 B8 DE 1F 0A F6 DD ED A6 E9 35 A5 1B AE 11
 92 23 E9 7B E5 A2 75 AB 9C 37 E6 DF 02 21 82 9B
 70 29 01 05 A4 7D 91 FB 0B 54 CE F8 CD F0 53 6A
 2D 8E B2 37 78 26 ED 57 1E F3 8B ED EF 22 BD E0
 1E 55 9D C3 7A BF 03 E9 07 EB F4 A4 F7 5D 9E 7D
 01 53 DD 13 71 85 03 99 6F BE 10 E9 74 FC 06 9F
 6B C7 B0 08 33 42 D8 1A 50 A9 C1 BD 81 B6 4D 3D
 7D F3 26 39 B1 21 EB 77 18 71 42 33 33 4D AA 62
 B2 73 53 8D FD F0 51 1F 96 2A 52 18 BE 91 DF 99
 20 E8 BE 4E 54 6D FF A7 5D 2F CD C0 18 ED F2 D3
 D1 59 F3 C3 A0 8E 6C 25 79 C6 86 2F E3 78 30 8D
 D9 84 70 99 27 80 28 27 A5 AD 9E 0B D6 AA 29 F5
 E5 5A C9 69 2B 4D 2E 76 29 68 BA 00 5B E0 A5 7F
 BB BC F6 7D 29 E0 B6 A9 5E 1E B4 2A 7F 81 9B D1
 7B C2 64 2D CB 75 62 B8 91 B4 A9 E1 B3 60 1D 6E
 BF 74 61 B6 1B A2 1F 1F CB 44 68 C0 4C 1E FD 44
 93 D9 D8 44 C0 10 48 BF A7 A3 C9 6C 01 88 C7 1F
 08 09 8A 8E 25 75 5F ED 06 C0 61 F6 5A 46 D9 8C
 14 6C C9 D9 C3 B2 DB 03 CA D8 6B 0C ED FD 64 06
 05 39 44 82 2C 5C 45 C8 83 89 B7 0A BF 91 F3 7C
 1E 28 9B 42 35 DD 33 7B 42 78 99 CD 81 0F 54 08
 3D 74 07 AB 5E EA F5 0B FF 83 51 17 7F 2E 31 86
 33 80 76 51 E7 CA A9 6F FD 70 BF 20 08 DD E6 B6
 99 C2 D8 85 C0 5C B9 B1 8D 69 4E 91 42 79 29 C5
 33 EB C1 EA 47 E9 9B 19 BE 54 F6 51 57 38 2D CF
 CA EE BC C3 8B 7F B8 50 BE 26 BF 76 DE 65 10 99
 B4 31 F9 CF C4 E7 76 A2 25 5A 6F F8 68 28 80 2B
 0B 1C DE 14 1B A6 F9 EB 92 1F 12 D0 C5 D6 31 05
 11 41 BE 94 A5 D7 34 C1 02 EF 07 94 AF AF 68 7C
 4B 10 81 33 D6 4D 60 69 13 C5 89 B3 A8 F5 DD 9B
 2D 11 DB 54 56 8F 60 21 D7 62 57 34 DF A8 27 16
 A1 AA 01 F2 24 A1 86 74 71 E7 24 73 5A 85 F6 3E
 A2 6D F3 5A DA FB 07 A1 5B 5C E6 FA 6B F8 00 E8
 E8 25 E3 8E DD 4D 47 5E A4 61 BD 75 EE 65 A7 E4
 AA 40 FC 6E 8A 48 75 7F D2 C5 17 C8 61 CA 34 3A
 C5 ED 9A 0F D7 02 5A D6 77 5D FB 4A BB 97 81 C8
 8C 42 67 DF DF 8C B9 3E 55 7F 19 08 A7 58 19 17
 99 7A A7 7F 0F 67 93 51 00 79 63 6D 63 94 0B D2
 92 62 64 D0 3B 09 6B 9D 26 D7 9B 18 7F 17 CD 22
 BA 05 98 B2 35 C8 35 C9 D2 FB 6A 97 60 A9 C6 AB
 94 D1 D2 DE 56 15 B6 16 0F 02 E1 A4 EE 10 55 94
 42 73 EF 7C 37 4D 34 28 09 11 DE CE EE 56 F5 45
 9A 33 8C 0A A8 17 A3 2F 2A 7C 1D 1A 8D A3 A6 1F
 C8 31 86 41 69 3E CC D8 A9 DA 8F C1 50 83 5A EC
 21 48 5C 2F FC AC 68 54 8C FA 7E 1F F1 B3 8B 04
 59 50 D8 E6 69 D3 84 6C C3 B9 00 C8 5C 07 A4 87
 1F ED 35 B7 56 E7 05 70 17 F5 01 F2 4E FB B2 48
 5C B8 15 06 85 7A 0A E5 83 39 30 76 9D 7D 3B 28
 47 53 49 A5 2B 84 A9 F7 3D 62 53 09 CF D8 D0 CB
 74 36 28 B2 E6 B6 32 C3 AF A5 A2 4C A3 34 28 65
 B4 D5 D9 1D 4B F5 E5 EA B4 9D 08 FC BB 25 E9 F9
 9D 3A 60 7E A8 F9 7F 25 C6 26 3E A9 4E 9B 7C 61
 5A A3 B7 A7 2C 58 B5 1F 86 D1 DE 43 F1 79 C9 C9
 1B 7F 19 9B B8 5D 21 B7 96 DF 89 1C 87 11 FE 0A
 DC 15 50 D3 75 24 91 27 BC 27 C4 EB C7 8E 07 D9
 D6 E1 CF BA F2 55 9A CA 10 05 CF DD CB 4D 3E 20
 F6 7F AE 55 A4 31 C8 F1 A7 5F E1 9E 29 3C 75 82
 5F 4D C0 4B DD 8A 8D 14 C4 27 9C 35 A7 0D 3F 93
 5B F2 57 BF D9 6C D4 85 7D 4B 44 DE DB B2 C3 FD
 72 54 A8 87 27 EA 87 0E 13 1B 5E 6E 13 26 73 62
 AD C2 E7 52 CF D6 B0 02 57 0C 93 FB 7D 64 E1 AD
 45 E4 E9 4D 29 96 79 D7 A1 EE 74 AA 3B 3D D7 A3
 A1 B4 15 A7 C1 17 B4 83 7B 72 89 F4 05 3B 38 45
 33 4B 2D 58 85 B4 D1 99 9F F7 5C AD A6 9C 60 26
 26 1F 72 38 74 90 B7 6F E0 62 6D 19 B9 87 B6 4E
 45 D0 12 8D E6 00 AF 98 1A EA 74 F6 F0 8D 60 BE
 D0 75 3C D8 29 EB DF 7A 15 C1 5B 50 49 99 67 AB
 3F 52 A4 79 79 D2 3B 05 75 E2 C1 9E D4 6B 6E D1
 38 CF D7 C6 CE C3 1D A8 1F CF 12 86 53 49 B8 DA
 8A 87 6A 6C D6 09 C1 74 54 39 B5 1F 83 D8 3D A1
 1A 54 5D F7 BF 14 A2 A8 89 05 90 06 92 1D 7F D4
 DF 76 D5 A7 06 6F A7 7C BF 9A 26 47 4E D7 30 E5
 4C 31 6E F9 7D 83 67 AA FE 84 F5 8E 9D 43 7D 84
 F9 B7 8A 3E 12 58 0E 45 24 3D 0F DF 81 D9 E0 5D
 E1 89 B8 B0 52 37 1E 40 E4 6E 70 2E 70 A5 74 99
 FD DD EF D8 C1 E4 03 4A D5 BE E5 5C 4B 9F 33 08
 F1 6B 69 1E 2A F5 FA 17 2A 94 9E 6B 88 A7 ED CE
 1F 11 61 2B D8 9E 82 2C D9 03 E1 B9 25 02 26 81
 7F 32 3C 87 49 7C FC F1 F3 DF 9F 42 17 06 16 EA
 BD 04 82 19 8F 69 0A 34 BA 92 80 35 10 E8 B4 BD
 C4 9A 61 77 A1 9D 58 09 D4 AF 5C E6 12 2F EB EB
 65 E8 82 51 8F 25 40 49 0D 92 D9 66 F5 94 F0 0B
 55 DA 42 EF 84 46 1E 44 F4 AD 97 D3 A9 03 47 D6
 35 90 D2 D2 48 93 73 69 1D D4 0B E4 DD D8 DC 40
 F9 CE 09 E7 4F 4B 86 1F B5 19 EA 14 6A D3 00 95
 B6 38 96 38 4E D7 B3 F7 D7 99 13 4C 9F 0E 89 03
 58 D8 8C 2C 80 59 D9 5F 00 0C D4 9A 9F 74 6E D0
 45 55 BE 91 B9 CB 67 5A EE 22 28 83 9A 14 24 B7
 15 DD 9A 94 BB E4 7E 2D E7 F3 3C 81 1A 16 08 8B
 1F 10 62 46 7A 16 C5 1F EA BC DE A3 B5 2D 15 4F
 73 A1 72 76 01 0C B3 42 5F F8 96 77 12 F4 8B 3A
 30 F8 32 F1 CF 75 AA 1F 8F AC 15 7B 63 71 1E F7
 E8 C4 CB FA 78 17 B1 17 BC FF C4 EC 9F 13 33 B1
 FC D6 9B 03 7E FB 72 85 9F 3B 28 7D 07 3E 2C F3
 82 D7 04 3D 84 91 62 DC 54 50 66 AB 56 BC 0B F9
 4B 33 0A D6 7F 3A C0 FA F7 9E E8 CA AE 7F 20 52
 E5 E1 6D B4 21 EA 3F B1 AA 95 48 48 BA 25 D8 EC
 29 CF 23 AB B3 74 62 39 8E C9 9D 08 A6 84 FC 61
 79 BE 9F 66 CF 88 B4 F4 FD 47 AC 06 C1 86 85 90
 A4 A7 49 D1 77 0E 52 C6 5D 5A 7B F0 4A 65 91 80
 8E C7 3C CD 28 B3 65 6E A1 F3 24 8B 94 FA C1 EC
 F0 D2 E1 F4 E8 08 99 41 F8 A5 A1 72 5D 63 E3 14
 8C 6E 0F FC 70 BA C7 C3 AA 4C 96 26 F2 4E A8 65
 FE 94 29 6F 55 D0 49 00 77 E2 42 32 E8 18 42 6E
 31 CA EC DA 4B F6 D2 7F 49 F0 D2 87 66 D6 B8 D6
 CD 33 86 62 69 A9 A9 A0 EF 3C EA 90 25 84 0B 30
 0A 67 D0 34 70 C6 54 89 D9 1E 35 70 1B 86 9F 46
 79 76 83 48 10 E2 FC 38 EE 19 7E C6 79 C5 47 EF
 F6 10 A5 1F 49 3A 4A 45 37 37 90 5D 98 97 04 C6
 0A 41 59 C8 62 7E B6 67 01 4E 39 F1 AC F5 21 E6
 9E 5E 14 FB BC FF 77 78 28 41 85 ED 40 82 23 3D
 67 33 C5 10 2B 9D CD 6B BB B4 E7 6B 6C CC 79 04
 4C 14 D6 5D AE 03 FD B7 3F 24 1C 2B E3 25 BB 9D
 FC 1D 5A 8C 67 FB 4E FC 19 92 22 EA 3F 83 FD EC
 C8 F4 77 C2 74 40 96 1D 0B 71 0F 04 14 3B 84 93
 01 6A 55 B8 CC 44 99 7B 6D 48 06 B0 74 80 EA 2A
 30 2C 02 6F 8F 6F BC DA 9F 8C 9F 78 04 FF CF 62
 99 5A CF 43 E1 64 86 34 27 7C 29 92 58 47 45 F4
 31 A0 6D EC E1 A1 B9 49 D8 18 3C 13 46 E4 95 57
 D9 EA D5 38 CF 36 2A 1A 3F 9A 8E 29 5A 0B DD 24
 E9 E0 E8 75 EF F8 00 E3 1E 3C C2 F7 7F 47 95 D4
 6B 9E 14 96 C7 6B BF 22 6F FE 6C 0F 1C 7A 33 B3
 29 12 22 F9 24 D2 6C 46 1E 60 9C A9 EE 52 52 76
 38 1C 5A 25 E9 57 B3 98 50 A9 63 81 45 40 5C EB
 25 33 C9 34 A7 05 90 39 A9 22 D2 6B A7 39 00 04
 8D 2C 27 6C 68 7F D0 79 FF EB 5D CE BD 45 A1 47
 EF DC 2D 17 B0 1E F0 95 1B B3 89 33 24 53 B2 FA
 9C 28 48 7C 13 F9 06 45 1C D3 CD 84 C5 1A 25 3B
 D0 C8 2C E2 81 34 73 C7 7C 2F F3 BF 2B 37 DE E5
 72 73 EE C1 1B EC 6F 92 D0 FC A1 5A E4 D8 02 1F
 09 5E F1 DB 8B E5 99 48 80 B4 DF CF 85 63 05 74
 9A 64 25 78 DB 0C 65 3B 0B 4B 53 E7 9B 82 38 58
 05 93 9B 4D 06 78 BC 4A 9D F8 41 C5 22 EA F1 23
 32 5F 38 6E 5F 98 16 57 68 CF 53 56 B9 B9 1D 58
 53 22 10 9E 1C 16 3E C4 10 69 DE 91 DB 48 3F C7
 E3 73 B0 5A C0 1A C5 D2 37 D0 6F 71 E8 98 C3 C1
 C8 D2 92 CC 23 D5 1E 69 25 D2 03 AE B8 7C 29 A5
 95 D2 9B 64 0B 39 85 D1 E0 41 88 AC 62 67 32 D8
 61 7D AA 98 3C C4 08 62 D2 2B 42 28 51 6B A4 46
 0F C3 77 DA 1B 33 62 3A 7E B1 AA CF 81 1C 33 2B
 E8 30 70 B4 95 A4 5B 5A 3E C4 11 7D 10 02 9E A3
 7E 37 92 45 CC FA 41 E8 FD 4A EA BD F5 57 74 F0
 78 2C 93 84 6E 1C 55 FB 68 90 A4 6A 59 AE 23 D3
 8A FB 64 A8 CA C6 E9 3B A6 0B 91 A5 FB D7 74 B5
 BE D0 91 A1 89 94 76 8B 3D 2C 42 B0 79 D1 4F 8D
 10 9C BB 30 07 8F 5C EA 9B C2 FC 57 F2 65 17 67
 EE 55 FC E4 AF 86 51 3A 43 77 A0 22 BE 03 55 7D
 B7 FE E5 F1 69 52 43 96 33 59 E3 F6 11 4D 38 51
 39 09 8E 90 02 54 31 E6 47 91 12 00 D8 D1 C3 49
 42 BC BA 9E FF 8E 74 76 9E 46 60 95 72 36 BB 07
 BC 6C EC 19 3E AE 00 D2 19 BD 7A 76 81 50 D4 BC
 30 E1 A4 70 BE E5 C8 74 AF 61 83 B9 5A 24 74 CE
 63 C5 34 38 2C 03 E6 6D 76 31 2F D6 B1 D5 23 CB
 E7 48 3B B8 FA EB 0B BB F0 DA 65 F5 EE 8D 2D 81
 F0 1D 44 6D 3E FC 7F 18 3F 3C 04 14 7B 8D 17 71
 DC 6B ED 5D ED 20 96 49 5A CC E6 C9 2F 07 46 DA
 8C E5 66 3E 79 58 5D D0 C4 E7 50 8F AE 34 3D 7B
 D5 39 6A 23 BF 05 C5 87 82 84 3B 01 ED F0 97 3C
 66 71 9C 87 A7 83 0E E3 05 D1 2E CD 5B 69 13 41
 72 FB A6 3E FF 70 A7 19 AF 20 36 36 71 32 0F D7
 65 4A 58 D9 07 2B 23 5D 2D 1F 3D 93 2F 9F C1 B5
 EE BF 34 A7 A6 E4 6F 9A A1 42 FA 72 B7 3D 0A 99
 1A A5 56 F6 54 F8 D2 C3 D6 89 48 AF FD FB DB A9
 3B DB 25 25 BF 2D 17 72 14 4C FC 34 E3 48 DE 83
 29 26 2D 74 17 2A BA E2 B9 E8 FC EE C8 90 B9 68
 9C 40 21 F1 5C 23 67 8B D6 E2 35 88 AC 92 5C D9
 98 AC BD DA E4 16 F6 79 55 6F 77 4E 20 0E EF E9
 09 42 C0 5D 0D 6D 3F B8 9B B4 A0 98 18 DC D7 52
 37 23 34 FD E5 2F 43 09 B1 56 6B 92 65 97 30 16
 A1 44 03 87 1B 4C 21 54 27 E2 86 93 0C 7B F4 A1
 8D D0 AB 01 16 A2 75 32 C6 9E C4 3C 52 CB FA C1
 C7 32 EC 22 4B AD B1 4A 8C 02 5C 39 48 68 37 08
 0D 18 58 E1 15 DE 3E 3F 44 D7 A9 BE 96 DE AF 6E
 4A 6C 13 5A B4 98 0F DC 0A B1 F7 43 63 6D 18 F3
 FF 98 9E 6A 76 CD C4 C1 FC 92 45 37 F9 BB 49 CC
 4C B5 0A BC CC EF AB 0B 6C 27 FD 32 7B FE 8D 74
 94 50 C0 60 2E 59 29 41 65 18 29 4F A0 0B 93 44
 4D F8 6B 68 67 96 9C 40 AA 3E 33 20 97 92 15 2C
 5C 14 E5 24 D7 4C 01 02 91 88 7C FA A8 B9 84 2E
 D2 BD 2B C1 A9 2B AF 8D 03 30 16 1D CA E1 BB FA
 B8 00 9F F1 3F EB 0A D8 1D 4B 40 9B 24 30 F9 56
 3E 0E C9 87 0D 5F CC 20 5F AB 95 44 0D C4 63 14
 8A E2 69 8E 94 86 DF D0 1C 16 6D 18 A7 F0 B9 48
 B6 5A E2 9B 65 AC 35 44 0C 92 F3 98 7C BF 63 DC
 BF 6E DB 15 61 FF 88 67 A6 34 3D B6 7E B6 8E 10
 C9 3C 94 3F D7 2C 01 B6 DC E9 26 13 11 E6 FD DA
 8E 09 C8 24 98 BB D5 72 CE BD 70 D1 2B 1B 49 4D
 94 28 C7 B8 70 DB 06 7E 5F 5D F9 8F DF 06 62 64
 9A E2 A2 09 27 CF 1C CC 0B 61 C0 5B 62 7A BF 93
 D1 A8 27 03 1D 7D 9F 44 34 7F 69 45 ED 4E 33 41
 0C 10 CB 0D 68 E0 4F 2D D3 01 70 91 8B C5 08 35
 0F 17 AA 05 B3 FC 04 8E 87 4B AF 28 E5 80 AC 98
 D2 11 4B C6 4D 09 ED D2 E2 AE B9 8D 4F AB D7 2F
 AB 67 A4 44 71 9F 96 2C EE 1F 34 83 84 FA 48 CE
 68 12 E0 34 A8 EC 5C AE 5F 34 29 EB 63 F6 F2 78
 9B 84 5F 6A B0 58 0A 6C BE 3E 05 2A 1A 15 8A 6B
 67 F5 C5 43 EB 57 08 C1 E7 40 4C AF 0E 48 B2 B7
 CC 11 5F E8 83 82 9D AC 75 53 48 87 FC BC C9 DA
 94 24 17 24 2A 9C F1 66 DE E0 D4 31 EC D8 33 C2
 01 9E FB 0B 83 8F C9 BB 36 BD 2B 76 8C DE C5 77
 11 B0 94 92 02 AF 7A EC 75 10 6F D9 45 71 A8 B5
 DE F9 29 60 CB 6E C1 15 26 88 B6 33 07 64 74 0C
 7C 2F 90 AD DF 2B 41 21 11 D2 88 E6 31 DE 60 95
 F3 19 BF 40 43 9C 04 E6 79 72 34 F1 58 42 6B 51
 04 AB 82 B9 D7 93 A6 74 DF 0A 94 41 2A 73 FE 86
 8E 34 64 E4 25 3A A8 B8 38 E0 C8 9B 8B FE 8B F9
 EB 5B BC E3 7B 35 47 95 21 10 F5 D2 FD 46 72 AD
 98 21 6D C2 D1 B9 02 97 B8 7F A4 F7 E3 E3 A7 1F
 66 64 B7 54 B8 B2 66 C6 D1 6F 64 41 C1 D4 62 18
 67 BB D6 3F EE D0 B5 38 E7 62 FD F5 7D 70 55 E6
 9D 02 76 81 83 39 9C D5 AC 00 33 BF 17 07 F8 19
 18 85 E4 5D 25 4F AF 7F EE 74 A5 77 3F 3A EB BC
 67 02 49 69 A1 D1 68 7D 46 69 72 5C 50 7F D5 B8
 A3 F2 59 37 7D BF 02 BC 1E 4D 5B 3E 2F ED E3 14
 61 4F E4 15 20 E1 30 D3 06 30 C2 A7 A1 C1 3C AD
 B7 93 65 E9 D0 F1 B1 7A A3 B7 30 1D 05 07 7C 79
 A7 04 BF 13 55 9E 7A 38 2D B2 4F 29 41 45 29 58
 6D C9 FA 16 AE A4 E9 A3 DF E3 D7 39 5D 5B 84 EC
 3C 74 19 FB 9A 07 47 0E 4F 25 25 3B 84 A0 9D 49
 81 3C 6C A8 0C B0 AE BE 64 90 A8 99 4C 68 0B E0
 70 B4 D0 F2 8D 26 F9 26 6E BD 53 61 61 AF F4 BC
 8B 06 2B D2 5C 44 CF E3 7B 35 C3 7E 29 94 F0 50
 29 5A 14 90 2E 8B F8 00 C1 D1 00 61 24 F2 B8 75
 31 61 E1 EF 0F 46 C0 C8 11 C7 2A AF 6F 79 C0 2A
 AE 20 57 5F C5 4F 8B 72 C1 11 DB 9F 16 82 D6 07
 76 3D E0 66 4D 52 B5 11 2A 83 22 0E 9F 9E 79 F2
 47 06 86 D1 85 C5 5D C0 C7 4E C5 CD 36 73 19 62
 CE E9 33 61 C2 0F 2E 06 F8 70 EA B5 37 A3 B8 5E
 99 8E 8E 14 E4 7C F7 B6 61 34 26 D0 0E 40 35 52
 B6 E7 FB E8 CA BB BE 63 37 55 0A 28 8E DC B7 6A
 86 D6 C9 AA 2F E8 81 58 11 91 71 E1 CD 24 07 EE
 ED 11 0E E6 45 7C D6 6F 1A EF C0 AF 5A 3C 76 E9
 0B BF C7 8F FA B2 EE E9 E0 59 20 C2 71 5E D7 46
 70 39 0D 77 55 1C 51 FD 27 E6 39 4A 4F C8 30 27
 F1 02 3F 37 33 E9 0D CF AC 41 BA 1D 23 1A BB 2F
 76 04 B1 B1 E9 E3 1A 9A EE 7C BB DD 98 CE 5F 4D
 9C 60 C6 20 4A FE 33 E5 B8 C7 CD 23 A9 CE FC 4B
 98 6D C4 5A 1E D3 88 E0 B3 BC 36 60 90 14 0E 0D
 1B DB DD F2 8A 2C A9 16 A6 22 8F 26 9C 04 AD A0
 89 32 A6 A5 79 13 BC B0 47 80 B4 58 0C 08 4C 27
 21 86 3E 5E A9 5A 02 6A 90 40 96 D6 1E D4 35 96
 A0 8F 40 45 35 B4 5A B6 49 34 8B 73 65 24 60 7E
 F7 7D 03 FF A9 CC 86 08 6A 4A 07 D0 F1 26 86 9E
 6E 3C 3A 40 92 CB 62 4F F7 12 16 8C 36 40 08 E8
 81 EC A1 18 E0 C3 5E 36 03 77 3D 4B 46 0E F8 78
 2B 55 49 D4 FE 7A 99 97 DC 89 93 35 1B 14 5D C1
 17 02 A4 44 67 A4 E4 B4 54 4A 20 58 8B FB 10 E1
 D1 A6 8D A3 57 22 11 03 64 2F D9 8F 44 3F 29 79
 36 89 CF F9 DA C3 A6 54 BE 73 44 A0 A7 D8 23 48
 52 D3 D0 3F 86 25 B6 22 41 45 5C B7 9B F4 0C 6D
 3E 7C F5 00 9F 1D 98 C3 D2 1E EA 9A 61 52 E8 2A
 96 4A CF 6E E1 7F F0 B4 DF 78 9A 09 E9 97 B9 35
 69 FE 5A FB 06 B4 59 92 57 8A 88 D8 B9 F4 85 DF
 3A 55 7E B0 C2 A3 DC 22 08 94 C4 AF E7 3D 46 29
 C2 F3 96 9B 98 FF A3 CC 34 31 6D D4 B9 44 D1 70
 85 BC 4D 49 2E A5 D7 9D 1E EB 0A CB 35 B9 D0 8D
 4B 6E B0 67 DD 55 C6 6E C8 24 72 D4 19 0C 6F A5
 3F CE 82 CF DA 16 9E 42 E7 9D 09 C5 02 37 48 24
 6B 7A 87 41 39 2A 85 5A 1E 3F 23 6D 87 49 D4 E5
 AF D7 31 4E FC 58 A8 CA 6C EF 69 42 78 56 57 A8
 C8 6D 78 78 1D 15 55 DD 3C F7 D7 0A 36 D7 71 DC
 22 E7 6A 67 45 97 B2 47 9C BD BC 3C C9 D0 56 AA
 67 44 89 D4 B2 A3 7E F0 B0 B0 F9 CE 97 49 A7 8E
 1B 7C 19 9B B2 FD F8 E2 98 7E AF 94 B3 86 7D 4E
 87 A0 07 1D D5 82 34 9C FF 74 7B 1C 77 79 63 43
 09 06 48 42 88 CD 05 62 C1 D9 A5 35 B2 0B F4 BF
 D3 F1 0A 04 31 C0 9B FD 13 24 9E 42 23 1A 70 15
 69 73 41 EE 72 82 43 39 FB F9 A4 A9 6B C4 3F 8B
 77 F4 FC 88 91 25 BA 63 6C 71 6B 2D 57 26 3C DA
 A2 65 33 E9 13 C5 2E 4B EF 2F C6 B6 E6 30 19 87
 73 13 55 0D 1F B8 18 26 24 7F CE 24 76 BD EF F3
 72 F6 82 B0 71 27 0A A6 DD 43 A2 08 4D 6E 42 70
 82 4A 93 AE 18 1F 91 DF DA A2 9A 7D FB CA A7 39
 C7 1C CB 8C 12 95 25 21 AB E5 32 29 D5 9B E2 49
 15 BE 52 44 1D 47 C2 5F FC 8A B5 C4 96 83 14 61
 F8 EA C6 55 E8 7B D4 F3 82 23 DB D2 0B E4 A5 47
 03 2C A1 8A 39 A0 F9 3F CF 89 4C 81 83 92 B3 FC
 0A E7 EA 0A 34 93 C6 C4 E1 B9 26 33 2D 87 53 1B
 4E C4 98 C6 F4 2C 82 92 55 93 F4 6A 8D B9 61 9D
 09 C0 A8 C1 B6 6A 29 3E 54 56 7A FE B6 52 3A D1
 CC 39 C4 08 EF F5 22 5E 2C E9 98 AF D2 24 84 1B
 D9 A9 A1 46 3F FE 61 62 6A AB E8 20 C8 F1 19 D6
 71 D2 FF 78 B0 5D 07 B9 EA 02 9D 79 E6 3F 80 18
 91 8F BD F7 A0 A0 F4 80 A8 90 81 C1 28 BA 37 F2
 8F AC E9 38 95 42 7D 3A 44 37 06 FD C0 5B FE 5C
 30 37 63 D4 1B 0C 5F 68 82 82 CA D0 85 8A 13 5F
 2B 2D BF 64 62 54 58 F8 EF A8 C4 FF A5 E9 20 85
 52 CA 03 DA C8 6C AE 9C 7C D1 0D 84 CE 33 7A 27
 F5 D6 7D C4 CE EE CB CF 6E D7 98 6C A0 8A AF 4C
 9A FD FF 93 87 03 DC 32 A7 C5 40 71 A9 22 53 35
 14 EA 2C A9 76 92 56 F1 B3 E8 43 BA 95 55 D7 02
 09 F8 5E DE 08 4E BC F6 C8 D2 2D 93 C9 4A 07 1E
 6D 8A 21 C7 37 C9 20 83 0E EA 0A CB 1C 8B A6 0F
 B9 B3 C7 DE 08 68 BD AC 3E 87 BC 0F 83 8B A6 92
 3E FB 3C B9 16 D3 62 D9 CF C4 FD 95 0E 34 A2 B8
 CA DB 2F DB 06 1D B9 3E E6 67 28 B2 AA 6C 16 BF
 0C C7 CF CC A5 B5 2A CD 52 7A 67 AE C9 82 E2 4D
 3C 42 86 15 4C C3 DE 20 50 59 68 D3 F3 EB 76 29
 89 E3 81 89 BF 62 63 BD C2 E5 6A 6C EE 10 5F A0
 1E 61 8C 09 C5 E2 B1 97 53 34 D2 FC A0 45 35 E2
 BE 54 28 61 A7 C8 36 BC AE C7 4C BC 23 D4 47 89
 3E D3 DE 2A D1 44 1B 84 3B F1 F7 D9 03 C1 9D 9B
 1E 38 2F 5B 40 A0 90 EA AE 28 21 29 27 59 C7 3C
 ED BA F2 69 D1 13 9C 85 9C 4A A8 6E 18 5E 8C F3
 F0 DE B9 20 51 AF FA 2D 9E 9E CF FA 2A F8 3E 99
 F3 08 E2 5F 8B 96 C8 F5 3F CF 39 91 4B 8B 14 AF
 4F E2 7B 8F 2E F4 5E 9F 05 AB E6 2E B8 48 7F 97
 1E 7C 2D 11 3F 7D 36 D3 73 F4 5E D1 AA F6 EB FC
 3C 3E 9D C8 07 57 59 8E 68 3D A0 CB 7E D6 96 C6
 E0 D7 A6 37 E3 F7 F8 B3 25 89 01 C5 BC E5 2A A7
 BB A2 86 8C 77 2B 72 A5 EB C5 6C 9C 7B 5F E7 CD
 F1 CF B5 A5 58 70 04 B2 72 31 7E 9D 1B 09 D4 D3
 0F 96 3B 82 EC A7 AA 05 F6 03 0E 6D 6E D0 FB 6A
 28 68 1F A5 6C 57 3A 74 6A 82 44 55 E5 40 0C A9
 19 86 3D 72 6B 34 EB 6F D9 56 55 D1 CA FE EE A7
 89 6B 00 2B EC 99 7C 19 D6 B0 D2 E2 6E 84 92 21
 ED E0 9D 23 66 00 1B 2C 7D 96 BC 92 78 65 48 C5
 0B 55 66 F7 5E C3 6B 83 CC 06 88 B9 D5 4C C2 03
 A9 83 93 B7 60 F8 9B 3F 80 E5 FC D3 43 5D 92 D5
 36 58 0D CC D0 7C FF 37 12 BE 0E 8D DB 7C D6 AE
 65 01 8C 32 D3 E0 25 1B 95 E3 99 C2 05 F5 74 49
 D8 63 64 C3 88 EE 8F 23 18 BE DB 7B AB EB 9D DC
 99 48 7E F5 4B C9 FC 26 E4 63 7B 2A C6 C3 91 B4
 4E B3 BE 63 9E 17 49 CC 6D C8 A0 2C 25 47 97 62
 81 EB FE 20 74 AC 78 CA 37 79 AF 37 A4 52 8C 8B
 51 8A 6F C6 89 CA 19 EC 51 2D E3 36 BA 23 63 28
 1D 3E A6 B0 42 79 52 D0 A3 73 2D 0D DF E7 40 B5
 EA FE D5 D9 E4 2E 10 32 7E E3 83 D0 27 62 1E 74
 0A F2 C0 03 2B F5 07 0C B0 85 EB 23 57 FA E6 0D
 24 9E 4E 86 CD D1 7B AE 74 58 87 44 0B 42 85 A2
 33 78 E6 2E 2A E1 F2 14 B9 CF 75 2F 48 61 DD 54
 4F 65 AB BF 4D CE 4B 96 5F 81 2B 87 5E E1 0F D1
 E0 28 21 35 28 B9 ED 5B 9D C0 39 41 79 4B 44 F8
 4F 23 CE B0 70 DC 89 86 5A 3F BE 4C DB F9 02 15
 06 38 55 51 4E 9E 3B 16 D6 84 15 56 89 1A 34 67
 6B BF 49 7C CB 1F 6A E1 69 6B D5 0D 30 41 BD 16
 EA 8A BB 1C 7E 64 A1 D7 4F F2 61 34 EC D3 C9 6F
 F5 73 82 54 A8 82 73 5E 6C 64 FF 50 F2 4F F9 8F
 C1 1A 4B 1F 51 55 4E 65 36 1E D9 7C A6 1F EA 79
 86 1B 51 C8 CE 58 96 05 65 A2 E2 BD 48 C9 89 4F
 76 D2 E7 1D 93 F4 B6 6F 5C 4E E0 B0 B9 17 6F 1B
 21 88 51 7B 2A 17 D7 72 62 9F 13 BA EF 76 CF DE
 84 00 11 AD D0 C6 CA 63 68 25 C7 F3 8A 5E A7 E0
 CC EF 66 23 65 B7 1F 8C 30 F3 A0 B1 CF C8 08 DA
 60 62 86 10 FA B4 3D A5 A1 1C 51 04 A6 5E D5 58
 75 3E 95 9F 73 5B 2B A6 7B E4 17 6B 93 CC B7 47
 66 0E 1C 75 04 9C 19 53 96 DC 96 3B A3 3D 90 AE
 24 C9 0A 07 9F 2C 45 2F 11 45 EC 0A 18 14 60 CD
 BB 2E A5 82 25 B0 13 F9 4D 84 BB A0 A8 DA 2F FB
 62 18 1B BB 45 50 69 D3 CD 09 6C 92 4A EF 8B 94
 BC CE E8 94 05 68 1B 70 7B 18 F2 45 59 CC 64 E5
 14 23 10 E4 0F D5 B4 A4 94 18 AB 68 DE 9F A7 68
 87 02 B7 D1 81 E3 9D 67 B2 78 00 EA 20 64 A4 3C
 18 79 ED 35 4D 0D 2F D5 95 BC 89 AB AF 09 DB D7
 4C 1C 0C 13 42 F0 9C D6 76 35 2D 74 DC CF FC 67
 1F EB A9 A9 B7 0B 7F B9 22 87 1D F4 DA B7 43 20
 30 11 6C EA 85 39 83 78 A2 92 B7 4E F6 B9 55 28
 B1 BB 8B 9E 29 02 15 45 CC 3E AF E9 CA 16 40 8C
 B6 08 A0 75 A4 D3 67 74 D8 6B 3F D5 6B 08 AD D3
 2A D2 EF C9 D5 BE 77 05 3D 0A F0 3A 4E BF 74 CE
 F3 CE 31 6C 99 9A A5 D3 15 3B 5E C2 BA 10 4B D8
 0D 2D 32 04 F9 4F 33 FA 73 CC 40 51 34 D6 DC 2C
 C5 A0 DB 72 D2 E2 F0 BF 83 B1 46 22 95 13 D6 E3
 69 D1 F5 39 8B AD 4E 6F A7 95 55 EF CB 32 51 09
 89 73 46 F1 7E CF 9D 63 C5 48 49 73 86 C5 F7 A1
 B3 2E E3 D7 2D 1B 5C 06 B8 2F E7 FD 6E AB E9 56
 4F 4B A9 3D B4 F1 A3 14 A6 9F F5 45 21 66 41 2A
 B6 F6 02 56 88 86 8F 72 F4 81 9D C8 28 AF EB 80
 03 4F D7 7A 97 2C 47 4B 31 C8 19 80 15 87 FE A6
 E2 01 21 25 50 B5 4E 80 77 33 9B C0 C6 F6 DC 61
 54 7F EF 85 8F 98 07 D5 47 08 04 06 69 65 F7 9B
 B9 EE 29 71 BE 75 2B 02 A4 A3 13 4B 66 CE F6 29
 E9 66 27 C9 6C 98 36 BC 3E E7 DF 7D 28 E5 74 E2
 3B F6 27 C4 A7 63 17 F2 10 D8 2E C3 74 3C C0 F9
 8A ED CD 5D 88 C3 E2 2C A6 14 B1 82 15 45 75 C1
 21 C4 0D E3 00 78 8A AC 53 43 63 2C 36 19 54 93
 AD 74 E9 D1 2B CF 79 99 54 27 3D C8 95 32 81 AB
 74 95 31 BA 9B 62 C6 93 EF 25 1D B3 AC 6C 1D B2
 65 C5 9A 60 B2 84 8F 08 59 26 4F D3 89 5B 72 30
 29 4F 89 4E DC A4 C1 71 AC EB 1C EC 4A A8 39 0F
 9B D9 AA 74 9D E5 03 C8 3B 93 93 1F 7B 14 6B BA
 54 1F D9 7B C6 73 36 54 C7 9A 9C 55 62 10 60 47
 7C 8F 72 D5 78 9C 74 36 D1 8B 22 68 E0 DB C7 83
 D7 5F D3 41 EF 9B 94 57 B9 56 44 E0 E1 E3 36 29
 FC 3A 35 71 4B B0 9D FF 2E AA 02 C7 5A 45 CE 82
 6A 65 E6 5A EE B8 67 2F 9E C1 A5 E5 F8 BC 47 6C
 31 97 8D 9E 9A 1F 09 EE 45 38 26 63 51 ED 61 4D
 A1 36 1B 4E 4C 4C 2A ED 95 D2 D6 9E F9 1C C5 9A
 AD 4D 44 18 2F E3 C9 9C B9 8B C2 28 58 C0 20 A6
 DB 13 22 AD 8A 98 3B 9E 74 97 75 A1 A0 53 58 34
 6A 06 1E 34 15 2B FD 1D 55 76 4E E6 95 79 C3 59
 43 DB EB 5A C2 6F 7D A4 EC AD 2A 54 31 F6 AE 6B
 BA 11 3F 19 59 D4 91 C1 DC CE B8 E7 D4 A9 26 06
 16 27 1F 16 EA FA C9 3D 8E 69 0E 90 E7 E3 46 49
 6C 76 59 EE 5A AA 9A 4C 95 77 AA DA 8E 02 67 84
 BE 51 B0 E8 20 F1 DA CC D0 D0 4A DE 0D 7B 57 20
 0F 90 28 06 2C 91 72 D9 3B 00 15 10 0F 8D 76 61
 B5 A1 6D 44 41 37 44 0F 81 83 E6 E7 40 45 B6 24
 68 B1 B1 F0 32 AD CE ED 4C 72 DE 2A 7F B7 FB 9A
 B9 6A D1 D9 49 9B 4E 1B 6E 25 69 20 43 4C 86 1F
 E6 6F A3 FC 8E D2 04 E4 77 03 80 56 79 F4 35 34
 46 42 65 E4 47 A3 09 28 8C 0B 22 E4 E5 46 29 39
 56 AE 97 29 F8 70 7E 79 7A 7A 0F E7 C4 7B 94 74
 4C EB 9C 8D D9 D9 3D A4 B7 85 85 57 E1 11 A7 08
 81 D6 C7 B3 13 C1 30 9F AD 8C 98 FF 44 63 67 9D
 01 AD 65 0A 1E CC 37 68 A9 00 27 FF 88 00 B9 1F
 64 9E AD 25 88 E0 FB 42 1A 02 2E 81 07 B0 29 37
 2D 9D C2 8C 71 CD F3 1E D9 F2 2F C6 7D 24 AF 71
 49 8F 06 17 DE 47 1F 10 E2 5E B6 B9 56 87 53 51
 66 36 34 9A 57 00 BA 45 49 63 58 52 B3 A7 22 57
 76 26 FA FB 23 5E 1E 74 7F 22 7C 26 5E 47 62 FC
 D6 2E 70 0C 69 53 4E DD 0D B5 03 EB AE 2E EF 3F
 5A E2 51 97 F7 E7 F7 B3 58 4D D8 96 3D 98 04 0E
 9C 28 D5 22 C3 63 8D 64 48 17 40 4D 59 D7 45 26
 06 66 CC 29 2C E6 33 B0 B2 F9 AB DA CC 3B 59 88
 2E 5E F0 AF 71 D4 B4 13 E3 80 42 DE 98 B1 A8 5C
 D5 57 22 7E 0A 86 EA 25 68 64 EC 10 80 DA 1F 0C
 4B BA F0 3F A0 F9 3F 70 98 17 92 E7 AA 45 E5 EA
 C6 7B AE 4B 4A 3E 74 26 E1 4F 1E 9A 45 27 02 7B
 78 C4 9B 0D 0B DC 4B 22 D2 C4 7E 69 39 D9 40 D9
 7E F4 8F 5C 2D 10 B9 53 B2 40 57 41 D7 49 80 8E
 42 17 EF 62 E0 AC 83 D6 DF D6 8F 87 C8 AF 58 86
 EC DA 01 E7 FA 11 7C A8 4A 7D 3B 12 DF 01 6C ED
 C7 13 D0 F4 7D 20 34 F3 25 B9 4D 04 FC 2C 6F 68
 E5 FE 97 7C 11 01 C8 49 7E CD C5 A9 F7 02 07 E2
 73 6A 6A 07 F5 E4 33 13 B0 62 88 71 70 92 20 46
 CF 9D 5B D2 83 04 85 E1 E7 26 50 E2 FC 61 8C C2
 49 61 25 4A 4F 5B 14 27 88 C6 8C 29 55 EA 52 F8
 F5 4C FF B9 3E 08 47 57 20 77 F7 E0 14 AC 17 81
 F7 B5 0E F2 82 D5 EB 82 5C 0A 82 1D FD D2 D7 8E
 F6 D8 93 26 B8 D1 FD 20 77 25 0E FF B4 EA E0 E7
 18 73 EA 7F 7B 46 A2 21 84 C6 75 B1 30 9D 52 F6
 2C CA 06 7A D8 32 03 FF F0 09 78 70 7C A6 F3 ED
 61 31 30 8A AE 7E 77 2D D4 11 BC 8C 02 6C 1D 3E
 46 34 FD 9D 0F CB 73 12 B3 B4 FE 18 F5 0C 5E 06
 85 CB 41 12 52 96 9E 60 FA FB BF 49 B8 11 50 A4
 5B BF 77 40 5E B1 81 A6 05 48 CF 75 C1 CE 8D 55
 29 6B 20 E5 01 C2 0A 10 DA 3D C2 13 85 29 A2 26
 E1 0D BC F2 C8 5A E1 78 D9 79 BF E5 C1 9E EB B1
 A5 F3 43 5B E5 51 26 91 A1 2E 6E 7A 26 87 17 2C
 7B 05 56 0E 7A 50 D0 16 B0 70 B1 9B 31 4F F6 7D
 91 42 96 CA D5 46 D2 2B B3 9A 39 89 6E BA C8 D2
 EB 3A 82 C1 1A 7B 91 E8 4C 29 50 33 C0 2E A9 45
 22 D3 07 64 11 E2 DF 2C D4 83 37 64 B9 FB 99 5D
 AD 6C A6 96 1C FD A7 98 4D E6 DC 95 8A 5F 92 0D
 A8 1E D3 F4 09 F1 38 5E 49 19 46 D6 43 3D 7B 10
 9A 95 55 21 65 28 26 8A 73 03 52 64 31 78 31 F5
 83 7C D7 68 67 B1 36 AB EC 07 BC 06 4B AC 96 12
 0F 87 BC 35 19 9D AB 0C 21 94 50 1B 4F CA C0 47
 08 D5 42 C8 07 7B 0B 26 96 1A 07 7F BA 34 B2 32
 31 0B DC 05 01 77 6C 46 FA 16 28 42 72 ED E5 92
 AD 49 A8 6F BF DA A5 35 3C 41 C4 F0 AB 8A 4C DF
 7C 3D 55 B6 CA 7E 2E D7 50 2B 4A 26 B6 B0 0E A1
 17 48 FA 3D 9F EC 4B 9B 42 17 16 F5 BD E5 7D 84
 EA FD 93 E2 DB 62 1B FC 73 4E 34 BD 34 AD 20 9C
 92 D5 42 61 06 01 56 A4 EC 2E D7 89 47 B6 E7 02
 7C 9B 94 41 A9 EF EF 2E 1D D6 DA EF 4D 05 FD 43
 9A 72 1A EC 88 A4 1E D4 E5 E8 83 57 15 DB B9 E5
 AA 7A 18 89 4E 9C AF EE 74 1C 2B 6B 12 34 D6 37
 C0 BE C3 82 6A 42 50 61 8E F8 B9 EC EC 17 40 26
 27 04 3C 9A 16 E9 2F CA 6E 03 95 5A AE 90 04 49
 14 B5 EC 75 15 F8 D7 88 70 24 37 AE CD C3 22 CF
 1D 82 AB 94 AD 2A 46 FB 7D 32 7E 94 14 80 CF 7C
 15 6D A0 D7 08 FF 6F C6 34 94 41 1D 25 47 BD F9
 A4 45 D7 0E 5A AA C2 5E C6 C5 15 3E DC AD 45 F0
 62 46 67 62 C9 11 68 E6 D0 41 95 D4 EA 61 D7 EA
 FF FE 73 FC F2 E4 D3 C7 EA 2F 23 D1 CF AA 66 08
 47 EC A2 6D 6F CC 50 B4 4B B2 32 AD C3 0D 09 0F
 78 51 03 55 94 B9 D7 73 03 A7 58 E6 1D B9 C4 84
 4E 7F AD 0D 08 F7 51 C5 15 FC 37 65 1D 3A FF 9C
 21 82 D8 E3 61 EC B4 88 0A A1 7B 75 E0 C5 01 A7
 FE F4 18 55 F3 2F F2 02 60 6F AD 1D B0 BE 98 56
 17 73 35 B8 94 4B F9 C8 B9 CA A8 3D F5 29 E6 EE
 73 F4 E1 12 99 7D 4F 8E 22 C9 80 46 7F 3F 9C 37
 EA 1E 13 12 23 D4 63 18 A9 C5 A1 82 28 3D 02 78
 FF 24 50 88 5B 88 56 58 3F D8 89 44 32 4D 58 7F
 A3 B5 90 EA 9F 96 BB 28 0B 20 37 DE 59 CC AA 04
 3C D3 A2 33 12 8A 92 E3 A8 E7 93 21 DE 77 A6 AF
 7A BC 43 7F 58 E6 5C 6F 8C 9F 38 EE F1 1E F5 BE
 F6 95 2B F4 14 B4 7F 0A 11 93 4A 8A 34 30 45 FF
 BD 79 6B 9A 76 C7 CF 5B 14 BE D3 4A A0 47 EC 76
 80 EE 1D 06 9B E8 86 8F 49 9A F0 5B EB 19 7A 6F
 A8 50 27 D6 6F B3 C0 2A 2E 70 7D 42 19 8D 6B 8C
 66 26 56 87 CD 7E 5B 78 E5 D3 6E 9E 73 90 6D CA
 05 D8 90 33 3A 6C 0B 78 B0 66 2E ED C6 D7 7D 34
 5A 78 BB 8F D0 7F 2A 27 B8 97 1C EE 87 31 43 0E
 D4 22 C9 59 0B 0B 8B 06 05 97 86 3B 10 7C 5C 90
 D2 E7 94 BE DC D7 AD 9E CE 46 C4 BA 97 9F 2F 94
 CA 4E CE 22 FE 06 2A A3 57 6C A9 D2 8A D9 FC 7B
 50 41 1D FF 6D AC 9A AB 2B 55 36 2B 98 97 C8 20
 D4 14 82 E1 22 D8 50 29 9F F0 FA B2 A1 55 62 A4
 A8 E4 6F 7E 9E 5F 0E 2B 6D 87 1F 2F D4 68 5B 77
 60 B2 20 64 A6 BC 05 24 56 A9 3E F0 36 C2 D8 DF
 19 91 28 EB D3 0F 09 C5 55 5F 2E 56 80 00 C7 04
 80 02 8B E3 13 3F B7 F6 6E B4 8D BE AE D3 CD EA
 B1 69 9F 82 B3 CD 67 19 9B 57 73 F0 81 21 FA EA
 2C 28 1D 95 1C 1A B1 C1 3A 93 56 93 4A D3 FC 15
 A1 CC F5 82 11 29 17 37 69 44 FF CC F3 9C 64 73
 A2 E6 A5 FC 05 43 F1 E8 76 E5 49 7B 9C 63 4B 2A
 9F 00 1F 47 53 BC 07 35 38 45 56 B6 C4 F0 4F 6E
 2E 6D E2 D3 56 C1 4A 44 1C 00 C6 9D 6C 1E 10 5F
 8F 9A 1C 89 B4 06 8D DC 3B A1 47 F9 8F F8 33 6B
 0E 7A 79 41 84 74 04 47 DF 20 76 38 DB 67 B3 C5
 AF 47 F7 E8 22 47 34 2D 37 75 1F D3 FF DD 07 CD
 E3 6C 3D 5F 88 54 4B 91 BA 1A 66 88 00 CB 67 44
 C5 69 58 77 30 26 71 D2 A7 C0 3E 81 09 F5 8F FD
 28 5B FC 78 AF 0F A1 7E 12 10 01 42 19 5D 3D 26
 D5 AA 74 DE 91 48 02 05 08 E3 0F 62 E3 15 C4 AA
 61 C4 9D 03 15 7D 02 8D D1 BF 11 64 0C A8 36 E6
 71 C2 71 FC DE B1 FC D2 B3 25 B0 8C B0 B3 32 36
 90 F1 0A A9 AB 56 79 3B 52 4D BF 0C 65 B3 FB AD
 26 1E 69 F9 D0 A2 12 19 FA AF 7D BB C9 ED 8D E9
 8D 16 DE 77 17 17 FE B4 77 9D 4B 1E 53 2E 81 5F
 20 B2 FE 8E D9 13 47 C3 40 6A E5 9B A2 E5 33 20
 14 CB 97 88 1C 70 FB F2 E9 7F D7 E5 DD 86 66 BE
 87 17 9B CD A1 BE C8 48 8C E4 A8 54 C1 3A CC 77
 27 7E 01 2C E4 47 B4 71 CD 0E 51 44 84 17 5A 01
 1F AE 43 30 54 A3 41 75 C6 5A 5B 36 75 ED 77 32
 A2 0F 8A A4 46 DD 39 72 C2 AD 9F 9D B4 CE 02 4F
 EF E0 45 69 36 AD C3 6D 82 8C 98 59 09 15 5D 46
 CB ED DD 80 6A BC F0 2A 68 80 5D BD 9C 91 D5 DD
 C2 BA FA 78 74 F4 7B 0E 25 0C CB 4A 48 DA B5 CA
 68 B6 D3 68 43 36 18 28 45 BA 3B D8 B4 8A 53 BC
 B3 DF 93 BB 57 25 C9 09 15 D8 AD 57 BE E4 6A 3B
 BD 27 AE C1 C6 2C EE B5 9C 36 83 C6 F5 27 D0 62
 A3 B2 FD C3 8E 87 B9 4C 76 C2 7A 49 0A 1E 1C 78
 7D 3E 69 7F 99 64 01 B4 07 E4 DB D8 D9 A7 DC 7E
 62 2B 42 9E BC AB 7C A3 E0 29 17 CF 1F D2 2A 7A
 D4 0C AC E2 9C C2 F9 2D C4 9B 17 FD 3C 42 E7 9C
 26 B2 68 08 95 FF 81 8C A7 44 E2 B7 BD AA 39 97
 6D F1 31 1F 41 C3 77 52 AF 0D BE E9 24 E2 BD 4A
 C4 89 6B 66 19 D1 5E 3B 7A 4C 44 0E 62 37 4A 02
 27 40 B1 5B 52 4C 26 04 23 B3 FC F1 84 49 45 4B
 BC 44 EA 34 AA 02 B2 81 A1 25 5B 0F 67 1F 4B FF
 7B EF 44 63 23 E6 75 0F B8 12 48 8D B1 62 02 20
 23 22 07 4F 35 5C 48 71 A0 9F 11 99 CD 32 5A AC
 E2 41 5C 6A AD 45 90 5D AD 97 57 8A 98 C7 AA 2F
 3B 88 E2 B3 D2 C9 3D 6C 8C EB DE 0F 46 71 0C 15
 A3 E9 F3 25 E5 18 08 0C F4 42 F1 B8 74 59 6E 53
 14 C5 A8 22 62 CA 16 69 A5 6C DD 59 E5 34 D1 2F
 62 88 DC 3D 4C CC DB E2 CB 95 1B BD 6F 5E 71 67
 3B 2F A2 66 BA E3 07 47 DB 62 07 68 E8 37 49 78
 DB A4 96 B5 74 B9 50 31 78 F3 8A 44 D4 3F 8A E0
 62 2F AB 42 0C D3 CC B1 4F 54 83 4F 92 8F EC 39
 A6 FA 01 CA EC F1 FA 23 1C 63 35 EB 50 3A 79 5B
 F2 53 52 ED 7D 27 E7 76 E6 BD F2 0C 74 C6 FD 63
 74 49 16 EF 63 1A 76 B6 61 F3 CF 21 73 3F AC 6B
 3D 3D FD 1D 4D 66 D1 0F 9B D7 CA 9F C1 1E BE 2C
 CD 08 B2 1C 61 3A 81 1B A7 6D 82 F9 E1 F5 13 CE
 30 EF B1 D1 E8 25 AC F8 46 CF 6C 06 3E 78 76 74
 F5 9B A4 AA DB 23 E0 7E 88 5F 75 D5 29 74 AE 70
 D8 4C 50 57 12 C7 EA D9 35 53 89 6F 9B A0 4A D4
 66 70 3F 08 F4 0D 6A B3 C3 83 B1 03 DE 3D D1 CB
 A6 9E 62 94 2F 5B BA 38 96 D8 E0 C2 E9 40 44 79
 68 18 91 FE 05 59 5E E3 5B 2C 58 17 D1 A8 66 2B
 CC 16 E8 6E 35 86 82 03 38 1F 4D 6A A6 10 B4 75
 47 B1 73 47 88 C4 C6 4A C2 F4 49 9A F1 31 DF 9F
 8B B0 13 BA 41 8E 9B D6 89 D2 28 DD 43 A7 F9 B0
 88 05 AB 90 8E A6 C4 CC 25 DC 69 C6 C1 AD E7 55
 A5 07 94 F1 41 9E 36 26 67 83 97 EC CF C7 ED C3
 9D 90 66 74 09 4E CD 5F 05 11 BD 6E 14 4A BF 72
 E2 41 1F 1F 09 A7 63 1F E8 F5 50 9F 4A 1E B3 0B
 33 5B 20 D2 FA E5 74 47 5C 3C 29 6F 8C 5F 3F 6D
 27 F5 4B 88 64 DE 64 36 DA 4E 6A B4 68 7F 3A 0B
 71 66 94 6D 2C 3E 15 50 27 F9 66 2D A8 41 8F 3A
 DB 53 18 6A 6D 17 2C 82 34 A7 FC 8D 6C 85 C6 62
 3A A1 55 07 1A BC C9 D6 2D 41 DD EE CA 99 A5 2A
 4C 26 79 33 FD 34 C2 E0 9D 88 55 97 DF 5B 20 2E
 90 7F FF CE 32 E7 88 B4 30 ED 8B C8 11 00 7E EB
 F7 A6 49 B5 1C CD AF 27 7E 4D 8C 0B 18 A0 81 5C
 45 9E 6B 4D EB 4C 59 24 66 28 93 11 DA DD 0A D9
 E8 16 92 8D F0 32 47 34 02 04 9C 35 E6 0A 65 4D
 CC D3 59 83 4E BB B2 6B 2A 9A 97 28 D9 64 9E C8
 B8 3A 3F 49 B6 35 31 0F 34 69 BA 58 FA 8E B5 36
 92 F5 24 14 47 25 38 4A AB CD E8 60 DA 25 DE 15
 44 2E 1F 87 C2 DB 59 62 D2 5F B7 70 7C D4 84 D0
 32 5C DF 26 98 01 32 09 A1 11 5C 9E 1E 85 02 25
 C1 E6 B8 83 B4 7A 1E CA C1 7D 8F 83 80 4A 5C E3
 95 1F C3 29 0F 52 B5 62 F7 B4 99 5C B0 87 60 75
 81 4C 9E DC 42 4B 6D 23 DD 95 EE 7D 4A CB 40 EC
 F1 7B 9E AD 1D 47 06 E0 CB 92 67 BA 88 C2 D2 7A
 31 AB 0D BC 0C 3D E0 06 94 E1 CD 66 94 53 3F 73
 06 85 0E A7 79 9F 96 35 A0 12 12 38 49 0B 75 CD
 C5 91 A3 46 94 8F B1 58 E6 A8 F5 69 EF 13 9A B9
 2F 9C 54 AD EE 0E 95 49 9D AE AF D0 DF 7D 3F 29
 B9 E0 B3 6F D1 16 13 C8 FB 91 F2 63 75 4C 90 4E
 30 E7 02 64 9F 79 EC 86 AB 34 0A 51 A6 AF F4 13
 AC F4 67 9C 55 62 72 62 E6 70 38 26 92 77 ED E8
 E4 2A 1C 6A 4A 22 BB 7B C2 11 67 73 A7 FC 3B AB
 41 93 21 9A 33 42 44 2C 27 CD 37 7F 4F 80 17 22
 A4 90 4E F6 37 F8 4F 60 7D 22 34 F6 2B 61 ED 64
 53 96 94 2D D7 16 C0 63 D8 85 01 AE CC D1 9E 01
 51 82 F4 57 62 A4 B8 21 C9 D5 30 A1 C2 38 E0 50
 9A A8 48 C0 46 75 5B 7C 4F 5D B2 FC 27 7F 98 A4
 1F 2B F5 0C 31 9D CC A2 5B B1 62 B1 7F 1D 6C 32
 2F EF AB F7 C6 02 68 E4 51 84 A4 7C C9 77 A7 15
 0E 9A E5 EB 29 01 D2 D9 76 8C 7F D6 BC 28 74 4F
 B3 FB 2D EF 9E 2A B5 86 BC 8E 8C A8 A5 B5 1B 44
 88 86 FA F6 D2 1F E9 E1 47 00 36 08 C2 49 5B 5E
 DD 91 71 94 D5 CA 75 0D 0D D2 10 04 2D A0 C9 AD
 38 70 FD 59 70 A1 EC 30 80 E4 3C A0 7D 72 79 B3
 54 89 15 86 FC 76 4F B2 D7 95 C6 9F 60 A8 09 49
 68 2C 83 54 3D 19 AC 74 2E 70 D2 5B 87 82 1C 09
 D5 AB 93 83 BC 11 39 42 84 65 21 BF 79 E4 05 0C
 8E 32 57 7E DB 7D 2F 90 B8 45 32 07 DC 81 3D 5B
 BC 8F D0 76 D1 67 CD 70 BF 59 BF 70 EF 3D EE 32
 2C EB 16 D9 1C 0A 61 72 06 0D EB F2 71 5A F2 82
 BB 97 5A 15 E2 56 1A 55 BE 35 39 56 CD ED 43 FB
 47 BC 64 57 61 90 E2 B1 9C 8B 20 9A DF FF 01 32
 3A DD 10 05 DE AC 25 90 B0 F9 59 E2 7B 63 2B 8B
 28 86 E7 2D 08 E4 81 8C D3 3A 55 FE A5 50 2D 3B
 9F 1F 4A B7 96 D8 8E 3D 47 91 ED 9A 15 14 35 E4
 E2 CE 69 33 1F C9 5F 43 D0 BD 38 DD 27 13 5D B5
 4D 94 05 E9 1D F6 D9 6D 11 3F 2A F7 8F 10 DA F0
 A7 CE B4 09 B1 B1 BD 33 0E 2C 92 6A 12 36 CD 6C
 FD F4 65 5B D6 B6 33 81 73 C1 C0 3C BE 77 AA 6B
 FC BC 04 54 16 E6 52 97 C7 42 F4 BB 56 95 FC 0D
 60 BE A4 E4 51 25 C4 E3 04 CD 9E 69 6A BB A5 5E
 4A 61 B9 6A FF 64 8E 35 3D D3 F1 DD D1 AC E6 F8
 B0 37 B3 17 E5 7B 44 75 86 88 B4 D2 EF EA D5 95
 B7 B1 36 9E A3 26 0F 73 36 2A C3 4D 98 55 6A EB
 52 29 03 D5 45 12 7C 02 8B BD E6 4D 45 6D 57 43
 49 EB 29 67 23 FC DD C4 07 67 E7 EC 2D F7 88 E3
 B5 FB 63 88 CA 5C BD EA 06 9F EE AE 2F FE 7C 8B
 1B 15 01 D0 F0 4B 90 F8 B0 A8 37 B2 A4 A5 A6 16
 38 30 1C 8C 62 1E 18 83 6A 5E 06 1D D9 1E 81 A9
 73 3F 17 2E 5A 40 DF CE 40 11 34 63 D0 70 8A 64
 D4 E3 65 00 78 4B E0 DD 01 C0 C3 09 4B 70 8E 8C
 B2 75 4F 34 5C 81 04 34 AA 13 2E D6 96 63 80 43
 4A A4 AC 7A B8 12 59 F4 83 3E 6D 28 1E 93 74 D5
 26 51 6F 60 A7 AF FF 72 74 31 6E 99 1C 09 AA 1C
 9C 5F 1E EA 50 F5 F2 FE 42 CE 80 C2 73 F6 53 E8
 7D F8 9E FE 0A 64 0C E5 89 24 E6 EF C5 12 A6 05
 91 50 2A 55 75 87 6B FC 18 E7 6A DF AA 61 82 FF
 A4 D1 17 75 C1 27 C3 C3 16 A5 64 56 6C 76 AB 8D
 1F F5 5A F7 77 86 74 28 D3 AB A1 63 43 0B B2 7E
 19 83 5C AD B5 4C 77 10 53 CA 3E 96 4D D6 D7 AD
 0B 7E CB 0E 3F AB C0 F4 37 9E 74 BA 07 31 53 72
 54 BA 84 BE 56 AA F0 1A 5E AF 5D 03 29 11 18 53
 4F E7 51 9C 10 AC 30 29 CF 2C 61 34 9C 8A 8D 47
 52 58 6A A7 AF C7 E5 9C 9E D1 D8 A5 BA FE 46 FB
 AA E4 83 62 DE C3 27 14 1F 7E F9 A0 9A 48 7C 6F
 3B 38 03 1A 85 41 A7 78 8C 9D 95 72 8D 01 2C E6
 A6 5F A6 04 DB BF B2 E6 82 8F 26 1F 1E 4C BD C8
 5F E6 DC BE 68 2C CF 54 FC CA 17 92 02 36 5B D7
 15 7A 0C 12 32 4D D5 1A 40 6C D0 01 B5 46 11 4B
 A2 55 C5 69 DF F3 28 6E 08 0D BE 7B CC 69 19 77
 7B 19 B1 BB 81 C9 A7 58 63 39 D0 6B F7 49 35 2A
 B9 8B E4 10 8A 4E 37 C4 09 01 7F E1 39 4E 96 CB
 1B 89 18 B8 B4 DA 01 C2 E3 1F 69 11 27 1F A8 8C
 80 B7 E7 AE CB F4 6B F5 CD 9E 2F FC 5B 7E 6D 74
 1E BE FE F8 52 00 3D 9A CE 28 F9 F3 25 C8 E6 18
 E3 53 0B 6D C8 2D F9 68 86 2F 04 56 B1 9E 0D 4E
 DA 46 F0 6E 96 E0 D2 96 01 5D C8 24 D8 58 AA 0B
 D6 A9 12 63 31 FA A1 BB 97 BD D0 52 9F 24 44 AE
 A3 0B 1B 38 16 29 76 34 68 43 01 0A 3A 46 37 BE
 2C 55 26 5F 2A E9 FD D8 BF DB 53 B4 FC 0C 34 3D
 77 82 80 40 5E 25 3A 0C 78 48 4D F1 14 95 C1 E5
 31 8C ED B7 3F 13 28 3E AD F1 CC 62 18 6F 5F 35
 63 E1 5E AF BF 65 6C 26 00 70 61 33 F5 2C 2E A2
 D3 2B F9 14 7E 02 17 D9 9B FF 7F 21 EA 31 6F 87
 0E FD 7E C8 6C 18 D5 5E 72 90 FB CC D1 18 0D F7
 45 FA 12 6B EB 0C 4A 29 44 B3 54 F4 3A C3 9E 1F
 EF 75 57 FA 38 6B F0 71 61 0D 06 5A D1 B9 EA A0
 D7 19 99 49 86 78 09 79 84 F0 04 5D 8C 2A A0 D1
 15 F6 0B B4 1E EA E3 8E 5D EF B7 E2 C8 5F 70 4D
 74 7D EB 93 43 19 56 DE 5F 57 02 EF 42 FC 82 0F
 30 EB CB FF 0A C3 D3 1F 53 D1 D7 CE E6 53 FA 99
 CB 6D 76 42 CD 1F 85 10 6C 08 59 CA BE 9E F9 10
 06 6E 4F 70 72 12 9F E9 A4 A9 65 84 8D 83 CE 24
 97 9E 8E 79 BF 60 37 30 45 CF 87 2D 90 E5 44 52
 48 08 05 5D 2D D4 5B F7 5F F5 E4 8B AD 2A 3B 26
 2C 84 97 AF DC 36 E4 3F 3F C6 8A 93 BE FC F6 F9
 0D 7C DE F5 F1 13 42 63 07 B6 D9 F9 A3 E1 BA 16
 B8 F9 15 9F AC 88 D8 65 C0 94 43 4B 66 11 9B 33
 8D DB DB 4E 64 79 27 8C 9D 34 79 0A 12 09 66 B6
 CA C9 96 6F EA 12 85 C1 9E 68 E2 51 23 A4 F6 FE
 7F 3B 84 ED 45 44 57 7C B1 46 1D 8C 49 2F 07 79
 61 9D 04 6C 93 04 98 D1 3F 59 DA B1 39 A1 48 64
 84 47 61 CC 2A 0A BE 17 AC BA 85 1D C4 FA AC C0
 9E 5F 0E 33 04 00 96 84 5E C5 FE 2A 8E CB BF 69
 0C 7E 6D E8 D2 14 0C 0A DB 24 D9 48 6B 8A AA 69
 FC 52 44 52 0F D4 B1 5C 68 CD 60 0D 2C BE EC 24
 3B 45 70 8C BD 2F 0A 1D 68 5F 98 13 20 0F C5 BA
 61 3C 8B 4B 78 B5 91 46 83 5E 85 95 64 0E 27 F8
 AF B9 B8 AF FC C6 51 37 CF 4A A2 EB BE 12 81 BF
 07 29 D6 7C 14 BB 58 01 63 7F C6 89 FA BA 6B FC
 08 09 1D BA 90 79 0E CF 4D 3B 98 12 DA 23 5C 3F
 6A C1 7D 4B 31 B3 FF C5 94 C7 03 0C 82 E4 6E 80
 80 CE 30 16 E2 25 E9 41 DB 66 77 1F B6 C2 9E A9
 F0 39 1D 8F 60 AD 94 2F 7F 18 8E 52 B9 83 26 37
 CE FD 43 60 D0 FA 45 E0 15 51 3B E2 37 B7 08 B2
 92 BC ED 38 73 E6 58 71 1D AC B0 FC 5E 55 6D 5A
 BC DC D5 14 17 36 07 38 F0 D1 54 42 7A 73 62 01
 01 D1 1D 0A 7D E6 02 35 E9 D5 B8 6D D9 D9 70 B8
 DB 64 88 15 23 95 C0 6B 65 A5 BA 02 4E D6 5C 53
 2C 8B 22 F6 4F 37 F3 DE 5A 06 E0 42 60 A0 42 EA
 FF FC AC B9 BC 5F F2 1A 89 97 B2 72 89 74 15 1E
 3E 7D 9F 8E FF 04 D0 A2 E7 BE 9B CE 43 C4 4A 11
 4A CE 6D 1C 7D 07 38 35 9C AE 8C D5 62 9F 49 1A
 92 BF 37 6E DA BC DA 44 C8 25 72 39 13 24 FF B6
 0C 71 75 D4 51 E7 FC 1A B0 66 2E 36 3E C5 FF 76
 43 F2 84 E2 2A C5 61 B6 F2 F5 94 5D E5 4C B9 FB
 3D 11 39 86 22 7C 98 8E E1 BF AB 4A FA A6 CC B4
 BB CA E0 52 60 8F 3B 52 F3 34 5B 60 FF 0C 64 EC
 99 5E 9C 88 32 D3 5C 34 8D DE 0A F5 5E C8 CE 8A
 9E E4 E8 59 1E 96 B8 EA 72 51 A2 2F 7E FC 3F 56
 DE 45 9C 65 AF 09 52 77 F2 BD 20 51 5A 4E 3D 04
 92 36 67 1B BF C9 4C 7C 3B BE 90 A4 E4 D0 F4 29
 C3 D3 49 AC F9 EB 0C 5F ED 38 2A 5A 79 71 0A F4
 27 B8 25 DF 99 1A 53 43 FE FE 65 C1 95 93 ED 16
 7D 50 DE AC 0D 90 19 2E F9 AC FE 3A 55 A8 F2 A1
 8E D0 E7 6D 0A 13 34 BE 2C 09 AE 8A 22 72 3B 97
 D0 8E 4D C9 34 1B 06 04 A8 9D 55 29 AE CE 3E 0D
 44 37 38 B6 53 8F DB 90 9E 78 9B 92 68 FE 18 C3
 0C 8D A3 56 22 9A 3B 47 D4 E6 02 34 BB 25 61 D1
 1E BA F0 94 34 9E 51 EE AB 1F DB E0 E1 B9 4D 4D
 1B 8C 2B B8 F7 D7 F9 91 53 CE C1 8C 62 8F 50 7D
 07 BA 42 6D 4C A3 BF A6 ED EC 37 9B 3E 9F 5B 7F
 9D 54 83 48 6F 27 13 70 D7 D1 A5 07 11 DE 41 3F
 C9 7D 80 FF D9 19 9D 0E 84 3E CF DB 97 26 65 4F
 51 A2 E9 18 B3 6F 2A 9C DD B9 91 9C 3C 28 CA F6
 50 A7 77 47 AE 84 F5 8C 0A 02 A1 A8 8B 20 18 21
 5F EA 1D 2D ED C7 46 39 F1 73 9C 40 77 89 C0 BA
 16 48 61 C3 F7 55 90 CA 6E C4 68 6C 71 3E 04 F5
 B0 5C DD 1A 29 0B 9E 7C 0F 62 1B 8D FE 8D F6 52
 16 F0 E8 25 30 33 F9 18 31 39 EA 46 F5 DA 80 67
 1B 76 4F 72 69 84 F6 09 25 6A F8 99 0C F9 0B 5E
 1E 8D BC C9 B4 9C AA D8 B6 04 68 0A 85 36 3E EC
 57 41 BC E4 BB 74 0E BB A5 F0 31 25 D5 ED 99 1E
 76 7B AF DF 30 3F 9B DF 77 65 8E C5 F5 D3 84 22
 47 3D 62 52 20 45 3F F6 F9 66 64 01 D8 B4 52 86
 75 75 DF AA 12 68 A2 99 83 BC 24 EE 15 C9 75 F4
 52 79 0A CE 2C 29 03 22 0B FB 8D 24 EC 17 BC 0F
 82 6E F7 3B 11 7D 71 83 7D 5A 16 9E 1B AE 34 39
 A4 E7 15 20 A7 0E 69 F0 F5 02 EE 98 BE E5 4F D0
 3F F6 64 B2 FE 50 95 AC 40 76 D3 F4 13 2D 85 7B
 95 29 6C 52 DA FB 98 62 F8 1C B7 4D F5 9B A8 CC
 F2 07 67 DC 44 B1 94 74 43 18 42 08 D5 79 2F DD
 B1 2D 08 A6 D9 5D 2A D7 F2 76 D9 B5 2E 23 E9 5B
 82 FE C8 A8 47 F3 94 96 06 EB 1E B3 5B ED 2C 63
 74 1D A9 B1 7B AF 9F ED 7E 89 41 31 6E 2A AE CD
 1F 9F 8C F0 5A D8 DE A5 0D F5 97 74 50 ED B0 9C
 71 DF 7A B8 23 71 50 7A AE 7D 03 04 A1 88 3F 9A
 72 16 6E 1A 96 28 3B 0C 94 DA B0 38 03 69 AC 4D
 39 DF EF DA 9E 79 A7 7B 53 09 88 37 53 C5 C1 43
 85 DF 46 A9 F6 FD 75 88 8C 1E 52 D1 20 EE CC 22
 C1 BE 16 84 C5 E5 C3 FF 9C 26 C9 0F A1 7F B8 FB
 D9 81 38 2E DF 1E 56 C1 8F 39 F0 39 B4 DA C5 01
 09 60 40 E1 85 D8 1C FB C0 B5 2C 27 85 22 37 28
 33 19 62 30 62 02 32 B5 F7 94 F9 9E DE 02 97 AC
 42 FE 8D D0 D8 11 72 3D 39 F4 68 F7 68 75 35 54
 68 0A 21 82 61 70 6F 2E 6E 0E C7 29 42 B6 E7 44
 32 BE D8 60 F5 C8 07 2B E8 91 34 A8 74 DB 96 53
 18 B5 CA 6A 45 3B 80 BB F5 12 A7 6F 89 0F FD B6
 5E C8 F7 FE 44 33 AF D8 8B 10 A1 87 A7 AE 2F 5C
 3C 6B F7 65 F5 20 7D D6 67 CB 51 D7 4E 66 30 ED
 27 8D A1 1A DC 06 CD E1 8C 00 F3 CC EB CE 66 0B
 A0 5E 06 5C C2 4D 1D B0 4F DD 13 B0 7C 65 34 ED
 0D 61 8C 1F 46 4B 8F FA C0 66 D6 79 17 B9 ED 3C
 FF CA C4 0D AE 0A 6C 4E 9F 4A 59 7F BC 5B 0D 35
 89 4D D3 43 F0 D2 CC 33 1E 76 18 ED A6 36 2E 66
 F2 DB 6A 09 82 92 14 EC E8 8A 60 97 E3 88 C0 09
 CA 05 17 60 13 70 E9 EC C9 10 1B EB E6 FE 00 64
 A2 25 74 01 0E 46 8D D2 14 20 3B FC 1A 2E 46 8D
 BB B1 54 52 D4 5C 12 14 31 40 A3 A9 D0 16 AC 6C
 1F 7A E7 B4 C3 F6 D1 43 24 22 20 9A 53 5D 37 0B
 EC AA 68 C2 F8 DC B6 10 2A D2 E9 2D 9A 3C 7E F3
 0C 8B 9F 64 47 AA D9 3A 0C 0F A5 45 84 E4 3A E0
 E0 B4 02 51 20 90 26 22 9E 19 0A 9F 1D E6 BC D1
 A4 A8 8D 5B B7 2B E2 B6 0E 40 7A 9E 02 75 0E 37
 55 BE A5 CC 6A 5E 1E CA 57 93 B7 2F BF E9 5A 8C
 85 63 05 E9 6E BA EF 1C 6A DE 0A 46 89 E0 18 FD
 85 12 B8 A1 DB FD 55 B9 DC 3D ED 28 63 6A 8F 0F
 38 6E 09 1B 93 44 0A 51 A3 BF CD FE AC E3 9A 61
 1C 22 83 07 39 8F 52 E5 24 81 AF 83 D5 6F D7 7B
 A0 C5 8B 25 9A 74 49 32 6A C7 2E 00 9D 74 2E B2
 0C 78 1B 3D B1 D1 A7 58 27 27 E3 12 36 EB 67 82
 91 07 BD 24 D9 3A E2 60 03 C8 49 82 C4 95 64 E7
 80 F0 6B 45 A8 1F A0 1D AD F0 18 DC F8 D1 D8 BB
 C1 9D F9 9C 97 DE DA 04 63 A4 63 94 48 5C D9 CC
 52 8D 01 1E 11 E4 1B 81 91 88 DF FD 5F E0 C3 02
 62 78 62 E2 C0 1D 81 71 34 E6 ED CF 5F 76 49 2D
 E6 49 F3 D6 0D 6D C1 C1 83 90 11 A0 A3 62 16 46
 C4 F9 58 8E 76 9B 77 2A A8 9D 0E AF 1E 19 63 1E
 D8 08 49 88 12 18 3D 82 A0 5C 14 80 EF 40 BD 79
 8E 1E 32 AC 14 01 4F D2 26 57 D6 74 18 1E 43 1A
 77 6F B1 53 38 34 7C 82 84 3B 45 55 FA CA 09 75
 61 08 D0 52 1A 66 53 34 A0 F7 20 9C F5 B0 F0 28
 3A AF 00 4E AB 23 57 1B 5C 44 1B 8B 43 13 11 C1
 80 63 15 90 CB B3 14 AD BE 91 E0 4F 84 76 1E 4A
 4A 89 52 3D 19 A2 11 E7 D6 7B 05 87 B8 91 15 37
 D5 FB 17 35 BD 64 22 1E E8 C6 69 BC 7E E4 C4 37
 A5 58 65 C2 41 5D DF B0 DC 06 1B 94 F6 CD E5 A4
 C6 19 2F C4 F8 B2 46 30 82 5F A8 9C 84 F7 AD E8
 38 DA AC CD A5 A3 35 DC 1A 71 2A C6 A9 D0 41 75
 0B 43 BB FF E4 DC A2 95 E6 5D 97 04 42 29 EB FD
 2E 62 B1 A6 CE C3 97 13 6D DE C5 A0 23 E5 8A 86
 A9 39 AF 40 01 2B 3B B4 CC 7F 83 AF 0E BA 14 E4
 85 D9 58 48 E8 C3 DA EE 8F 2D 23 A5 BB 9A 6F F4
 72 9D F2 11 10 CF D8 E1 0B 0E EF 88 5B 0C A0 43
 22 40 1C B6 9F BC F2 CE 0E 96 51 B8 12 12 B4 FF
 30 E6 9A 60 05 BA 9A AC 9F 7B C6 0C CC F0 80 5B
 D6 0A C2 E8 F5 9D D3 99 D7 E4 DE C2 A8 42 7D 5D
 5B 50 7C 1B F8 AE 5D A4 A7 FA CE 23 7F 8D 7F 5D
 1F 70 66 BF 98 55 51 B7 13 94 0B 63 75 5D 73 36
 74 29 27 A8 B4 6A 5F EE D8 74 E9 B2 F4 F9 39 1B
 41 00 C5 5D 08 FE 40 70 76 B9 1C 91 06 A4 3F 49
 BD 92 16 14 1F 10 5C B2 13 1B ED 7E D1 05 13 46
 87 93 03 83 BC 62 D2 A7 58 EF 90 C2 E5 1C B3 FB
 55 68 D7 74 32 4B FC 5A 11 7A 4B 2D 7A C6 97 F8
 08 D9 4C D4 B1 25 F2 79 75 CA DA C1 B5 D4 0E 9F
 17 26 87 9A 43 04 61 49 2F 2C 7A F0 1F 84 26 B8
 03 9B 50 D9 DB 43 3C 2A 50 AF F3 B0 AC 52 45 5F
 5A A8 39 A1 D0 BB 0F 4F A7 DF 3B 2B BE 74 FB 3D
 8E 14 45 07 79 62 3E BB 14 E0 94 EB 0A C6 1F 66
 BE C4 6B B5 5A 93 57 49 B3 19 BA B8 EC 68 3A 4D
 D2 1A 1D 89 B1 CF EA 13 B6 2B B4 D0 ED EB D7 19
 18 35 5B 76 DE 87 D5 72 B1 14 0A 37 F5 85 A1 23
 C1 80 B0 66 7A 0C 81 BF B3 95 46 FE B3 7E 21 FC
 8B AC 70 7F 04 46 55 77 72 83 11 D2 7C 5C 1B CF
 A5 4F F1 13 7D AC 16 3E 1B 72 1E 5F CD 58 1A A2
 AA 1F 57 8C 50 1A FA E2 D7 40 B3 84 70 D1 49 2B
 18 11 FB 0D 34 43 6D E1 09 34 D3 03 5F A3 AA A0
 16 E8 E2 D4 74 78 92 EE 8D 06 56 65 2F 28 AC 8D
 11 D8 FE CE 83 C6 87 CB A1 BE F4 74 12 70 29 9B
 FC 48 1B 6D 27 73 5D 85 5F 3C 31 93 EF E8 82 8A
 6C 39 CB 44 D8 24 28 12 D3 6F D7 52 7B 93 EC 2C
 7A 7F 23 99 92 1E B0 8E 75 02 96 04 B0 D4 FF 97
 BE 2B 62 52 BD CE FF 08 47 5E 32 18 F6 A3 98 E8
 97 6A 47 6F 81 03 1B 06 98 71 21 CE F8 00 EE CB
 D3 3E 2A 5F 72 51 0E AD 8E E9 94 36 6D 73 82 E2
 02 E5 4B 80 62 EA 22 78 E4 27 F7 82 F4 3B 99 58
 D6 24 54 31 1A 5F 2A E8 34 A9 99 B4 F7 C6 74 DB
 A3 F5 C3 E0 AA 11 86 18 E2 79 65 53 5C DC C1 4D
 2A AB 4A 48 03 4C B2 08 A7 9A B7 8F FD B0 4B 62
 58 10 B5 FD E6 83 22 85 11 D4 0A 8F 03 AB 5E F2
 74 C1 E3 4D C4 18 A1 64 9A 2E 97 E3 9E F4 B5 3E
 18 74 5E 65 8D 6B 1C FF 25 30 27 96 7A D7 EE DA
 97 58 F1 A8 1F B9 7F A8 AC B4 CF 16 3D 83 11 C5
 7D 0B 11 12 2B D2 B9 0D 0E 0E 31 DF AA E7 CF 65
 97 06 D8 5C EF EB 6E 71 6F 24 F4 DA 40 BA E7 4E
 6E 7E BB E5 D0 48 95 8C BA 27 00 D6 3E 32 8F 17
 AF D9 A2 FF 32 A2 43 07 6B 9B AF 77 98 C5 0E EB
 5A 7B F0 2D 32 50 8E 38 E5 C5 20 6B E8 4A 92 B6
 DD 6F 1D C7 90 89 68 98 63 0B F1 17 B5 AA 4C 65
 4E 98 C0 8B 63 16 8E 94 3B 51 53 04 0E 8B BA 76
 F3 9F 71 29 D6 18 06 BA C1 70 92 20 4A 2A E7 41
 D4 E6 3B C8 29 D0 1D 23 C9 4E 9E 05 A6 D1 D9 73
 DE 76 A1 00 32 30 58 CC DC A7 73 6D F1 74 1D 73
 6E 8D 93 89 11 49 7A 87 4C 27 61 9C B5 01 A3 30
 B9 9C 2A 9C 93 C7 36 BC 6C 63 99 53 90 AE 79 56
 B8 2F CC 99 CB 9C 8C D9 58 B3 00 54 D3 1D C8 0E
 1C BA 3F 19 28 38 20 91 2F E3 8F F2 BB 58 83 90
 0C 17 D5 B8 52 1A 03 6C EC 43 2A 47 01 DE 9D 38
 41 13 B9 F0 2F DD 3B 1B D8 B4 A0 AD B5 2C 04 6B
 C3 8D 3A 12 75 74 CD 3E 27 45 CD 60 7A 42 D0 E4
 D0 3E 5D F3 7B CB 11 62 17 6F C5 CD 55 4C F2 F2
 6E F6 63 DD 65 E5 72 12 8D AE FC 66 4C 70 5F FC
 9E A9 0F 57 1D C0 84 39 D0 A5 76 39 58 69 FD A3
 0E 44 F7 FA 09 AD 43 00 95 B2 E6 1B 06 FB FF 05
 68 76 6C 23 D0 B9 BC 74 A7 77 EE 00 6A 07 26 08
 8E 7A A5 38 7F F6 E9 B0 69 14 73 04 F1 D5 CC 71
 DF 91 81 C8 CA 18 EB 22 F8 BE 46 78 A6 34 04 41
 FE 9E CD A7 A2 24 47 2C 3F 55 42 D1 84 38 5A 88
 32 85 94 7F FC 21 E1 16 CA 85 25 E5 F3 15 0E 8F
 80 01 4C 83 FC CC 1D E0 8D A6 38 A4 88 9F A7 71
 BE 7A 05 99 08 00 4A 4C 27 7E 57 9D D3 3A C3 80
 4B 92 1C FA BC AE C2 35 FE F1 FD 04 66 A4 A1 C2
 7F BD F9 42 B8 3A 00 43 86 83 2B 6C 79 04 FA FE
 6D 39 4F 16 AD BF 59 A6 E5 6E 37 BF 33 88 4A D6
 07 0D 5E A7 FD 2C E4 EE C7 40 80 B5 B7 99 D8 58
 33 B0 DA 1D E9 C5 52 42 20 AB E0 37 AD ED 81 0E
 BC 31 50 00 4D 6F B7 14 2C 92 A8 F7 B8 DA 97 3C
 79 9E 6A CD FC DC 9B 3A F4 CD D8 5C 83 94 4E 3A
 BB E1 DF 9D CB 46 85 8D 2D 85 3A 19 AF 72 BE 1F
 00 51 24 19 DA CF BF 4F 93 E1 6A E0 AE 0B 06 16
 4E 09 65 F6 9B 07 4D 0D 8F E4 AC F2 A8 7F 04 FF
 4E 10 60 2E 39 8A 19 3B 38 16 A3 C6 82 1B 43 D6
 4D 97 62 13 0A E8 8A 57 64 7F 56 43 CD 22 73 A2
 DF AD 85 A9 35 34 1D AF C8 55 C8 57 21 9B F5 0C
 19 C7 7D BF CB B5 2B 5F E4 25 53 3A D4 D2 A4 0F
 BE C6 5D 00 54 18 33 25 6A 4C 38 99 13 20 3E 2A
 A2 26 80 9F 1A 05 77 03 75 82 9D AF 45 7C 51 4E
 91 18 17 26 89 D6 21 5E 3C 7E 19 BB C0 02 B0 98
 77 4D 2B E9 7F 5C D1 63 7E 01 F0 20 71 AA 63 07
 FB 0F A5 2C BF 2A C4 6B 32 48 1D 47 2A 9A D9 C1
 C6 C5 5E 5C 6F 0F AB ED 4B 54 17 FB 74 9E B6 B7
 7D A6 75 31 74 10 6D 5F AC FD 39 6D 56 79 1B 0E
 26 49 97 A0 14 2A EC 58 E0 CF DB 8F 0D 87 1A 9A
 14 52 CD 32 F0 0B C9 6F A1 63 62 28 7E 7E 10 4F
 60 2F C5 24 64 6F 2E 93 7E F7 31 08 0B 7D B5 9B
 FD 49 01 0B 20 0D 40 15 49 C3 EF C6 A6 A9 A4 72
 17 68 F4 20 EC B5 96 60 86 C5 4C DB D3 CC 22 50
 B2 3B 1A F6 C0 BD 93 23 98 7C B7 A8 4F C9 7A E8
 D0 9A DA A6 67 25 EF 40 FB 4D BC 1E DB 33 95 BE
 C4 AA 43 14 2C 41 FA 2A 83 B8 46 8F 87 26 4D 76
 8C 87 AE 2C 87 EC 21 2C 5B 1F 44 63 67 F1 9F 0E
 12 DC 55 B7 E6 90 59 3C BC 11 95 44 6A 55 FB 73
 5F CD F1 AA 65 DC 70 90 3C DA 23 55 32 0B 59 79
 D3 85 D3 57 23 E1 17 59 5E 1A 2C CE 44 A8 2C 07
 D8 E6 83 D8 3A 56 88 82 2D 29 3F C6 83 2D 56 7B
 A4 D7 51 FB 1D 41 6E 30 50 9D A4 3F 34 2E 91 CC
 46 C5 17 37 63 1C 09 D2 DF E2 C4 49 75 E6 9E E5
 34 F2 B5 7D 0A D4 96 70 55 E5 E1 57 91 10 24 C3
 5C 5D DD 4E C0 BB D5 CC 0A 9B 9C 95 4E D7 42 E7
 1C 69 B9 4A 4D 48 44 1E 75 CF 51 08 98 D9 2E CA
 A2 E7 25 CA 26 53 A0 D4 65 27 86 EC E4 2E 2C 22
 CF 2B 48 60 79 65 55 2A 17 AC 84 1B 64 6C DF 72
 66 60 50 34 21 FD 2D CD 2B F9 A0 E6 BF 83 B5 4E
 5E 42 11 70 0B EC 72 4A 4E 99 13 8D 46 25 61 DE
 13 80 D3 F6 38 FC A1 79 89 3E B6 20 6E 87 DE 2C
 4D 74 2A 67 6B C5 5D 21 38 24 5E 86 7A 55 DC E9
 BA C3 6E 73 65 1C 85 58 87 42 26 FB 7B B5 C0 D2
 13 76 5C E1 11 46 82 CD AC 72 2D F7 3F 08 5B BE
 27 30 D5 FC 63 88 85 FB A5 CE 74 96 47 8C 80 46
 F4 4B FB F1 08 CC 22 8B 62 21 E7 55 24 F9 B9 C6
 BB A1 D5 2E F6 60 D3 D6 C5 8F 8D E0 F4 67 0A 76
 A3 A4 1A CE B0 E6 C3 5B 7A 14 88 A7 37 43 E5 F5
 AE B6 A3 1E 42 8B 46 EB 43 67 0E 93 92 4A 50 4D
 50 61 E2 C9 F5 9F 89 6A 47 F0 2F 7B D8 85 2C 7E
 9C DB AC 50 F4 FB E0 EA 28 B9 7B E6 9E 21 B5 E8
 55 1C 7B 2A 4E D6 22 22 D6 D5 67 39 E8 09 F0 F7
 94 68 A8 2D E0 51 DB CD BD E1 24 BE 62 9D 1F 8F
 E6 49 C9 5C 84 5D 20 A8 2A 80 89 EC 41 A8 7D 82
 B9 C3 05 2A 2E 91 D6 C7 4F E2 F3 7E B7 4D F5 F9
 48 7D D5 75 43 4D 5B 0A 90 85 34 C3 EE D1 B1 16
 23 AB EF 57 67 B9 4F 32 49 DE 06 97 D0 7F EF DB
 DC D7 38 41 C6 13 D7 4C FA 55 1F 2D 3E 35 D7 60
 53 EC CD 53 5F A1 FD C4 E8 B7 7F D2 9B 05 E9 02
 2C 2B 42 33 90 C7 84 F1 0D 93 6A A7 4A B7 23 85
 4D 76 72 2A 9F A8 1C F3 10 4A BD 66 A2 A3 18 3C
 BC 65 16 06 89 6E 35 B2 80 4C 7E 52 95 EA 9A 48
 F0 1C E1 CF A4 A9 73 DB F0 22 F3 AD 0F CC 52 92
 0C DE A6 23 F7 26 A2 D1 35 8A A0 E4 5D BE 51 04
 32 91 49 A0 25 B8 46 EB 66 B3 95 39 11 D4 CC 9F
 26 F8 EB 2C 5D 69 B8 8D 99 1B 0E 31 A5 FA 77 7E
 E9 F7 89 54 77 DD 02 A8 2B B5 4A 6A 79 BD 99 2C
 3B 61 9F 79 05 52 BA E9 09 3A 30 0D F2 0C 55 F0
 26 20 AD 6B 13 90 AC 15 2E C0 CD 0A A3 64 4F 1B
 70 56 36 F0 70 BC 8A 34 67 62 C8 BF 95 32 E4 91
 FD 07 CF C2 16 E6 BE 9E 9C 29 0A 2D EA 94 10 A8
 43 B1 FE CC 07 95 7E 73 A9 DE 1B 65 B9 35 09 0E
 9D 77 EC E5 9C 40 E3 6E 8E 8A 0B 56 81 D5 AC 1C
 1D 00 59 0A 23 62 39 0D D5 D6 A6 34 94 43 4C 62
 40 6C 79 9A E7 BD 3E 40 80 70 6B EC A3 3F 10 26
 FE 9D 92 BD CE 5E 0C 28 2D 78 66 A1 F8 92 F0 CE
 78 6C EA B0 BC EB 92 86 BA 61 3E D2 5F E4 6D 0F
 B6 15 D1 22 EE 1D 12 E7 98 49 E8 55 0B 2D 4F 74
 41 6A A6 F9 7D 76 CC E7 67 BC AC E2 71 56 12 B9
 2D 16 4E 02 3A 8A B0 20 6B A1 CD 5F 98 DD 86 CF
 4B 6A 58 DD 09 A3 C5 DA A1 A6 DC B1 1E AA 27 BF
 33 39 CB E5 95 9E 1B 92 F2 5D 93 18 BA 00 59 5C
 1A 64 33 D4 46 6F 17 1E BD 00 AF 5C A1 3C 48 0A
 49 6D 8A 35 F8 D6 67 14 F3 81 77 E3 79 8F 6A 60
 AC 11 9B 82 75 28 4C 7B A2 97 10 4C 22 E6 4D C7
 C2 98 D6 B2 0D 4C E3 C9 01 28 3D 28 8E ED AA AD
 0A E2 4E FB F0 71 1C 1B FA 04 31 29 5E 0A 6C 9D
 DD 64 18 B1 09 5C A0 CD 2B 48 67 E8 C4 E9 0D 5D
 68 5A 49 E0 51 A9 9A 7B E1 81 70 8D 08 D6 91 B3
 5C F2 4C D1 09 CE 2D 4E C0 CF CF 7C D9 41 CF A2
 02 18 AE 6E 15 44 28 73 07 76 5F 9E 40 F0 63 6C
 77 E2 5E 7A 53 0E E6 AB 13 33 28 8C 57 5A 9F DD
 75 75 D7 0F 0E 54 5C 54 11 CD EC 20 95 4F 70 6E
 0E 0B 88 84 25 FA B2 AB 70 C1 9B 6A F9 F4 B8 6F
 02 76 21 2A 94 5A 56 5B 93 4E 72 32 3C 7A 9A 0A
 EF 0D 78 21 95 50 20 A6 95 B1 C1 8C AF DE 1F D7
 0A F3 90 5C 5A 3A 42 A9 C4 9F 6B 64 D4 E7 04 BD
 6B AC C1 5F 3E 15 3F 2A 78 07 7B 94 54 D3 1F 85
 AC 00 D9 59 78 90 BC 91 4D 62 88 23 5C 89 3E 33
 20 93 FD 2A B1 35 73 03 16 FE 1C 54 3B 99 AB F4
 0F CB 60 BE 78 AA D9 E2 04 75 F9 30 8B 3E D1 24
 93 26 7A B0 84 1B 47 33 10 11 C1 D2 1D 94 B7 54
 2F FF EC 62 16 B2 B2 E9 47 20 23 05 7E 42 82 5F
 8E 6B F2 AB 73 84 91 33 55 05 08 16 51 D9 C5 F8
 23 A2 B3 10 45 7C AF B4 D4 72 C3 28 DC 62 DF 27
 2E 3B 48 DA DB CA 12 31 D4 72 C9 53 5C B3 62 74
 3B 28 1A AA 71 D7 EF D0 EB BE DF 0C 4A 80 8E A4
 F7 5D 84 E1 26 FC C8 5F DF BA 7C 23 B4 42 8C FC
 4D 6D 63 39 AE 17 FE ED DF B1 5C B9 17 2A F8 6E
 F2 40 86 AF 6F D0 52 F3 71 9A 0F A6 5B 5A 43 84
 50 66 6F DE F1 37 CE 7C 20 38 23 D8 DB 5C B4 A2
 98 3D 48 45 30 33 6B 4E 86 DE 7C 00 6A EA 41 A9
 DD 70 93 BC EF 23 88 F8 70 59 C7 E3 B7 95 E2 EF
 DC 5B C4 58 CF 48 CD 9B 77 C0 72 52 77 9A F0 59
 B1 FB 36 BF FC A2 5A C0 6F 8D 24 D1 02 26 DA E7
 FD 06 11 98 66 15 4A E3 AB 04 24 D3 02 DE 5A 9A
 33 A0 53 C5 BE 39 C3 D8 56 32 F9 80 BF 1B B5 CB
 01 26 86 A1 94 72 82 C1 1D 62 CA CB B9 9E B8 6D
 A4 57 7C CE AB C1 B5 49 B2 4C 9B BA CD 77 63 CD
 39 1E 0E 00 24 D2 4F 20 A4 CA 37 99 1A 7B B0 72
 60 00 AA 83 1E 0B B1 FA C7 A0 21 78 4C 51 74 B4
 87 77 DF DC EE 6D E6 6D E4 D9 91 1F CF A4 65 CF
 1B E9 0B 74 36 9D C1 56 31 8B 3B 01 94 22 DD 30
 07 88 DA 45 98 DE 48 3F BB 0D 51 C8 EF B6 AE 03
 9F 73 61 A5 82 FB BC 4B 3A 39 FB E8 AF 4C 15 DC
 10 7D F1 86 FE 9C A4 16 CE 4E 5D 96 24 65 08 39
 F8 04 BA 40 D3 84 E7 C8 55 95 EA F7 81 3E FC 16
 44 37 B4 60 5D 80 F8 F7 94 70 3C 14 F6 89 59 DA
 10 40 AE 5A 3B 62 53 1D 20 4D 2F 5A 5F D3 68 38
 BE 97 8C 1B 7E D8 5D 2B F2 1A A3 43 D1 C7 AE 4B
 C8 B8 A8 CD C9 5F E6 71 9E 4C E0 3C 99 6C 4B 93
 70 52 A2 7A BD EF E5 01 2F 23 50 CD C2 9B 57 EF
 FF 75 9D 37 9B 77 85 50 35 1C FE EF D3 79 C4 B0
 7E 38 CF 6E BB B7 67 BB 2F 3D 49 88 BD 17 EF 5F
 3B D0 2E 91 23 7D F8 5B 36 8C 50 18 46 55 23 4C
 55 39 F0 B8 CF 75 D6 B3 9A B5 DC 83 8A C2 07 84
 36 56 02 66 C5 B8 AD 86 45 B2 0D D7 2D C6 8C C5
 53 13 30 D4 C0 27 BB 52 28 29 6C 9C EE 92 C5 F4
 AA EE 96 17 59 68 F1 FC 4D AA 2F 7D 83 9B FB 22
 D6 D0 2D E5 11 AD 58 93 57 BB B9 43 42 DD A2 F9
 F1 16 81 64 DE C0 B9 ED 03 AA D5 A8 E2 96 C2 80
 13 DF AE E7 CB 56 FC 66 9A 7D C8 C3 37 D5 55 D5
 55 B8 5B ED E4 F8 75 97 CD DD 57 7C 9B 52 0D EF
 71 05 33 72 0D 0D 8F 30 9A 06 6E 5C 9F F1 97 A0
 E8 9D 53 98 19 68 A5 F4 17 E2 41 8A 28 D1 0B 19
 62 CC 25 14 80 50 C5 D4 05 FF EF FF 09 2F 00 CE
 3F 93 19 23 66 7A 79 42 AC 8F 1D A3 2D 11 C5 89
 39 51 81 3B 4D D9 8E BC B7 33 FD A0 E4 F4 F3 E5
 0B D8 C1 92 97 91 21 AC A7 14 19 F1 1D 9A 22 88
 7A 58 AB CC 8A EE 0F 1C 1E 7D 7C 0E E0 20 D3 FB
 08 5C 49 ED 46 B5 A2 D3 9C C4 41 8A 41 B4 9C A0
 8D 5B 96 71 3B E1 39 9D 5D B8 05 E4 58 6F 5C 2F
 8A 27 0A E0 2D 6B 53 29 83 41 22 BF 79 5A 96 18
 15 2E 0A EF 49 9C B4 0A 70 45 D5 EE DA 79 9E F6
 FE AE 48 3C DB 5A E4 48 44 DC D3 85 23 E3 7C DA
 B8 2D E2 69 89 FC 1E 4B DD 5D 35 EF 66 EC B7 41
 7F 8F F1 CD 43 5D EC 24 8A DA 4C 7E 31 DC 35 8F
 1F C0 18 62 F2 93 93 D3 24 C8 DC CA C8 F6 A8 87
 44 51 C5 2C AD 98 48 F7 22 1A 3D BF EE E8 4F 5C
 7E 38 C4 8D DE 8C B2 47 C8 A2 75 B8 68 A3 2C AF
 59 57 A2 30 BD E8 D7 C2 F7 5D C0 E0 3C DF E8 C5
 C6 A2 8F 16 48 1E 2A AE BB 46 F2 A3 69 DC A3 30
 54 FA CC C9 67 C1 CD 86 FF 73 24 16 E9 5B B4 CE
 66 47 C2 FE D8 3E 01 58 6E 6C 59 43 E0 11 21 66
 21 E5 41 DC 0C 78 3D 7E 8B 4A 60 64 8C 43 22 07
 82 19 DD FB AB 7E 1C 5E 65 BB 5E 7E 8D 6D EC D1
 D6 9F 0B F3 71 E9 D3 B3 D7 49 F9 C0 09 E9 7A F3
 E5 3D 06 BC A5 9E D8 E6 FA E4 71 7B 34 40 B8 D7
 81 DA 00 59 F8 6F 38 3E 9C 58 93 39 63 E1 5D 80
 2E FF BB DB 08 34 1A B8 DF 27 80 5D EC EC 81 F9
 CB 57 BF BC 84 98 1A 12 62 73 A2 C1 54 31 CB 41
 2C B4 AD 28 5A 57 46 1B 6F 2C D0 EC 64 67 74 07
 6C FD E4 B1 AE 4F 01 5F B7 B9 13 0C 1F 2E 1F 4B
 19 F8 0E 15 73 EC 63 EC 05 67 7B 80 C3 D9 C5 75
 F4 F6 79 72 31 24 DA A4 51 13 1A AB C2 9A AB 54
 FF F7 7A 1E CA 03 E0 4E 03 9C 1D 90 CE A1 26 31
 F9 DC 4E EE DD 43 CD B2 F1 47 BA AE AE 17 9A 35
 F9 C0 F7 6A D1 2B E1 18 E7 13 4C D0 9E 17 AD D1
 B3 16 86 E5 7F 5F 19 F4 85 7A 72 B2 5B A4 1E 6E
 E4 3F DE 7C ED 56 A0 54 9F C2 A7 F4 83 81 40 78
 0A C8 B7 4A F5 EB 7B 1F D1 5A 26 56 75 66 0C 4C
 44 64 83 B4 19 A4 98 CA B4 0A 52 DC A1 C7 5F 2E
 42 FB 4B 88 C6 A1 F0 CD 35 C3 7C 72 0C 34 BD B2
 55 5E E4 80 FD 1E 14 9E 4C BF CE 5A A9 D7 9B 17
 7B 3A D2 67 0E B9 F2 7E 62 6B EE CF D5 9F 61 BB
 53 48 F8 8F 13 E3 C5 B3 B3 EE 8E 56 42 60 3E 58
 F3 AD E3 3D 1F B4 B0 45 8E F2 44 DB B5 94 6A C4
 99 96 76 CE 39 69 FF 35 EA C9 86 82 8F DC 7C EB
 E3 62 7A 22 09 19 E1 26 4D 2B 11 53 19 12 BF BF
 CF DD AE CD 4A E0 CF D5 C5 23 20 70 16 59 E0 1E
 25 48 27 C6 F4 0E 4E AD 43 BA 5A A8 8B 3E CB C9
 BE 93 44 AE 3E 9A 8D 2D A9 8D 5F 22 09 A1 70 3E
 A6 90 03 14 6F C5 2B 73 60 49 85 22 3C 68 C8 92
 1E 75 5D 6C 0A 59 93 D5 DA E9 15 E9 11 2F 93 A9
 87 4E B8 BB C7 5C EE DE A4 0E 1C 6B CE 4E AB D9
 34 1D B2 0F C4 C8 8A 15 CF D3 97 3D 74 E2 E4 76
 D9 B7 96 FB 2E 70 BF 67 5C 21 92 24 BC 6B D2 58
 44 D7 7D 8C BA 8D 48 C6 C5 01 73 11 7A 2A E7 44
 88 9C 08 99 4B 79 71 AA 05 E7 F5 99 25 C7 B4 C2
 E3 C0 4B 3D 2F 36 8A EC D5 75 56 6E F4 01 87 14
 E1 47 31 13 A0 A4 0E D0 6F 0B 79 2F 3F AE 1F 70
 D0 90 A7 FF C0 A6 2D 73 6A E7 B8 45 AA B0 E0 69
 E8 25 D8 51 09 04 1C 7D F9 C4 75 89 09 DC 14 F2
 7B 04 4B C0 BF 12 80 6D 93 79 12 96 AF A2 A3 9A
 13 85 0B 1B 0D B4 B4 5C EA 36 84 B1 2C 85 06 7D
 DB 7C 9C 36 4A C1 B0 AB 2C DF 16 1D 19 9C DB 7B
 13 1B 13 36 5E EA EB 71 1C E0 19 74 C7 E3 C7 BA
 01 1B C1 10 C5 F1 2E 0F BD 43 87 42 47 EC 9C AA
 C8 37 8E 9B EE 40 F4 95 16 31 34 8A B2 4E 62 76
 BF C5 D8 C2 71 B4 C7 35 45 99 65 3C DA 1F CE 04
 06 F3 19 DC 2D D7 FE 5A C1 EB 90 22 3D E4 36 41
 79 05 FC 97 E1 F9 6B B9 C6 FE 02 49 FB 05 8C 9B
 E3 E2 47 E8 E7 CC 2B C6 FE 3D 6D 2D 3B 9A 33 9E
 03 26 B0 19 AA 80 68 04 60 0B 33 3B 4C C2 1A 2C
 55 88 21 76 30 8B B4 64 9F 39 71 F7 AC 88 4E 7D
 0A 2E 5E 57 EB B4 A6 1E 20 57 68 F5 25 D4 F5 86
 27 10 6B B0 16 DB 94 58 2F 4B 3B 03 C3 6D 73 B6
 D0 6E E4 AE 5B F6 7E 4E DA 22 19 71 7A DB 9B FC
 20 B3 A2 4D F1 E0 A3 94 96 C0 AA 2C 38 B0 73 86
 62 34 F8 98 40 32 53 CF E0 A3 92 93 EA A8 F9 6A
 64 38 10 D4 36 DF D2 9E E6 DA 33 B4 A8 64 8E 22
 7C ED F5 92 E1 16 67 DF BE 5E 16 A0 77 87 DF E3
 FB 4F 6A B6 15 C5 C6 4B 01 B1 44 81 A5 97 8E 1D
 FC 16 93 CA E6 09 9F 2B BB 1C 9A 1F 01 27 31 1D
 26 81 EB EF 3C 41 C4 C4 08 DE 83 26 FF 08 6C 8C
 75 91 EE E5 58 73 7A D7 8C B9 38 F7 1A 97 79 4B
 1E 37 F6 D8 2E 48 F7 47 1F 75 28 CC D5 F1 DD 23
 F2 90 09 97 AE CB EF E4 12 6A CF 2D 63 44 6E 5C
 88 2B 44 82 6C 60 E0 A9 F8 8D 00 DB E6 50 5F 83
 D2 FF 5E 3E F4 48 D9 C4 FB C3 89 A2 59 A9 04 16
 15 70 13 3B EA 18 97 2D 93 38 D2 F1 99 78 5A 31
 EB D6 B4 45 53 37 96 83 77 33 16 98 A9 B4 40 1D
 0F 91 41 D2 08 CD B1 B4 A3 D6 FB 42 6A 88 B2 A0
 0A 33 6E 91 2E 81 CC 6E 8E 65 E8 04 13 95 79 15
 32 39 56 D2 3D F8 BE 77 D7 70 19 1B 81 E9 62 30
 8D 6C B5 91 FC 3B 9C 45 BC D9 EA 54 58 4B 5B A7
 BF B4 88 21 E9 9E E1 02 08 F9 AF AA 4F 86 00 AA
 9F 28 31 CA FA FD 33 56 C4 62 56 00 58 17 43 8F
 FF 3F 62 DB 45 F8 31 87 5D 28 D2 CB 7E CB 46 3E
 AD 28 1C D2 E3 DC 7E 69 C5 74 05 93 E7 E6 0D B0
 34 D2 E5 66 6A 2F 0F 3E D3 DC 65 0D C4 1A 65 A6
 3C 76 37 BE 31 92 02 86 25 30 CC B8 73 95 3F 29
 D8 7C 04 95 3D B3 B5 71 17 C1 BD F7 4A 66 1E 0F
 37 A2 F9 5D E0 5D 5E 28 04 D9 15 AF 97 5B 5F C1
 AC 18 A0 BD 4B EE AF F6 F6 25 4D 50 6D 10 29 55
 EE 6E EB B6 1C 76 E0 DB B0 D0 F7 24 55 D0 49 6D
 3F 8D 0A E1 14 E8 B9 DE 08 12 79 04 5E E6 33 F6
 1B 35 C6 26 D8 C2 67 05 49 58 05 7A 8D B8 6C 7C
 88 3F A0 5C FA 89 5D 70 13 36 E0 65 35 E7 4C 17
 09 40 53 42 FC 2D A6 18 C7 E4 CA 03 C4 C1 2A CA
 04 E4 74 54 53 CB AE EA D4 3C 54 6E A4 86 51 30
 1F BE 12 18 04 7C 36 76 ED 45 8D 92 6F CF 2A 14
 6F DF 87 B1 9B 12 59 A9 B4 66 7A ED 02 10 3C 25
 8A 13 57 C6 74 68 26 01 38 54 49 AA FA D3 FB 17
 B8 FC CB 84 07 DE 06 3E E0 E1 6D 6A FC AF 95 28
 51 3D 0E 1C 38 9E BC E0 6C 1C AF 80 13 C3 81 B0
 E6 98 E9 E6 FE 7F 15 41 2D 99 9F 52 F0 BA 00 AE
 AE FF AC 2D D4 CE A6 75 3E 27 FC 82 52 5F 26 66
 9B F5 C9 89 EA 07 EE 31 96 F5 F1 08 E7 CD EC 01
 55 F0 68 06 01 4E AF B1 83 61 C6 0B A1 5D 5B F4
 68 7F 03 2F D0 CB B3 57 0E 86 E6 D7 79 E4 98 41
 12 1A DF DE 84 B0 2D ED 44 83 11 AD C8 F0 3A 6A
 5F C7 E4 72 EE 2B EB 9C 0A 22 37 0A 10 80 AD 84
 92 B7 17 4A 06 88 2C 3F 36 F8 49 1E 30 23 B3 2D
 20 D8 AA 1B B3 40 10 15 1F A7 DD 73 A4 E6 A7 3D
 E8 5E 8A 15 80 1A A6 36 74 AA 02 4A 94 7F 37 EF
 37 4E 79 14 09 1F CB 7D E1 E0 CD DF 1C 24 7C 4B
 9C E6 D5 10 19 E0 EC D4 71 F7 36 D5 CB B2 1E 35
 24 EC 1C D3 B1 95 84 F9 6D 68 46 61 D6 F0 0E F6
 68 4E ED CB C7 9D FE C5 E2 41 3C 9A FC C3 96 96
 29 1C AC AF 8C 72 4D 92 34 29 C2 03 FC 83 A8 9B
 4F 67 D4 F4 6E 5B C8 E6 47 71 4B 85 29 43 11 2C
 F3 9E 39 C7 2B 18 5E 08 2D 53 CA 0C 09 F5 70 61
 C3 D8 EC 07 59 E1 8B F9 99 73 CA 3F 26 5B 00 AC
 C4 4B D6 A1 A7 18 88 01 CD C9 3F 1F 60 CE 20 85
 7D FE D3 14 1F AB 5E 54 F7 E2 DB A7 4E 58 25 8E
 B3 6F AC EE B5 06 44 98 D4 3D 4E 80 76 D4 6C 6A
 E9 3E 1B B0 E0 FE 50 2E 55 2C 4F 7F 45 ED 6B 63
 E4 94 B2 A7 C2 79 B6 FF 97 69 E8 33 C5 65 4B 54
 CE C7 54 7D F4 11 02 59 56 15 A7 24 9A D5 45 A2
 C0 B5 98 0C F6 D1 B2 58 CE C0 64 C0 14 2A BD 0E
 42 A9 99 0F C3 CC 17 70 6A 94 08 8B F5 22 13 8F
 28 2D 55 90 13 E7 2D F8 5A 29 A1 99 7C 78 AD 8B
 5E 7B 62 4D B0 8A 6D 6D 59 A7 CB C5 29 2A 38 16
 AF FD D0 27 BE 12 F0 85 1A 5C 6C 7E 00 A7 89 C5
 A4 2E 83 F9 F7 F6 02 34 77 FA 76 73 BA 59 96 42
 1A E7 4E D7 A5 C0 B9 52 8D AB A8 40 C3 F6 66 A7
 EC 12 CD B7 25 2B 0A 51 5C 70 5A DD 94 18 8E 0F
 34 95 6B 23 F9 45 3C 40 8F 5D D1 39 0D 78 F0 7B
 AF 0C A4 B9 7D 0F 50 2D 8A 02 BC 4D B1 9C F1 63
 E1 65 8C 92 94 55 91 18 B2 CD E0 FA C9 2D 83 67
 D1 5D DD 42 44 27 F0 AF E5 CD BA EE E2 A5 D6 73
 99 45 A3 EC 5B D7 22 E2 9E 99 37 B9 71 46 AD 06
 0F 8C 2E C5 A6 97 B6 A1 8F CC 3D 83 C2 61 E3 01
 BF 13 CE 05 85 05 E9 D4 A3 9D DB D7 99 29 52 D0
 25 25 4C C5 6B 4A 54 AC F7 0B 5E EE 35 8D F3 9B
 8C B9 36 E7 93 CE F0 D6 41 42 56 09 B9 A2 7B C2
 AA 86 51 96 F2 8E 5B 3F 0A 7D E3 DC 8F 15 E3 D7
 80 89 EE 9C 8C 47 84 31 2B 10 51 51 FC E0 84 92
 8B 84 79 9E 30 84 B2 81 94 F9 3F 2C 0D 33 96 82
 0D 2F 5C 39 8E 8E 27 E3 38 A4 AE 6A 0E 9C ED E0
 23 E6 2C BA C6 3A 36 12 55 9E C9 33 E7 6D 62 67
 04 80 B5 26 5F FD A3 FE 47 8B B8 46 F5 62 EB C1
 C1 CC 48 C3 54 59 96 9B 5A 8F C6 5F D5 DA 1A CB
 AA B2 DB 38 ED CC 6B 2C C6 96 2C 2B 40 6F 0A C3
 F6 A8 CD 33 DD 34 46 D9 23 1C 15 8E 2D AE 9C 8B
 5A DA 70 7E 54 1D 9F 99 01 AF 21 D4 32 88 3A AF
 A4 E8 B2 97 D3 37 99 D7 A5 AB FA EA 5E C8 24 82
 2C D9 66 06 22 1B 0C F9 E1 22 70 B9 92 E4 5F 5F
 F3 53 C4 94 CB E9 23 15 5D 8B 54 0D 6F F9 B8 24
 97 FD 6B E4 66 FA 62 FD 30 C9 63 6A E0 FD BD 1C
 A8 FF F7 28 24 6A 13 49 75 FE 94 5F 2F F1 DA 20
 16 47 6B 43 90 F8 85 93 06 44 7D D6 73 05 A0 98
 AB F0 CF 20 D0 04 8B 05 7D 83 48 88 3C 6E 61 8D
 62 57 E2 83 B6 5A 51 2C E9 D6 FC 2E EE 6B DE 12
 6A FA FD B5 54 BA 8C 11 85 68 4E 5C EB DC F5 5F
 84 25 BA 1E A0 77 7C E3 DB 4D A0 53 A8 19 9A BF
 84 39 65 08 80 B4 C2 0F F5 B9 58 36 2D DE 4C 20
 A7 C0 EE 98 0D 16 9D E0 61 73 29 F7 9C 83 55 DD
 43 7E BA 96 D2 D0 4A 2C 2E 68 9C 9B 45 C5 5B 24
 83 BA C0 EA 83 9F 11 CD FD 38 31 DE 7B 28 C2 8F
 FC 38 34 E4 88 82 CC E0 C8 08 F1 02 B6 21 ED 4C
 FB B8 4E CC B2 68 69 90 14 E9 B2 C4 7E 29 C1 2B
 C5 5C 60 1B F7 1B D7 D2 F7 86 DE DB 0C A8 50 F3
 CF 70 9B 7A 78 45 86 4D 7B 68 A2 D9 42 BE A9 00
 40 C1 5E 65 BE 8C CA 10 F4 47 5F 3D 97 2A 72 AC
 BF 3F 32 87 B1 2D ED 8E 86 AC 7D AB 67 47 90 6D
 98 45 57 3D 42 C2 19 A5 E5 05 41 99 55 C6 6D 2B
 CB 24 20 CE 76 EE 81 E8 31 93 2C EF E9 51 75 24
 10 10 EB 42 BA FB C0 83 82 64 04 FC C8 A1 15 6B
 0F 46 41 AF A5 EB 04 69 D4 D8 DB 36 80 0C 30 AE
 E0 90 E4 BD 23 CC 29 12 BE E2 6B 6B C8 20 F7 11
 DA DF 82 83 DE 02 21 B2 D4 CC B3 61 4B F0 43 3F
 83 63 D1 E3 1F B8 58 31 5F 04 F0 1A DF 4E 69 38
 50 18 A6 2D 40 99 C6 68 75 9B 36 07 9C E9 39 DF
 80 33 FF C5 2C 33 E8 0C 90 0B 49 2D C5 0E A9 01
 FA 86 AF 2D 15 39 61 0C 7A 41 9F 1E B0 AE 24 2D
 AD 3A 1A F3 21 16 C9 1D 3B F7 E9 D5 18 74 90 E5
 ED 94 56 58 D3 40 E3 97 00 78 38 26 7F 2F AC 04
 A0 F9 57 12 71 F7 D4 CA 8D 8E 93 76 79 D7 7C 58
 19 E4 70 36 29 EC 92 AA BD A3 BA 13 7D 1D 8A F3
 CE 28 23 35 A4 50 42 56 8F E9 D0 01 30 F4 E3 07
 00 9E 41 0F 13 49 A2 B8 A5 6C 15 2F 8A DF E0 C6
 56 13 4F 0A BD D7 7D 9C 08 CB B1 D2 A6 40 2F B7
 C0 9F 83 3E C9 AD 6C AC 94 4E 3A CB 1A 98 A0 78
 F7 8C D2 5A 5B D5 C2 05 0D 88 48 C3 7C B3 4D 11
 43 39 E2 2F C9 D0 C2 4A 41 33 B5 A7 1E 4D 63 8A
 BD F9 2A 21 16 96 8E 45 A6 A1 9B 78 5E 4E 5A 68
 01 76 1A E4 CE 30 E2 82 57 FA E0 A5 D5 2B A7 C1
 F1 F2 39 74 0C 22 3C 19 67 A2 89 27 5C DC DA 1D
 0F 46 AF 98 E8 48 72 50 1F D8 5B 1D 67 11 D1 FE
 4B E4 D5 90 90 FB 67 6F 98 C3 19 F1 8F C6 95 74
 43 27 CA D4 30 A9 C8 50 7E 6F 6F 68 D6 1B D7 29
 85 19 79 FE 07 A8 D2 EB 57 36 E4 77 68 E7 00 64
 E0 A7 80 ED 10 B5 37 5B 7A 83 17 FA 40 46 1C 80
 63 A8 5C EA 1F D2 98 69 EE 9E BC 89 88 86 98 9B
 00 DA 51 DD 4D 47 32 E4 34 C8 FD E4 29 FB AD E0
 4F F7 6C 94 46 58 C7 F6 A0 97 87 ED F7 F1 55 16
 B3 59 CE E5 63 B4 7E A3 45 B8 69 1C 93 A0 75 8D
 8E CD 49 E2 8F E6 63 13 3A 8E 28 5A AA 9E 6C F0
 0A 63 82 F3 64 23 9D D2 9A FA E6 65 2D D8 3A A8
 12 2A 55 4E 01 6E E2 45 67 95 BD A1 61 08 4A 15
 E9 09 A3 FC F4 DA A5 EF 3B DD 23 F4 DF 99 09 9F
 A0 B0 15 00 89 1D 3C A6 71 97 CB FE 15 79 EE E7
 65 1A 03 36 2C D5 36 40 0E 97 80 0A 4F A2 80 7E
 53 AB E9 30 E4 79 ED 73 B9 95 D7 E7 24 10 32 E0
 D4 06 76 41 A2 D2 0C D5 16 C0 53 B5 EB 82 79 EC
 5F CC 6A 4E 3B 77 69 A6 5A 4D 43 FC 27 BF CC 62
 D8 0E 08 A4 D2 44 21 DE 62 69 53 B8 0D 70 94 7E
 A0 0C 3E DA 1D 00 51 60 28 A6 D6 E8 3C 56 F6 93
 B0 EF A4 0C 8D 37 98 AF 63 0D EB 53 0C 59 11 5B
 A8 7E 80 9F 43 50 66 05 0E F7 F0 B6 EC 14 64 05
 50 1B 08 04 41 BD 4F 31 7F E1 2B 56 02 AB 1C B9
 FC 58 55 1F F4 B2 12 0A 27 33 4B 4A 59 80 BD 97
 D6 1F 1B F1 87 21 DE DA C3 98 99 24 D1 27 35 9C
 3E F3 C4 1A 1B 1C 9C 62 29 72 E8 02 66 88 14 CE
 20 0B 46 16 8B 21 49 B5 DD 8A E7 8E 26 C5 E4 82
 7C 69 F6 92 9C F3 0C 45 5A 41 C5 02 AA 24 36 C6
 22 BF C9 A6 8C B7 F2 81 79 96 A2 B7 F1 9D 17 96
 E0 7E 52 82 F0 94 63 B7 62 71 8E D0 8C 7C 10 46
 F0 63 44 DA CE C1 EF 4B 8E 78 F5 E1 33 63 3A 32
 E8 C5 50 A1 D5 79 4C 9D 86 27 9B 2E 93 45 27 E1
 4B D6 F3 B7 96 64 4A 44 39 C6 2A 7B AC BE 14 57
 10 33 10 FA 09 0C C7 68 3E 52 6C 7C C6 29 95 C3
 22 B5 68 4F 04 E2 EC 6A 63 D6 75 D5 2D 7F A5 A8
 C2 5F F7 43 B1 98 D0 F9 CC D4 C4 DE 06 36 B0 0F
 AA 43 25 0F C4 8C C4 D4 31 0A 5D A1 0E C8 76 73
 10 4B 80 69 4E A5 68 2C 3A DE 25 44 81 D9 7F 7B
 12 99 EC 15 82 46 8D E4 45 98 AA B7 95 73 96 38
 58 1D F7 69 54 23 75 DF B8 AC 88 06 53 25 DF 90
 04 84 D5 D1 06 31 48 E7 82 C7 25 D3 19 9C 04 97
 76 9A 5D E8 A6 48 5F A9 55 1E 19 19 19 CA B4 1E
 7B 32 57 BC 84 62 5D 8F 22 F6 94 CF 83 16 7A 97
 F7 EA 98 AD 67 AA B3 B6 F4 D7 16 05 89 55 04 AA
 4C AB A3 B5 2B 63 15 CF BB 0F 39 DC 89 01 86 83
 92 86 7E 0A 68 45 8B 03 25 3D D2 33 D8 03 7D 21
 A5 72 E9 CB EA FB 3F DF EE 1E 67 37 3D ED 43 62
 39 BB EB 23 51 D7 6E 58 6B 7C A4 C6 2C 1A 9C 37
 29 A3 B8 33 4E 28 B9 2D 35 F0 2F E6 BB A3 6D 75
 E7 B4 01 AE A3 9E EB B2 B1 BD 4B 1D F4 A8 F0 AF
 7B 2C 8D 91 80 B7 28 36 3E C6 BE 64 7A 3D 21 0C
 B7 3F 53 BC 50 AC A9 7C C4 96 42 DE 88 1A 47 2D
 A9 A7 BF 25 58 0F 61 2B 4C C0 03 4C 43 3A DA CE
 78 BA 40 76 10 F2 C1 58 AC 7E A8 D4 57 D8 3A 05
 87 2E 2D 4F C4 74 5A 88 70 D7 C5 AA 76 03 35 FA
 0C 9F F1 D1 53 52 FE E3 96 90 04 30 02 62 44 5C
 7F AB B4 6C 44 A3 5F AB 8D 90 B8 AD 9C 3B F8 36
 B4 D3 97 9E 70 F2 02 36 47 E5 1B 5B B0 91 BE B5
 2C C2 23 55 A4 A8 20 B5 29 FB 2D 2C 1A 25 ED B4
 44 AE 26 A0 64 23 E2 5B C7 49 3B 08 7D CE 44 F1
 AC F1 73 95 ED 61 2C E7 7E 8E 44 10 72 EB D4 4D
 57 29 77 6E 55 BA AD C6 E2 33 84 E2 A8 E5 25 F4
 53 EB ED 96 A9 8E 00 A8 99 0E E1 39 3A 9B 3D 21
 76 C3 CD 48 BB 7D 52 02 A9 5F 86 95 AC 2B 38 97
 69 64 FB 73 C4 1E 37 84 09 BB CE 1B F1 3F 2A A8
 8A 60 52 E7 12 F4 19 3F AD 11 E1 10 BC 55 4D 1E
 5C 0B 5E 68 FB 2F 83 DE 86 2F 2E B5 98 23 F4 0B
 88 AC AA 47 97 78 A5 4A 86 AF 53 F4 B1 A8 37 3D
 1B BF 13 3D BF 20 DD A9 E7 A2 B4 3C 50 AC 50 AB
 A4 F9 A1 4B BF AB A7 68 1F 04 2D BB 10 58 7E 6F
 EA 7C CF 82 A7 02 1D E3 DF 7A 98 4F 8B 56 C2 30
 AF 00 49 98 7F 25 4F 25 1F 4D DA D0 52 76 F6 DA
 2F 03 B1 8E DF 3F 46 01 47 29 2F 39 B8 B6 42 4B
 79 A4 75 69 E5 F0 10 DF 94 CE E6 AE FC 2A 58 82
 22 A4 E1 CF 67 B0 94 7D 8A CF AC 23 9B 3A E5 DE
 6C 56 E7 CC 2D 5A 65 3D 22 73 69 33 35 A8 5B 06
 59 0B 0D 17 C5 EE 49 5C 9C EB B3 A9 3F 63 A5 44
 45 8E B5 F8 C2 10 00 4D D1 DE F2 10 01 7B 7E BE
 83 E4 02 6C 70 95 0D 32 5D E5 C8 4C B5 DA 30 AF
 19 1F 68 27 8D 85 D4 C2 1C DE D3 59 79 EB 39 9A
 7B 7C DA 78 68 1C BF C3 DD 43 41 1A 97 DD EA 82
 AC AA 3E 84 7E 9D 77 48 E9 17 12 FD 0C 22 CF B7
 5F D5 CB B3 DB 65 50 2E E0 AC 26 5F 08 F7 1E FF
 5D BE 3F CF A6 DB F8 30 01 91 58 7F 2B 2F 8E 67
 70 18 54 85 28 23 9D 0D 0C 3C EE 32 E1 E8 C7 35
 6E E8 6D D0 30 26 48 83 FA D9 FF 2F E4 C4 BC BA
 4C 00 B4 1A 1E 04 10 62 DA BA AC 51 96 EC 92 59
 1F C5 EF 13 6F DD 2E DB AC 73 B0 B5 B7 82 01 2B
 BF 7A 15 D1 CA AB 38 52 EB AE 9C F0 CE CB 7E F9
 2C 41 58 CA D6 23 0E C2 E5 F2 C5 8A 7E 23 EE 9D
 53 92 CA 69 84 F6 2B A5 E4 5D 53 28 40 49 95 FB
 F6 CC 0D 8C 1A D2 4A 2C 39 21 E7 47 25 8E 73 52
 1B F2 96 19 58 ED 1E 9C 04 8A 50 AA 5D C9 52 F1
 04 00 95 73 D9 F0 AC F7 7D 3F 3C F2 54 49 7D 80
 E0 10 23 54 A9 6F DF 12 8B CD B2 C6 95 F2 73 6A
 C8 C6 AE 43 7E 43 98 11 7D 50 9B 0C 78 76 73 7C
 66 35 09 21 06 3D AB 5E 75 2F C6 DB BA 69 6D 89
 83 DA 9F 80 66 C5 D5 EA 3F 84 07 31 85 AD 4B 6E
 98 77 D0 03 01 EE 5D 54 54 41 56 04 FE CA 72 C0
 BA 3F C3 6F 25 C9 48 99 74 63 1E FC 37 CD 8E 2E
 E6 E8 39 B9 90 4B 7C 88 E6 CC FD 3E CD A7 FC 2B
 12 E5 E1 EC 00 E4 B0 6B 03 17 AB 04 51 E6 C9 0F
 58 5F A9 34 E0 92 F1 65 4D 33 15 88 F1 86 4A 16
 8C F1 38 20 52 04 EA 4E 3B FC 48 64 84 BB 05 27
 E8 57 7B 66 7B F8 E6 12 7F B5 A9 AE F4 37 AF A7
 9D 87 FA 11 CD 76 44 19 A6 5A 76 F5 76 04 BA F1
 31 BD ED 1B F9 9A 19 A6 18 B9 B0 3A 0A D5 F6 A8
 9D 98 10 ED E6 FD 28 CA 73 1B 36 85 A9 EA A8 79
 70 82 FD E6 6F 82 EC 4A 08 3D BB 5E 01 7F 28 15
 69 13 43 05 16 D6 9A 1C 7E 02 5B 33 82 A7 BA 02
 01 A6 C4 F8 16 24 CD 50 87 49 4A 6E 5C 6F AB 4F
 20 F9 21 C1 B3 43 A9 BC 40 5F 8F 24 BC 3B EC A3
 01 3B 02 14 4D 1A C8 F1 8B 59 D9 28 1C E4 95 68
 10 97 88 A2 90 3E 50 B7 DF C7 6E 6B C8 06 4A 04
 74 FD 8B EA 1B 16 EE 7C 47 D0 B0 6E 35 57 E5 37
 78 64 CF C5 11 6B 71 EB 3B 68 11 E1 E9 BC 68 98
 95 4A 50 33 9D A6 39 77 FF 31 9B 71 B3 32 57 6C
 CD 22 80 2A EE CA EA 75 E6 ED EE 1F 6F 77 AC A2
 0D 24 40 FB 60 99 05 D9 63 75 8B 87 7D 3C C6 82
 E2 76 4C 28 80 0C 9A 39 CB AE 32 1D DD 7C E7 A3
 B8 AB A6 6D CA 62 85 A8 4C AA 1E B2 43 61 99 3C
 12 05 BA 52 78 72 23 DD E2 1C BF 95 68 49 C6 17
 55 B8 3C 7C 9C 26 DC B6 9B 4A 32 76 57 5B CB C0
 0F F8 2D 23 04 14 B9 BE 66 AF B8 09 29 33 7F 04
 9E 2B 68 D2 02 42 2A 9D C4 15 18 59 FF 55 DA B4
 8C 28 E8 69 4F B5 BA E6 F7 71 10 23 1A 5F 7D 19
 79 8B A4 71 8B B2 56 11 5E 61 D0 C0 20 F4 22 AA
 E2 EA 7F 9D 38 4F 2F F2 AF 07 E2 EB 20 74 24 C5
 23 53 CD EE B6 2C 8F 59 97 69 EC DC F4 C1 C1 26
 BB 61 D3 FD 94 19 EC 9B CC 32 0D DF 3A DD 4C D4
 8D 54 9E E0 EC 5E DF 4A 92 93 95 87 52 9E AC 52
 78 07 1A 00 ED 72 75 C1 96 66 E2 54 91 A9 B8 5F
 6C 7B C9 AC D2 59 CC AE A2 E7 A2 C5 FE B4 FD 36
 BD DA FD B5 9A 95 4C BF 8A C4 06 D1 7C 4A 62 6A
 5F A3 1C 6C E8 24 32 C2 46 D0 FF EE 34 6A DB C4
 5F E8 26 68 0E 6A 47 19 36 04 93 16 ED F1 B3 22
 4A 3D FA 22 B7 B5 E7 A7 C8 4F FB 7C 7F 6A B6 0D
 1C AE 93 05 89 C7 DB 3A A7 6E 94 52 4C E4 D0 D8
 CB E2 D2 73 AD 1C 68 3A 4D 92 90 A6 66 3D DB C6
 FD 9E B7 CE 30 D9 9D A1 AB 40 4D BC 31 A2 96 F8
 0C 46 67 8B 70 78 1D 33 43 A3 7A 19 38 05 CC 41
 CB 8A 6D 88 AC 9C CB C5 F4 70 38 A3 A2 E1 D4 64
 60 34 FD 54 3D 65 63 43 35 7A 4C E6 B3 D4 55 03
 2A 01 81 1F 24 9D C8 99 D5 F4 55 81 8E 47 0C 2A
 BA FC 77 D3 03 C5 27 6E A5 22 AC F8 FB 15 A6 9F
 42 07 B4 07 F9 B3 30 37 66 D1 28 1D 32 CA 7F 8D
 43 F1 66 FF 79 51 3D E2 F4 2E C9 4E 2E 4F 72 03
 73 BE 4B CD 11 A2 90 E3 E2 AA 77 69 C7 6F 33 FE
 D1 E8 3F 0F CE 66 5B 20 4E B3 B6 58 D3 42 04 1D
 25 2E 4E 38 EF 9D 5A BC A8 3C 49 46 B2 45 7E 81
 C2 B7 63 EB DA 63 55 94 51 68 77 18 95 89 0D 81
 0B 3F 8B 79 EF 61 6B AF 50 EF 70 E6 5F C0 27 6C
 1D 42 D4 E8 7A 97 0B 2E 53 C8 F3 55 10 1D 51 46
 D0 FC 37 B7 85 AE 58 1B CD 2D 82 BF AE 1E F2 44
 3A 8E D8 E4 5A ED E8 65 4D 64 20 D9 B8 DC E4 C9
 3C 31 BD 00 EF 9F 7B 38 61 3F 8D 5D 21 D5 33 EB
 8E 36 F2 19 21 10 04 6D 05 74 24 72 A6 21 55 B3
 8A D6 EC 12 56 C1 8A 3C 3C 7E 1B D8 36 0E 20 EB
 A7 22 C7 36 A1 E6 E6 AC DB 35 8E 68 24 1E 93 FC
 0E 6E 2E C7 8E 96 AB 8B 5A FE 98 9E 7A 46 65 21
 C8 07 82 66 46 C0 21 7D 42 0C 82 79 38 F5 CB 1A
 C3 64 68 DE DF 44 CB 49 FE D9 CD 75 5A 97 DA C9
 2F A0 D5 16 66 EF 79 D8 1B 6C 88 57 A2 73 C6 41
 FF B4 91 F7 E5 B0 0E 92 E9 2F 70 76 EA C1 77 92
 B4 48 65 FB F2 DC 42 79 DC B1 0A E6 2F 1C C4 96
 34 80 28 26 0A FA 28 ED D7 99 C7 36 3B F8 DB 8D
 F9 A3 4E F5 F9 6F 02 3C 33 FD C3 4A 9B 5B 3C 64
 7A 9E A1 D4 44 95 2D 2C 17 19 D4 E9 A4 31 0D CA
 D1 24 55 C2 AA C1 B2 40 FE 21 D7 B6 B1 8C D0 66
 6D 3B 2A 0F 42 5F 3D E9 3F 47 3E 4E C1 35 70 89
 87 93 E0 9C 34 1F 6B 60 EF 7F 8B 66 53 22 C7 53
 46 B0 88 C3 B0 04 E4 96 BC 07 A2 80 A7 62 7C F0
 AF 67 BB 6E 76 98 66 D7 E5 A6 33 07 D5 D4 CB C3
 D7 F4 F8 E9 DB A2 93 70 D0 F5 91 17 B7 C7 52 AD
 61 94 0E F4 2D 69 DF B6 88 13 E7 FD 6E D2 BC D8
 DD A7 23 DE 07 85 7A 1F CB 19 77 4D 60 45 38 52
 CE B0 AF FD 04 4F A6 56 B6 69 57 C8 61 E7 A0 AF
 9B 1B B6 18 33 3E 22 91 95 E6 78 5A 94 94 8E 02
 F1 93 91 B2 8C 29 52 2B EB 88 5B 8D EC CF BC E4
 5E DF E8 D9 1E 8E B2 F7 AE D7 9C 1E 2E 29 87 CC
 B6 EC 9E 40 5A 82 25 58 84 D9 AC FF A8 59 52 76
 6B 75 21 49 DF 2E 03 98 46 95 2E 6A CD 12 1A D3
 31 9A A5 0D B9 E6 E9 7D 9F 83 1A 92 0E 79 B1 7C
 DE 63 EA 18 96 BC 82 A8 77 34 11 CF 65 A7 BB 12
 1D 41 02 C9 BE DD 4F 58 F0 9F 3E EB CE CF F8 B0
 09 8B AB 3D E2 17 B4 37 71 35 41 59 D8 4B 69 07
 AA A7 11 2C F9 A9 6E A6 BC 1B A2 D2 AC E7 DD 61
 6F AE 3A 97 89 AB 38 5A 37 80 14 C9 7F 4B CD 00
 C9 BA DF CB 77 A4 99 97 1F B5 AC F9 CF F2 95 52
 96 D6 7D 55 89 CA 14 D8 F7 7E D7 14 45 A6 9B 3C
 2B 56 04 52 29 0E F0 48 D1 5E 1C C0 C4 37 1C 96
 CD AF F0 F7 76 DA 76 8E E2 E5 23 23 4C A7 DA A1
 F7 16 87 D1 5F F7 DE AB 56 5A 31 2D AF 13 2D 4A
 96 88 10 C7 BD 8B 18 C2 E3 A2 DA 8C B7 90 BA 18
 92 BF 1D 8F 28 58 27 5B 71 A0 3B 4A 89 A7 90 7F
 BA 26 CB 9E 05 49 A2 3F CD 82 BC D8 0D 9A 3C 52
 45 33 F5 9C 9D 7B 1A 8C C5 C3 DC 44 96 1A 5C 6D
 05 BC 79 9E 32 BB 37 0B ED AB C6 BF 07 64 5C 86
 17 DE 1B 46 74 E8 39 D3 26 E6 99 29 B2 B6 FA 38
 2B 64 C6 70 9C 62 60 4D D4 00 2C 76 D1 4D B1 8A
 FE D3 30 DC E3 2B 24 9B 09 26 C5 50 15 69 83 D9
 72 01 2F DA 99 B8 89 C0 97 E7 D4 9B BB 31 03 60
 AE 10 E4 F2 1D DE 76 DD 20 C3 D5 DE F0 A9 CB 04
 2E B4 FE 0C F4 08 D1 61 40 5D F3 D0 8D 9F AD 7E
 DD 4C E6 35 57 8E 04 60 F5 52 51 BF 36 F0 1B B8
 FA 52 50 4E 45 4B 2A D8 E9 C5 D0 48 AE 65 26 C4
 B3 92 D4 3F A5 CC 0C 69 40 5B 6C 18 0B 26 B4 67
 03 6B 6A 26 44 FA F9 39 A3 19 ED E5 4D 1C F5 C3
 CE 76 BE EE A0 EF 89 A9 A1 C3 84 31 EE B0 2E 48
 14 74 EC A9 F4 AF 88 A7 15 AA B0 62 64 C3 8F A9
 49 E1 91 7C 9D 01 FC BD 63 78 16 40 94 0F 9E FA
 61 32 E0 09 34 D5 F8 C3 8B 18 6F AA 8D 52 74 88
 B0 33 EC FB 21 99 75 C6 FF 40 12 B0 A7 D0 77 C3
 CC 00 46 9C A5 76 6B 80 76 60 A5 82 9E E9 C2 A1
 6F 93 98 B3 67 2B 96 10 50 F9 FA F8 27 6E 62 2D
 76 D1 52 3A 27 AE 16 99 A5 E4 FF 5A ED B5 B0 57
 60 A0 E9 21 A8 83 8F 93 3B 0E E7 09 95 49 41 FF
 D7 D7 49 AD 17 41 AE 5F 19 50 07 27 83 7E DD 5F
 E8 8F 56 04 3E 6F 1F D9 6D 3B 60 28 EA 24 D4 AF
 27 4B 56 05 F6 F1 44 AD 2E E6 AD DF 88 B0 09 A6
 79 50 E2 54 29 89 69 93 B9 E2 CB 5D 87 92 C4 73
 EE 78 51 B8 CE 7E 21 E3 BD 9F C1 3E AE E6 95 B1
 94 02 CE EB 10 DA F0 4E A6 F0 71 BB 38 6A 1A 3A
 15 7A 14 05 5C 18 24 60 DB EA DE 47 9D 16 B5 59
 D7 2B 33 63 D4 2A 80 C0 1B 87 82 54 A7 BC 04 EE
 FD A8 21 B4 E9 57 F1 56 F1 79 C9 04 C8 07 66 93
 9E 1A B3 A9 78 C0 28 52 C5 1A A1 C4 AE C1 BE 3C
 69 04 9E 9E 15 67 14 18 B7 4D 8D 33 79 AF 4A 22
 E8 D6 F2 6B 26 45 4F D0 BD 0A F5 5D A6 A6 65 00
 7F E6 39 1A 58 0D 33 30 6A 71 F4 EC 57 5D 31 AC
 2B D9 21 39 BD B7 64 ED 7A 0E FF E3 E7 60 7A 16
 08 3A 22 BD D3 2F 07 71 3B 77 2F 5C 4E 3E D2 54
 67 05 CF A1 19 47 9D 1C D2 E0 BF 35 A5 F5 68 60
 D5 01 40 DF DF 10 F8 35 FA 0F A3 3B 9F 6B 91 36
 E2 A4 99 04 D3 B9 59 A4 DB 9E 83 21 75 45 6F 67
 89 39 AC BB 29 A4 B0 EC 07 FB 3D 1F 3F C1 35 6D
 CA 26 13 D6 B3 4D 49 DA 0F F3 08 7D 20 BD 4E DB
 C0 3A 20 50 BA AD E8 F3 F9 36 2B 73 BD 17 55 7D
 43 C1 2D E4 B9 8E 07 FA A6 E5 81 FB A5 D7 3D 1D
 5B A9 30 46 9E D5 30 6C 22 03 A4 BD 33 BF D2 C6
 92 DB 6B EB B7 B6 0B EF 86 25 C9 1B 9F F1 0A F0
 C7 37 92 EF 2F 58 E4 52 BE CE 3E 3B 1A 4E 9D 83
 63 D1 3B 3E C9 93 74 67 F4 7F 54 23 90 06 2D 87
 F0 77 FB CB 5D 03 7A BC FB 5C E8 4F 88 9A E6 93
 BE 66 23 07 2D BD 77 24 C7 61 21 8C 69 3A 49 81
 1D 9C D5 E0 8A 82 24 05 6B 31 EE 83 0E E3 80 42
 72 75 D6 FD 31 CC 83 7E E7 54 2C A4 3F C4 E6 0B
 1C 3D C8 3A 4C B3 54 A9 85 1F D7 E7 B5 44 17 21
 96 34 F3 61 CE 36 A6 53 9E 87 89 73 70 F7 AD 3F
 E2 B2 92 58 A9 F0 EE 25 55 08 D6 DF 9B 9F 97 9E
 55 A7 3D 4D 5B 5E DF D7 AF 1D 8F 2B 97 5E F8 C5
 5F 38 64 EB 71 6F B3 B7 80 4D ED BD BF C5 0A F2
 B6 A4 08 DC C4 20 77 CC 59 96 05 88 C6 9B B4 F2
 81 4C FA 5B 7C 4A 16 7E 9E B5 1D 50 81 1F AA 4B
 B8 55 1C B1 67 60 19 0F E4 3F 75 2D 6B 0B 35 61
 91 A9 1D D0 5C 3E 71 EF F7 BF ED 75 71 09 87 05
 09 33 FC D0 B7 AE 39 CC 4D 85 B2 B9 06 E3 E1 5B
 8B 16 5F 9A 7C CE EC 9D D7 22 4B 05 F2 C6 61 65
 70 04 B9 2D 22 43 C1 17 E9 73 72 4F C9 97 F7 F6
 4C FC A3 DC EA 03 E1 11 B6 BB FA 9E 12 FB 59 D7
 B1 D8 82 F0 9A 0A CE 09 29 35 46 CF D9 FB C7 CC
 02 7B D8 C7 A5 64 A9 CC 0D F8 BC 41 8A 53 A4 11
 67 AD B9 5C DB C5 C2 7E BE F0 75 01 4F 6A FA F7
 02 E2 12 DC 20 F4 62 D8 A0 A9 BE 45 1D C2 66 E2
 8B 27 64 25 D8 E4 4E F2 10 A9 4C EB 7C 60 BC 09
 9A EC 56 30 41 C1 D4 14 21 66 98 1D 07 E9 AC 46
 43 5B 4D 91 A3 D4 69 38 C7 B4 87 A3 67 30 4D 36
 85 C9 57 85 51 F3 9E 62 26 07 A9 91 A2 4C D4 16
 5C 2F BA 09 CC ED 54 4C 4D 06 CD DA D8 FF 90 61
 9A 47 3C C2 E2 22 58 9B 49 AE 0D 7C 0B 5A 50 5D
 AD 77 2F C4 2E 09 F4 E3 19 58 32 C3 5D 90 C3 9B
 A2 CF 09 BA D2 22 47 1C 4B D4 F4 50 21 D4 13 EE
 A2 B2 AB 08 7A 66 40 44 1B F7 56 CA A7 31 01 B7
 1D 38 CD 62 38 A6 0A 37 AD AB 15 4A A9 2E A3 04
 4D 80 D6 39 4D 14 1D 6D 27 0B CF 5B 7D 08 ED 44
 B7 F4 DF B3 4D E9 D6 BF 36 99 B7 DC 9C C4 D1 F5
 35 F6 A8 53 0D 7B 53 EC 28 D9 64 2E 47 74 AC F7
 E7 6C 52 F9 35 F8 7B 97 7C 53 7D 66 22 74 FC 23
 6E 75 E6 9F 62 36 27 AD 19 CE E5 00 BB F3 CE 15
 E6 FC 74 D7 8D 4F 54 7A 54 F6 AB 42 8A 42 2D 2F
 46 BD 1F 2A D9 32 17 16 6A A5 63 06 D1 A9 0C 82
 81 B9 19 08 A4 D1 5A 59 52 BF 6B 8E 92 68 C9 50
 1F F5 02 6F 8E 67 FD 57 BB 73 1E 5A 3D 21 40 4F
 E7 89 56 0A A0 7B 63 2A 53 A1 7A 27 7C BF EA E8
 4F CE 77 4E F3 0A FA 8E E2 E7 23 30 AF D8 12 12
 AB E7 CE 05 17 04 79 D1 89 1E 85 DB 6C E2 DD AB
 EC F0 79 FB EB 79 DE 3C 2D 3B 1E 2F 33 6E 9E 7B
 8E 05 D4 BE 1B E0 D3 76 23 A5 C4 F0 91 E4 33 82
 FD 25 07 6B F7 3A 3C 98 EA CC 2C CB 9C 07 D3 82
 FA 7D 42 3F E6 22 19 43 95 B0 3B B9 BC 62 06 A8
 D0 B7 BC CB B8 C7 4F DC A6 18 CD 9A 43 6A 56 1D
 E3 F1 8D BE E4 6C 2D 55 7F 83 85 C6 41 92 26 11
 56 40 F6 E7 DA CD E3 34 FE EC 79 10 BE B6 C4 25
 AF 10 18 74 17 72 54 52 4D F5 F8 1D 29 10 98 BF
 7A 2B 9C 01 39 B3 51 9B 62 A2 59 BC F6 16 EA AE
 8D 6F 81 F1 1F 95 30 49 C5 F3 EB 15 FE F6 DF 2B
 44 A6 4F C1 E0 8B 73 D7 25 9C D6 13 8B 19 CF 85
 58 97 D6 3D 46 90 09 EA FF 13 F5 77 36 0D 10 F6
 8F 88 DC 0C 15 6C E7 E1 EF 58 29 71 D9 5B DF B5
 AA 32 81 3E D7 7E 41 03 A3 CB 68 DD 60 4F A0 46
 12 C4 F1 2C FA 02 D8 95 CE 78 D7 CE 27 26 1A F3
 AA BA C6 EB 4E D8 08 D4 3F 94 4C 56 6A 05 5C 9B
 BC 27 17 25 23 D7 8A E0 CB BC C2 D1 71 89 BE 75
 B5 19 74 A8 43 22 62 07 DF 82 3E C5 51 92 DB EB
 91 A1 9C 77 CA B1 AC 77 BC D0 E0 AE D3 64 A6 86
 CB 6C E3 A0 4B 8A 5A 69 A9 9F BE 96 79 3A C0 51
 90 8C 2A 2A 1E 3A F4 DB 38 39 4B 70 76 6D B8 59
 C2 78 C9 C1 E7 AB 68 D6 81 93 B3 C8 27 42 7A 4C
 CD 8B D2 DA C8 9A E8 14 AD 85 31 D6 BE 69 64 3E
 9A 61 EB DB 22 A5 DA FA 94 A8 7D 57 65 16 A8 1B
 48 9A 5F 27 B0 6D FB BE C2 C5 65 82 C3 94 20 FA
 3E C3 88 31 BF A6 3E C9 18 31 8E 2E 7A 80 DC 08
 36 67 D4 02 14 FC 86 56 D0 3D DA 9F 0C E8 DD 7D
 56 FD BE 90 59 D7 1A F0 DA 70 B6 DD 12 55 7F 20
 F2 FA F9 A0 1B E1 FF AD FC EF 70 83 98 16 50 86
 FF 52 47 05 E3 58 B9 C4 B3 D4 7E EA CD 21 08 1B
 70 9C 2D 49 6C D4 E9 A7 97 97 F4 28 14 78 1A D8
 CE 46 CF 37 30 41 53 08 3E 57 D5 76 EC E6 2C FA
 F6 36 C2 E7 69 41 1C D9 22 E2 51 58 40 2A 9C 0C
 B6 09 80 C9 E4 33 00 58 9B 3B 4E DA FA 1B BF 0A
 C8 33 31 11 94 70 E3 5C 5A A9 4D 1E 9B B1 01 8F
 7E 1C E4 B5 F6 86 BC AA 13 55 A9 33 A0 85 99 CB
 CF B8 61 F7 8C 42 19 F2 86 01 E7 02 EC 78 75 D4
 E1 D8 B1 CB 15 79 5F 07 3B 9C FD F5 13 1C EE 82
 BF AD 84 DE CD 03 1E 20 85 64 A4 E5 A6 24 D8 B4
 8C BE 12 2D E1 E7 8F C2 7D 51 FB 9B 51 62 9C 70
 B0 0C EF 13 01 41 E1 2A 1C 38 53 B5 22 6C 10 81
 F9 99 FC 23 F6 20 2A E0 F0 D7 B7 3C 7B AA 8C 5C
 C4 3E 02 96 30 DA 9F A3 CB 78 76 EC 8C 66 60 89
 E6 B0 53 70 A3 41 2E 03 35 21 3C E4 4C B1 B6 FE
 F7 8A 0B 2C 0E F1 17 FE F9 B5 D3 C4 FE FF 06 BE
 37 97 3B 8F 57 C3 C4 9A 46 98 81 76 17 15 0C 86
 6E FA 12 9B 8D D0 9C 05 AB DA 70 33 11 E6 38 C4
 BD 05 98 39 8B D2 39 38 B0 8E 36 12 8E 54 11 90
 30 AE B1 16 E8 E3 D3 5B 4F 98 FA BE 47 A8 17 5A
 2F 46 42 69 90 87 0A AD 4D F1 74 9A 1F 80 C4 93
 57 17 3E 9E 86 C8 B3 78 6D F1 2D 22 27 BD AA B6
 30 72 F3 7C 79 33 82 1E FF 3A 0F 42 35 4E 05 03
 82 76 B6 2F 15 A8 B5 4E DB 8D B4 D8 12 6B E9 03
 E8 E9 EE C7 46 D0 88 4D B6 53 8E 3E 82 69 57 10
 73 23 44 B1 AD 4B CA 76 D1 91 D7 5F F5 1E 95 5B
 96 6E 8F F6 CA 30 57 F1 3C 91 86 74 9F CF 9A F4
 E0 20 40 0A D7 1B F6 79 D7 B1 7E 2B AE E5 0E B5
 56 34 8E 1F 62 21 A8 1A 4E 9B 90 39 E7 E2 3F 83
 E0 29 82 D5 0F 82 B0 5A D5 6E 55 3E DF 2C 26 BC
 37 DE 16 0D 2F 4B DD C3 10 24 F9 83 34 FD C3 BF
 B6 2B 1C BC 36 06 DD B6 B5 67 3B 0C D7 E8 BF C7
 08 8F 2B EB E4 83 19 C5 FD EE DC F6 C9 06 75 7E
 D9 C7 B6 1A 61 C9 1E B7 57 C0 98 DB DE 91 6A 0C
 90 83 B1 52 FC 38 0D 0D 26 2B 65 23 C6 92 78 92
 8D DF C1 D9 02 49 CB 99 5D 70 21 B1 1D 5D 91 71
 98 B2 3E 4F 47 F0 E6 2F B8 A0 90 4E D8 08 59 26
 51 75 7A FA 59 7F FE 9F 8F B3 F5 3E 4E 4C A7 CD
 80 CD 76 E1 1B 3D 28 C4 3D 65 7A 23 34 56 DB E5
 30 AF A8 01 4A 95 AC 71 1B 4B 47 77 7F 41 84 E2
 7B FC 19 4A 4C 2D BB 55 C3 CA 61 EB 22 BC 93 4D
 86 92 D7 0A 47 6C B7 27 4B C8 2D 19 9D 37 25 E5
 9F 04 A3 59 EF E8 11 58 54 D7 E0 DD 21 B1 36 83
 AF AA 70 B5 A8 50 8C A7 78 8C 19 2B 3B 9E 6C 2B
 BD CF 36 63 F3 AB 1B 4B 76 CE 90 E9 F4 4F D0 0C
 78 77 77 ED 9E BB F3 A1 42 71 C7 4D 55 0A 54 AB
 71 0F BE A3 3D AD C2 84 07 45 00 7C 18 50 48 C9
 4C AE 12 25 E8 93 01 6C C1 3E 89 34 01 78 56 79
 3E CB 70 E0 5E 30 6E 2D F5 E3 13 14 95 07 35 6A
 5A 79 17 46 1F F6 CD F2 62 17 6A E3 70 2C 54 A7
 95 5E 8A DB DE FF 8D 43 BE C8 BA B7 F1 16 08 39
 09 0D 18 73 37 24 30 02 0A 35 A5 7A 52 27 0B 57
 DC 6A 1F EE 17 98 C1 DD 81 93 94 ED 7E 5C 79 64
 6F 65 1A 6D 9F CC 5A A3 A1 DE E1 18 C4 77 75 17
 16 6F B1 64 9E BD 29 F3 C2 3C 75 BE 54 5C 97 47
 0A 4B 2A 16 BF CF 79 FB 64 11 F7 22 F5 4F 73 EB
 D1 6F 3C 58 6E F8 B1 61 E2 59 4C 74 05 C0 F3 49
 D0 D7 28 10 60 BE AA DC F2 7B 51 83 93 54 E8 4A
 09 8A 51 1E A5 D5 5F 53 B8 25 5E 17 DD D1 93 98
 97 F6 B5 75 07 1D 8D E3 D0 20 6F 8F 5A 25 F9 CD
 D2 06 AA 70 44 D4 43 A0 C4 E4 91 A9 AB B6 AB 29
 90 D1 42 21 8A 60 31 CC E3 7F 7F 42 18 48 AA B2
 06 C3 3E 72 6A 5E BA 30 E0 42 97 CD 61 70 3F A0
 62 FA 7E 88 90 52 38 CA FC 9B 8B FB 14 06 4E 6B
 6F 30 79 C0 9B 58 0F 89 DA D7 E3 4D 6D 79 EB AB
 09 67 70 C1 1B 2D 33 2E C2 41 40 C3 DC AD 4E E8
 24 68 DD 43 68 1E B8 F6 37 EA D3 8D 4D 72 25 24
 DC DD 0F DE 4F 83 E3 27 26 AF 34 15 A6 84 40 96
 48 23 75 33 76 1D 0C E6 ED AC 7E DF 39 D6 3F A1
 5A F6 D5 B6 13 13 46 85 63 41 B0 9E B8 89 07 34
 CB 0D 3B 75 93 EF 19 EE E8 F9 33 8C C3 D9 54 D0
 6D 72 1C 0B 3C 86 9C A0 B4 2C AD E6 11 EB B0 13
 3C 7D 56 21 76 BE F3 FF 5F 2C 6D 08 49 4E 91 79
 03 ED 6E 1E C2 9A 5A 7F 24 F8 AF 85 B4 33 AB 7F
 09 C2 4B 4F A4 CF AD 7F 03 A6 62 41 87 33 08 8A
 02 BB 74 8A 7C 76 97 40 73 34 13 66 35 E9 F5 34
 56 94 DC EC 75 9F 79 05 9D E4 CF A4 7C B2 92 9B
 4B 2C CD 1E 8F F5 22 91 E6 D0 E7 5F 5C D6 8C 79
 7D 0D 57 B5 4B 6D C3 31 0B 8E 8C 26 D1 6E 0D A8
 28 72 CA D5 83 B5 CA 19 E0 33 D8 0E BA 4D C1 CD
 B9 50 45 03 63 99 7F C3 38 46 A3 8A 0B 99 0D E6
 9F 9B DF 92 C4 B2 D6 18 6F 52 9B E6 27 4D 64 88
 65 D1 4F A2 5A 1B CE 5A B9 B6 13 0C 17 D7 B9 61
 CF F0 B5 30 BE 6C 39 E0 BD FD 61 38 50 5B F9 8A
 91 E9 D3 CE B9 DF 0D 4C C5 DF 6F 8D CA B4 DC AC
 F3 65 A3 0A 98 31 BC 78 84 FA B2 9C 36 13 EC F8
 A1 83 62 A9 C3 D3 86 2A 6D A3 FE 58 76 E8 4C 12
 CD 1F 74 92 86 4D 60 69 D8 26 D0 30 A1 7B 63 0A
 B9 82 0C 65 8C 8F 3B 10 A8 47 7C B5 44 3F A8 80
 1D CA EE 14 D3 BB 08 C2 56 2D 7A 6B CC F1 C6 25
 38 13 C8 13 53 2A 9C 38 D5 20 AE 44 94 80 81 9E
 34 50 4A F3 0A 82 C1 B7 90 49 1E 61 5D 76 C8 73
 72 5D 71 27 23 A9 EF 7C 47 CF D7 89 C6 B8 05 6F
 00 88 64 56 BE 3E 4A F5 5E 80 FF 28 AA F0 B2 60
 A8 56 FA 4F B3 01 58 17 57 E6 B0 3D 52 73 93 E7
 CB 15 09 FF 50 29 32 E6 3F EB 4F 75 99 7F 05 4F
 EC 47 80 AD 9B 8E E5 6F 62 E0 F4 34 6B 87 FD 29
 A5 DA 3B BE 67 8D 61 EF 52 75 FF 57 48 8B D3 35
 9F 1C 11 C5 D7 11 98 1C 73 C2 09 66 7C B0 15 D3
 0F 8D 1B 54 00 D7 09 33 A4 3B EA 0B B7 45 AF A9
 00 EB F7 CE BB 36 F6 04 1D 67 FD DD 08 9E 1C 65
 B1 F6 AE AB CE 3C 5F DF DD DA 84 B7 6A 64 08 B3
 6D F4 2D 14 7D E8 86 FD 9A 0B 5A A2 61 74 B1 79
 8B 14 A4 68 8E 61 B5 E8 CA DC AD 58 07 21 23 4F
 21 08 A3 55 8C A2 F4 C6 08 99 3F 22 1C 71 1C 27
 EC A2 58 AC DF BA B8 C3 B4 3B E5 8D C1 C3 42 BC
 75 78 88 68 51 A5 1D 9B 1B 19 95 57 52 1C A4 4B
 75 AE 63 59 30 66 C3 42 5C 17 B7 AC 0A D5 6A 35
 4F 97 C5 7F 7E 72 17 9E C6 71 16 36 13 A3 6F 81
 07 4E FA DF B8 48 6D 07 A2 63 04 1B 80 CA 2C 8D
 11 D4 7A FB C8 5B 25 97 1C CE 1F 96 7C D7 37 DC
 0D D0 C6 08 0F CD 4E C0 9F AF 00 92 9B A6 1C F5
 A8 7C 56 87 FB 30 9B DD AE 57 9E 9D AA 15 95 95
 82 3F 17 1D 79 D6 9F 4A 74 42 44 4B CF D8 B9 39
 F7 14 A8 7C 20 AF CA 95 87 3F 03 E3 3C 28 2C 78
 7E 5E C3 4D 7B 33 92 0E C1 9F 7E C2 6A EC 58 D4
 CB FC 68 75 85 39 CD C1 7C 33 1A 32 19 37 C7 5B
 7A 37 83 7D 05 67 F9 94 24 86 07 F6 54 33 3D 78
 A9 57 4E 02 07 C4 30 8E BC DC A1 9E E5 7A B4 70
 C8 91 7F 36 76 7F FE E0 A3 EB 51 A6 D7 55 DF C5
 3F 1B 25 AC 78 23 21 14 7B 97 BB FC FC 2E C8 9C
 3F 97 8A C5 D2 C9 B1 FF 26 27 84 E3 15 56 25 AA
 51 61 4E 2B EC 32 70 86 AB 5F B6 BA 75 A5 39 2D
 5A 5E D4 6F BD CE 03 14 0C 96 86 8D 06 8C 8D 41
 0A AD 95 5E 89 4F 62 1D 0D 65 CE F6 C4 21 F6 BD
 70 C6 32 84 C5 DD 20 38 35 34 6F B0 D4 35 A0 22
 0D 23 9E BB D2 78 06 2C C3 45 8D 8D 94 08 64 8F
 D6 12 96 22 4F 4F B0 46 4C 03 85 21 43 4B A6 EE
 E3 87 4B 1E CD 5D D8 16 60 FB E5 BB E1 E9 73 DF
 FE E0 F3 F3 84 CC 43 A6 5E 6A F8 02 C6 9C EC D4
 26 91 B8 A0 B8 C6 AF AB 6A 5B BA 95 95 CC 92 81
 E1 06 8E BD 43 36 27 C8 42 F4 53 C6 F1 41 4D A5
 C9 97 24 EE 28 A4 F6 B4 31 23 E8 F6 76 B7 84 CD
 49 DA 57 E7 80 15 03 F5 D7 D0 7E 5A BB 05 CD 7E
 2A 17 D4 76 B3 CD 2C E0 7F BE FF 15 15 70 59 1A
 43 32 DF 2F 21 A8 AB 00 2B DE 20 C8 D6 5F A2 91
 6C 53 2E 25 21 C7 43 F0 B1 B5 AA F1 D5 FE 7F C6
 F8 28 8A FF 15 E2 EA 71 77 80 C4 5F 0B AB 60 55
 FA D2 C5 10 64 9D 63 74 AA E3 DE 47 F0 D4 AC BD
 3C 12 85 DE CF C4 8F 75 CC 51 20 B1 72 61 AC 6F
 90 78 43 8A E7 FE CE 13 E7 53 36 07 1A BB B8 92
 A2 9F D9 67 1C 86 F2 52 61 CF AD F1 91 89 D4 AC
 7E D3 D8 D7 9F ED 67 C5 C5 B5 F0 B1 F3 B1 52 F8
 7A 6E E0 C6 1D 65 B5 BD CF 2B 6B C3 25 F2 E7 57
 8E 17 3C CB 8E 59 2F FD 9B 08 70 A8 5C AC 52 F9
 F3 CC C8 C9 98 DA B6 40 11 74 81 2C F3 70 98 14
 D1 79 D6 15 B0 DC 6B 6A 20 6F 5F 64 29 8B FC 38
 33 A9 71 EE 12 0F E3 CF BE A8 EF 9E 02 DF FC 4C
 7E EC A9 94 BB CD 27 CF 1D 99 02 33 68 1F F0 63
 A2 C2 D1 77 A0 C1 39 F6 56 34 32 F4 62 EA AA DF
 09 1A 69 A4 08 13 A4 38 C7 CA 3D 97 8C AA 17 6D
 25 AD 7C 4A 25 9B 59 24 75 CE 41 6A AE 54 44 74
 70 FE FC 54 CD F1 68 EB E0 AD AA C1 AD 4B E2 65
 D2 B6 17 A5 2A 10 5B 15 47 BC 75 24 7E 37 60 13
 64 11 37 96 14 F1 68 43 25 E2 E8 55 4D DF 7A 8F
 0C 58 9D 9C 54 97 FE C9 0D 8C 45 D3 4F D0 3B A1
 16 79 96 3C E6 E0 AC F2 FB 45 4D CE 01 7A BB C6
 82 0E 91 E3 B4 68 9B 35 F0 1E 8F 0A DF 52 80 14
 CA 0A E2 1D AA 07 09 12 94 20 3F 72 C2 F0 0A 9E
 77 01 34 86 F8 A3 FB 0B 3F E8 9F C1 67 11 58 D4
 DE A6 EF 69 FF 4B B8 C1 4C 5E 0F 4F A2 EA BA 38
 01 F4 CD F6 B9 0E DD B8 56 BA 21 70 D1 CD 46 72
 9F 94 4B B2 76 F6 FB 9D 8E D0 0F 46 55 92 DC A3
 11 62 36 1F E5 BD 73 32 5C 1E 02 70 C4 E1 D4 E8
 35 14 95 9F 94 F8 30 28 68 C6 68 38 80 24 ED 5E
 54 CD EF 6B F1 17 86 A4 76 54 38 94 33 23 FE EE
 10 8A 4C 71 EF CB AE 0B 60 69 FA 07 C9 94 2C 9E
 2A 6D 89 EA 36 45 6D F8 0C 17 9F EA 14 24 C8 21
 66 F3 37 9B 82 16 B5 8C 99 A6 72 4B 2D 3B E5 F0
 A7 49 E6 39 03 68 04 08 5A 1E A0 16 88 7A 70 F8
 40 C8 2B 01 0B 62 02 1A 2A 93 E2 45 BE 8D 95 94
 15 C3 1F 5B 55 B7 46 7E A5 65 1E 8B AD 21 62 ED
 95 65 13 08 CA FC DB 20 8F C9 88 7E 6E DB 6E A9
 C7 A0 D7 14 7C 0D 00 24 BB E9 93 CD D7 22 BA 1E
 39 13 64 2A 33 29 4B 12 02 0B 9E 77 2E 76 B2 2F
 B0 08 EB 50 C1 15 2E 8F C9 24 AA EA 29 EC 30 F3
 66 C3 50 B5 A1 28 9E C5 41 B2 A8 20 60 FA 44 FB
 39 61 A9 51 A5 9E 52 C8 73 6D 92 F3 84 34 B1 7B
 46 FF BE 68 B4 91 0C D8 90 B4 A7 25 74 13 61 59
 D2 8D A7 37 4A AF 34 F7 1C 92 C2 B5 F9 A3 97 4F
 07 A3 1E 3F F0 11 CC 39 62 08 30 0D E7 84 DE 9E
 32 84 BE D2 82 D0 D1 86 38 E9 CC F7 9E A4 0B 31
 3E D6 58 E5 41 B1 36 7B 07 6A 0E 50 0F 16 CC 56
 D3 0A AC 58 6A 1B AD 87 84 23 38 B0 9E E1 20 D6
 85 DA E3 D2 ED 07 C8 12 66 45 E3 FC 9D 5C 1C 2E
 4F F1 36 32 07 5E 2D EE DC C0 D8 CE AE 39 1F 59
 F2 CD 8C B2 AF D4 B9 8C 9B E8 E2 05 12 E8 A8 CE
 3E 1D 09 E1 F1 24 1A C7 38 C3 3D 36 DB FF 56 53
 10 AA AC 59 17 E5 BA AE A0 D8 3E 3C 2E 6A 18 AF
 22 E2 80 B5 AF 52 1D C8 CF 4A 1D B5 8D 3D 62 70
 73 5E 9E 66 30 F9 AC 19 E4 94 4E 49 76 DE 70 D0
 21 97 26 72 AF C9 8A B8 D2 F3 A4 32 B9 B0 61 F1
 FA ED 39 BD 3E F4 C0 3A 14 D2 B2 97 E6 52 18 91
 6D 9C 3C FF 37 24 D5 77 85 59 1D 1B B9 A5 FF BD
 F2 56 24 0A 70 0B 94 4F D0 17 65 C6 68 91 53 1E
 4F 10 26 BD 24 30 9B 24 3E CD F3 50 8D 23 75 A8
 9E 25 7E 4E B8 B5 4F 1B B8 5C 72 80 40 55 05 41
 14 14 15 99 5F 0A FC AE CB F4 68 28 58 34 7D EA
 E9 EC 3E F3 2F 7D D9 5D 0F BB A1 CE 8D 84 59 E9
 D9 19 CF 03 C8 62 E6 4D 3A 1D 2B 3A 6D 65 37 AE
 DD 9C 7F A8 B8 99 16 03 7C 8F 94 B1 4E 1C 8D 32
 37 B9 B9 02 BF 0E C2 5B 54 89 F4 C8 1A 60 EC 85
 57 10 0A DF 55 05 08 CD E7 35 62 45 95 0A B2 29
 21 7D 58 48 3C 73 91 5F 59 80 FB CC 40 ED AB 17
 EA 5F 2E 30 78 71 9B 29 72 65 03 68 30 A3 26 FD
 AC 6A 75 95 9D 72 F8 54 83 EF 2A C1 64 50 68 08
 73 6F 17 AC C8 71 59 90 C4 1A C0 D1 C7 BC 6A 0B
 24 01 DC D9 5D CC 41 F5 D3 51 BF 0D DF 9E 32 F5
 95 F2 97 5D 2B 9B 4C 7D BE 41 53 F0 D9 C1 93 77
 8D 7B 18 0E 25 42 70 B6 19 5F E4 97 20 63 41 9C
 8E 4F 59 53 B8 38 21 28 C6 7B AA CE BD 56 5C 56
 FA D0 AB 1A DC 37 83 2B B3 47 12 93 B9 01 39 CF
 5C F1 DB 31 BA C5 D3 4B 16 02 A1 E4 5B 02 B0 20
 F9 57 91 F3 DE E4 ED 8E 05 3C 83 42 1D 8C 48 27
 FA 8B CE BA 23 8F 94 99 E9 95 26 C1 64 91 E4 3D
 FB 77 7B B7 F2 BF 0D 2F 1D 22 B2 0A 20 CC 6A A9
 76 A1 FB CB 49 3B 24 23 DC 0C 3D 87 21 CE D1 27
 8E 37 08 BF 96 3C CC 8E C2 2E DA 53 DF 7A 6A 70
 AA B0 25 B7 83 79 65 53 8D 2E 62 3A A2 56 6D 1E
 EF 8A 78 B6 D5 DB 61 18 49 19 50 63 A4 76 66 25
 B4 3E F8 8A FF 82 F7 2D 24 E8 8A D7 E3 5A 46 9D
 D9 71 89 C1 20 5D 69 6B 34 FD 10 34 29 F4 57 C7
 88 03 CA A6 B5 BC BC EF 2C 56 DA CD 72 58 59 80
 48 05 C9 11 4F 3C D0 1F 2B 41 19 D5 CE 95 1F BE
 E4 E7 62 B1 D8 10 9C 44 85 04 40 23 28 6C 19 D3
 A7 37 1C FE EE E3 A5 98 B2 97 A3 56 DA FD 32 34
 D3 B1 F8 F6 47 66 4E F3 18 77 30 AE 49 39 E8 07
 1B E1 39 59 2B DD E3 CE 23 06 12 DB F5 07 5C 3F
 C7 CA AC E7 ED 8D B5 BC BE F9 4A F8 FA 54 31 E5
 2C 73 7C 86 27 B7 50 E1 9D 10 E7 BE B7 45 54 40
 F5 52 45 49 C5 E0 8E 62 72 EF 81 B9 3C EC A3 81
 B9 D3 2C 46 65 26 ED 38 E1 C5 C2 51 14 D0 39 F9
 2B 75 BB 59 E2 B6 06 02 6B 41 63 29 12 3A 9C 24
 DC 24 29 1C 2E 47 F3 A4 A7 4A 75 CF 6B 33 02 FA
 87 DC 42 69 E3 43 0E DD BF 23 4D 24 11 13 3F B7
 48 C2 3A 3B 39 DA 12 9F 1E EE CE 1F 51 BE 3F F5
 24 4B 9B 57 27 B4 4E D5 4F 0B B4 18 D4 7A 1B 8A
 4A 98 1D 84 73 69 1A 86 E0 2C B5 33 26 DE 22 51
 89 41 62 71 E7 8C 3C E5 F6 AA 85 2C 50 7D 2A 0B
 CE BC 09 4B C7 63 E8 50 CB 4C 8F 93 D1 A6 D8 15
 92 65 02 AF 1E 74 E2 93 17 A8 8D 1F A4 B5 CF D8
 70 AA 37 77 B9 31 DE B4 B4 50 83 03 CC 9B E3 F3
 9A 06 E3 EE 20 70 4E C5 6E AD FD D2 02 6E 96 CA
 9D 1D 3E E4 0F 97 8F AD 1A F4 8C 8F DD E7 A8 1D
 5F 86 95 74 5A 2F 30 9B AC 71 B2 2B 82 F1 AB 57
 76 FB E5 A1 F2 79 D2 0A 3C B3 C9 AB 1B D2 C8 F3
 AB 7D 68 54 3D E0 3B 98 FB 0D D7 40 9F 8D DA F4
 83 04 9E DC A2 7C 73 F2 A6 4B 0A A9 6D 7D 0B 5E
 C7 F6 4C 4D 29 5B BE 04 D0 AF 0F 5E E5 B4 FB FB
 17 D8 49 4E 00 98 B6 9F 6B 06 70 8B 87 B8 F2 A2
 86 7E 0D FF F7 27 A6 E4 66 CD 17 B8 2A C9 7F 22
 2E 07 5F DD 03 C6 69 E8 AD 23 01 E8 D8 03 7D 0E
 1A 90 87 B1 73 AF 45 87 D4 14 BC 4F 9B FC 73 83
 41 46 77 6F 66 E9 5E 8A 8F 3E 88 30 44 2E E8 65
 BA 60 B0 3F 5D 7F 95 77 60 7F D9 2F DC B6 3F BC
 80 9D 59 E5 E0 87 B1 A5 FF 5C 72 3E 40 0B 32 84
 BB 11 86 17 4B 4D D7 79 A9 A0 62 A1 56 3D 83 E4
 16 B3 97 BE 19 63 55 13 8D 97 56 21 0F CE 2A D6
 5E 82 35 C6 0B 22 34 EE 74 D1 11 85 D3 7F 32 2D
 03 32 BA B6 44 E1 8E B6 41 13 40 FE 7B 13 D3 2E
 3F F0 8E 2C D6 69 8F 60 67 CC 9B 0E 6B 38 11 0A
 16 E9 4E 99 47 AD 20 4E 32 FE 12 EF F4 17 E7 F6
 34 57 A4 7B 19 23 88 9D CF 98 E2 A5 EA DC 82 40
 54 7E 5D 51 CF FA D8 3C B1 6F 06 22 15 0C 51 66
 6E 10 11 7D 8C 59 F5 5E BB 04 13 18 F2 A4 85 F2
 58 50 C8 59 3E 6E 03 F5 26 BA 0A 03 DA A2 8E 29
 94 76 1F 51 02 23 FE 1D 7C B3 72 33 CF BF 08 5E
 E1 E9 8C 60 02 DE 74 F2 8A 7D 3E 96 72 EE 75 D9
 2C A0 19 29 32 A5 38 39 A8 34 D3 64 0C D6 40 D8
 61 C3 16 4F AC 5E 17 1A 4B 7F 1D 99 5D F0 2B 15
 92 6E 52 95 8E 54 72 CB EE 54 83 30 79 E1 BC 4B
 4B 0C 05 04 FE E8 25 2F D7 64 44 72 23 4F 39 88
 9F 19 1D 59 28 AB C4 38 9A A4 12 E0 51 EA 17 14
 29 FE 2A 91 B4 7E 7C 6E 49 67 43 8D 11 3A 5C 33
 18 FF D8 CF C7 48 A8 5B 85 DA 79 BE A2 5C 09 A3
 21 71 82 77 5D 18 0F 0D A3 80 F7 62 BE 1B A0 70
 26 65 D1 CB 5A 97 AB 0B BE 2D F0 73 FC FA 46 17
 B8 8E 25 45 F6 4E E6 BE 18 0C CC AD 70 08 D9 82
 4A 72 BB 32 82 3C 2B D9 73 74 4C 02 85 4D 67 B7
 97 C2 0A DB AE B0 1C A0 03 FD D9 90 F4 40 FA BD
 24 7B 12 BC A7 50 4F A6 5D FC D1 36 B1 4F 3B D4
 70 10 77 95 D2 A2 6A 78 99 92 99 DD 8C 2B AB C6
 21 1F 2D 84 20 0A BC 7B 10 76 7C 1E 11 46 76 F5
 7D 9F C5 2A 99 30 8E E2 CE E0 E7 F4 82 3A 26 09
 8D 6C D1 48 B7 70 A4 D0 10 B7 F8 0E 2D 77 EE 4C
 1B 0E FE AD E3 1A B6 8A EE 63 3C BB 24 8C 18 47
 6F A8 DE F2 7B B9 B0 8E 0B 84 1A 22 99 04 A6 38
 4A EC 96 D1 6F 6C 3C 74 F2 E3 12 4F 4E 58 EF BC
 22 91 C0 A2 0E 87 9A F5 FF D5 D8 D2 75 6F DE 0B
 5B 8D C2 98 79 6A 49 14 86 13 C2 A6 67 58 CF 5D
 B9 45 A0 11 F0 13 7F BA 03 7A 1E 45 46 0B 8C 92
 7B 21 E2 50 C5 A1 DA 4A EB E8 DA 97 65 A0 25 6E
 64 E6 F4 54 7B A7 FD BE D9 54 D5 12 B0 86 B2 61
 66 DD E1 8E CF DA 9D 89 08 74 31 DC 7F A0 8C B1
 89 8F E1 51 6F DA 15 70 49 7A DB EE 9B 62 59 13
 21 47 A6 08 86 A0 48 93 46 6B 78 71 C1 99 25 B8
 98 38 52 99 C6 FD 9A 1E F5 BD E8 FD A4 BA 8C 87
 C2 22 4E 26 50 2E 1A 3D 02 67 C7 BC E6 EA D8 16
 80 64 17 76 6A 31 80 19 A6 2B BB 68 4F DB 12 0A
 3A E0 B8 3D C5 D0 26 EA 91 62 D2 F0 37 D4 FF 15
 35 D5 7E 77 68 52 E4 97 7F 71 9C A8 10 49 03 0A
 AF 76 AD E0 17 F9 1B E2 72 A1 0E 1C 32 62 3E 27
 36 DE 93 87 9B 29 E4 91 38 9C 0F 73 AE 34 0D 46
 97 D2 68 B4 6E 2D 06 BF 4E 98 4F 0F 70 E0 AA E6
 CC 82 BF C3 E6 11 91 3D B2 3B AE BE 56 43 84 3D
 F8 C2 76 17 41 48 55 89 D9 95 F6 95 AC B2 7D F1
 86 9B 16 36 C8 62 7B 90 F7 CD 84 0B C7 3C AA EC
 36 5B A8 2A 70 63 C4 95 2A CB 3C C9 A3 49 56 1D
 B2 4E 8D 50 79 F1 E9 27 DA 78 CA 76 E8 DD 13 1A
 A5 97 B9 5B C1 2E EC 2F F2 3F 97 DD 13 6D 89 15
 D1 05 82 D7 45 AE 5D CE 12 71 86 42 7F 5E A0 61
 09 FA 54 03 96 80 42 59 84 B5 03 19 5F 76 82 9D
 27 34 DE 99 A7 DC 66 54 E3 93 97 11 96 FA 1C BD
 85 A5 5B F7 6E D5 37 61 B9 FF 92 CC 62 E4 89 AD
 96 78 DD 5E B5 67 FC 06 27 48 52 7A 5F 8D 25 49
 9E 57 B4 F5 53 45 F6 C9 E4 77 60 53 0B C7 3D 22
 31 09 6E 5B 1B 8E B8 B3 7F 89 ED 6F 62 03 8F F0
 1E 95 0D C3 2A 47 46 B5 6B FE FB 8D 83 B1 D9 52
 EC 98 4F 9C 34 A7 B9 82 50 89 CA 48 45 F6 BE AE
 C4 36 C8 10 0D 14 06 02 F5 2F CF 39 5A 4C 4A 4D
 E7 52 FA 75 59 86 8E 37 3E D3 7B 24 40 81 DB 8F
 2F 00 2F 52 21 FC 4E 16 28 0D BE C5 69 6A 25 C4
 7A 83 25 B8 E6 D5 19 06 57 5B D9 18 57 21 7F 27
 0F 91 04 23 E5 18 D2 5A B3 72 0F E4 16 96 74 A8
 39 D7 E8 32 89 B6 96 EF 2E 54 49 45 5F BC C8 E7
 7D 70 40 6D E6 21 B2 9F FD 59 42 CD 7B E6 B6 81
 4A 53 C1 20 82 F9 A7 89 1B 07 1D DD 8B 41 A2 0E
 70 D1 8C F6 CE 46 7F 35 1B FC 25 00 A2 A1 E6 AB
 0A 59 4D C6 40 52 9A 30 3A 3C 36 10 32 1B 68 D7
 16 E5 12 1F 4F B8 78 57 8F 64 9A DE 30 64 43 93
 20 1B DB 31 03 97 76 36 82 78 B6 D2 94 25 B4 50
 9D 25 9F AF AE 63 90 ED 76 1A C6 C3 74 F9 1C FD
 6B 01 3F 9F F4 9B A8 D9 0F 8D 45 F3 32 C7 EA 13
 52 36 B1 18 03 EA D1 0D 97 9F 8B 2B CA 53 9F A7
 25 FF 3B DB 11 E3 AC D7 B0 89 E4 0F 57 20 D2 EA
 25 5B 3C EA 31 7B 65 88 81 A6 13 83 79 09 EE 74
 A9 86 72 96 69 C2 C8 F0 41 FC 3D 0E 87 F9 C7 4A
 E1 15 32 51 1C 3D 87 79 BC DA 96 B1 10 3F E1 FD
 49 C8 31 B6 27 85 27 89 7B 46 02 A3 78 49 BC 74
 4B 63 B7 D2 3E E2 73 2F 83 A0 18 09 63 A7 8E 50
 E5 00 B0 11 04 81 9E 12 2B A6 DD 61 5E F8 D4 09
 82 E6 D8 6A 82 16 49 0A E9 EA 94 5A 5C CF 00 03
 F2 A8 75 E6 55 83 97 44 0B 34 A1 9B 5E 90 1A 1C
 C1 8E B5 E1 A0 1A 0A B8 56 81 BF A2 1D 20 59 31
 37 96 34 14 1F E6 42 10 12 B8 88 59 4C AF 61 D3
 CA 36 BB 9B B2 11 D5 C4 50 BD 83 4A 79 6A 00 52
 14 51 04 26 64 2E A6 F1 77 15 A3 36 0F D4 48 EE
 1E 99 7F A1 4F 90 66 E8 BD 3D FC 53 6D 8F 15 59
 4C B5 B1 3C C9 6E EB 01 DD 90 15 E0 77 CD 20 D9
 5F 55 1F 0D 7B C1 C7 F1 29 D9 6E EA A8 CF 6B 46
 AD BF B5 30 DC 26 29 94 BE A1 BD CF 30 A7 2E 29
 D9 0F F7 58 D1 39 BC FA 25 A6 B0 26 38 E9 6B C6
 78 C9 C7 8A 3A 93 74 93 35 95 48 B8 68 5F 46 66
 A7 9E 5A A3 DE 13 80 2B 4C 03 4F 80 67 6A 76 3B
 A0 0F 98 11 80 48 46 2A 51 87 4E 71 B0 17 55 AB
 10 F8 41 E9 38 B2 78 EF 77 F4 27 AD 91 20 54 1C
 82 BB 3F 52 2E 68 EF E2 E5 32 44 6A 8E B3 35 1F
 33 30 A6 E4 C9 48 91 A0 99 7B CC 0F 6D 5C 33 15
 AE 28 A8 C1 96 B5 E2 6D 46 36 8A A2 8C F5 4E 57
 B4 F3 22 6C FF 9D 42 03 3E 06 E5 DC 16 F6 D2 1D
 FD FD 94 31 E7 AB 45 DA CD E8 C2 A7 47 7B AD D1
 21 9D A4 5F E3 76 A0 85 E4 0A 4C EF 2E E8 CC EC
 AF AB F4 6D 5F 99 FE 0D A8 2C 70 A2 D0 EE 88 42
 80 53 F0 B5 E0 BC E1 E1 A9 37 30 72 F7 E0 0F 86
 AB 4F 62 FB 0A 3B 6B 5C 6E 0A 0A 02 C3 E3 69 9C
 C4 05 74 5C 4D C0 0D 94 E9 45 3D 02 D4 37 AF D4
 C7 03 F1 58 BC E6 65 71 A3 20 76 42 5E E5 9B D7
 7F A2 96 D4 19 73 19 C4 C0 B9 FA 2F A9 DC 83 01
 BF CC 37 2F CA 20 57 5D D1 D1 BC FA 98 59 3B 01
 75 24 D5 43 83 B6 5C 33 CE 7B 56 39 E1 21 F5 CD
 79 4D A5 DE 7B DA 28 68 33 CC 67 2A A6 CB 6B 9F
 30 52 2E 75 41 40 A6 E6 E5 56 88 2F 64 23 6F 46
 0F D9 CE 25 FB 97 8C 1B 13 88 B9 4C 2B 71 44 DF
 C3 06 EB C8 91 CF 72 32 55 15 F5 66 DD D8 28 B4
 EF 6F BC 99 87 E3 F4 AB FE 49 9A D2 59 97 5F 62
 75 0C E6 D4 E0 DE DF 9E BB 56 61 1C AD 9B 59 95
 C8 C2 34 A0 01 87 9D 60 99 FF CD FC 79 4B 46 9E
 0B 40 10 20 4A 14 98 91 AE 15 2F 82 BE C4 F7 CD
 3E 84 AA 79 96 0A E3 23 3D AC F6 D5 96 81 91 54
 94 B1 EA A2 8D 83 85 CF 58 5E F5 5E 12 F9 49 C3
 0E 3B 8F 0C 06 5D 2D 31 CD B7 8B 00 06 29 24 23
 1E 20 C0 F3 61 D4 61 91 80 91 30 2D D1 8B 01 49
 E1 A4 C8 99 FD 36 3C 38 DE 56 36 3C AD CF 73 84
 A5 BF A8 D7 16 29 B7 6F 5A 62 6B 71 03 2D 94 2E
 43 6B 01 40 12 90 77 1A 5F BD 1C DC 59 5D 05 BE
 A6 12 94 C9 13 79 17 EB C4 8B 9E A5 33 87 FC 9D
 DC B1 21 A6 4F 4C CE 87 80 B5 FF 03 3E E0 23 7D
 1F 23 F6 A6 AE 36 A7 68 20 CA 39 0E 1E 77 47 BF
 2A 95 DE FF 05 E5 00 A3 A9 9B 68 1B E2 6F A3 56
 BA BF 97 06 ED 63 83 E3 D9 FB B2 2A 2D A4 09 E7
 51 51 D0 CB B9 E0 09 CC 0B 69 D3 9B B1 C9 F0 91
 8E 37 77 CB 61 FF FB 5F 35 C7 B4 5C EA 20 91 CB
 1F 79 B3 CC 40 0A 7C 02 7A 2E D4 50 6D C0 BD 4C
 B3 36 7E C1 ED CB 7C DE C0 E6 E0 16 B0 B7 A1 ED
 B3 9A 79 4A F0 BA 9B AA 46 5F 11 AD CB EF 61 36
 C9 7E FD C1 EA F1 A8 EF F4 6B F4 92 61 6D F6 AA
 BB 9C 26 49 21 8B DC 7B 4F 5C 09 C9 5D 5C 1C 4F
 12 3D 12 CF E3 D4 A5 49 22 64 99 68 8D C6 F8 E2
 8A 95 79 0C 9F 24 45 86 FB 83 3E 74 45 D7 A5 09
 50 FA EB E0 7F 21 43 8F 40 56 57 47 34 96 5B AB
 EE 4C D8 52 3E E4 7D 58 91 60 AB 2E 2F 23 1D 8F
 BD AC 67 53 B4 4F 3F 76 39 D9 A2 86 A4 15 B4 4F
 C7 3F DA 1E B5 06 4B 51 D5 59 C7 C6 1E 96 A3 59
 28 AD 99 07 96 41 5C 15 83 93 8C DF 28 DB 7A C6
 5D 6A 4D C9 B4 D7 62 0D E9 EC 34 CB B9 09 B3 27
 6C 2B 5E 15 9D 27 A4 2B 1D 23 EA 5E 39 02 D7 45
 DD 35 CE 17 A9 7C 27 2D ED AD B3 8D 8C 4C A8 83
 86 2A 65 54 B0 54 29 7E 8A F6 F0 F1 F0 85 F5 B4
 F0 ED 82 25 5E 25 59 32 2A AE 35 3E D3 DD D2 B8
 B3 13 64 A6 83 30 36 F0 48 97 81 A3 2F 42 94 DE
 91 C9 6E 4F E3 9C 38 33 AC CA 58 37 04 58 A3 4D
 B5 EF 0F 75 43 EF 23 47 15 C4 D7 E8 33 CB B5 59
 7E 05 BF 37 69 18 9A 33 3D 42 49 1C 3B B0 6D A5
 8C 16 B0 BE AC 89 1B 79 43 F5 A8 87 C4 86 4D 88
 0D 93 87 B9 4F F1 70 1C B9 7E 0D 08 52 5E CA C8
 94 2A A5 07 B5 4C C9 5D 04 BA 10 BE FF 6F C9 92
 25 38 80 4E 9C 03 6E 22 32 98 EE F1 13 14 D1 C6
 29 57 88 D6 A3 4C A5 BD 5F 22 E0 FF 46 8E E0 81
 C9 D3 D5 E4 B6 CB 27 4C 83 1B 0A B8 C7 23 C6 3A
 A1 22 95 77 05 B0 93 9F 6E 9E 1F 36 98 87 BC 0A
 88 96 41 A7 BE 52 4E D4 AF 56 AB D1 D2 E1 F3 E7
 2B EC E5 E8 0F C3 E3 04 12 C1 AF A5 A0 06 EE 6A
 A6 12 4A D5 C6 58 47 07 2F 08 76 6F C5 3D 69 35
 1B B1 5C A7 EC C0 9F F3 C6 38 0A E0 FD AD D5 2A
 7E EE 3D 19 79 89 0C 4E 26 AF F9 B3 49 4F 77 1D
 CA DC B1 71 1B 30 1A 97 A3 89 D6 6C A7 65 4B D7
 EC 05 E9 19 FF 72 BD 83 91 CD 05 DD 19 8E 23 37
 32 1A EE 37 C5 E0 8E 4B 07 98 2C 79 A6 59 AC B2
 63 7B 96 74 21 DA 4F C2 F8 EA 8E 39 52 3A 3A F8
 BF A0 91 58 97 63 20 71 80 9A B1 4F B9 AE 27 3F
 1F FB 38 6D E5 0A E6 2A 27 F3 F0 78 EA 3A 11 11
 33 F0 F7 84 EB A0 80 76 5C A4 66 1F 2C B0 B7 59
 8B 96 26 5C 48 51 13 3F 6E 73 69 5A 48 D6 81 C2
 A7 32 88 88 2C 8F BF 9C 3F 55 F8 DD 51 BB 28 90
 E2 D4 28 43 7A EF 4D 95 6A 3B 93 E4 96 78 83 D1
 52 64 22 17 F3 27 F0 E6 43 FC 0C A5 01 1F E9 CF
 C7 21 91 4A 00 0C 05 20 A8 82 85 8D 91 B9 DD F2
 6C AB 21 C5 E8 21 FF B5 07 02 A6 E0 7E 91 CB BF
 79 0D 64 42 1C 77 FF 37 D0 6A 15 B0 CC DE 95 DF
 0D FE 5A C8 D9 45 8D D4 09 AD 08 7D 0D 68 6F F2
 9F 98 89 43 61 EF 43 98 77 05 C0 33 13 30 25 22
 04 90 A8 50 A2 6E 88 D6 A1 FD F8 DD EA 19 C8 C3
 29 87 C6 04 E3 A3 39 84 30 40 E2 6B D1 78 DD 02
 54 29 37 C2 7C 76 AA 58 25 A5 00 5D B8 21 57 55
 0F 63 5E D1 8C 23 F0 A3 CF 05 62 A1 22 8F 95 96
 B5 22 A8 CB D3 BD 3A BC 8F FA D9 B9 D0 6E 13 01
 04 91 11 E9 A7 9B ED 09 A2 8C 49 EB B4 BF 5F 58
 D2 F3 80 D7 98 5A A6 DA 23 B9 79 41 F8 D6 40 A0
 A3 26 EF 65 DA 1D A0 38 27 4C FF 3C 27 F4 A6 88
 BB 02 23 12 B0 9E 50 5C 4D 9C EB E6 A4 1D E0 A0
 81 F1 B3 35 B5 EC FB 71 35 B3 68 05 E0 B2 3C B1
 D3 B8 96 E5 24 33 D2 45 2B A9 E1 9E A6 56 6F DA
 F7 0D 0A 3C EC AE 4A B2 F5 BA 29 65 CD 84 F8 0A
 D6 F9 B4 86 AA DC 05 F7 B4 48 1F 02 AA 70 3A 6E
 B5 59 C3 45 61 D1 44 BC 18 9F EE 97 E1 3F 79 E5
 8F CE BE B8 6B 03 CB C5 CD 3E 98 D0 86 00 AE EB
 E1 01 25 31 E1 D6 FE C6 0D 70 BB 90 C7 A6 C9 0A
 1E 7F FC B3 7A D7 4A 73 8D 1E CC 33 2B 13 D9 E7
 1C 6A DA 3B 99 B2 AB 9B D8 9F DE EE 6C 90 77 26
 70 8D 67 1E 3D 3B 92 59 D6 78 F4 F6 BE B3 8F AB
 79 91 CD 83 8B BE 49 68 E0 40 91 A6 B0 0F F1 39
 33 01 8F E9 15 09 A4 6F AA 34 0E A8 70 19 40 4E
 A9 CB FB 2B A6 AB 07 C3 84 F9 87 36 92 C9 C6 97
 86 8D 4B 73 D4 FB CA 78 FA 7B DD 36 C2 20 7A 2C
 64 5C FC 90 3A 40 0C 4A E5 11 AD 87 64 D1 53 60
 EA 28 56 44 4F B3 F3 16 25 46 7C DE 99 FC B2 CB
 53 D3 CF AE 9D B6 8C 40 EC AD 1B 06 EF E7 7E B1
 28 D2 69 5E 32 44 81 85 BF 7B 44 69 52 10 2F 0A
 E2 4B FB 6E 4D E7 06 1D B9 6C 17 81 A3 7D 1B AB
 45 3F C0 BA 65 A5 D7 91 68 8A 5F 4E AA D5 89 BB
 08 BA C7 1A D7 19 31 AC 25 EB 27 ED 59 F7 92 77
 19 55 34 4D 41 C4 A8 B5 3A F0 0A 9E A5 5D B9 39
 9C B2 56 A1 7B 24 8D 19 0B C1 EA 96 D1 35 BB 55
 47 F5 1A 64 CE 52 CE EB 67 A0 9E 27 DF 47 F1 A9
 51 E7 78 0B 2A E5 3E E9 BF 5F CB 00 5F 88 A5 94
 CF 94 4F A8 48 F2 E0 8B 0A 3E 9A 4F FC DB F2 6B
 E1 5F C6 FC 82 DC 3D 0C 66 31 D9 FF C1 65 C6 31
 5A 28 5C 70 1F 99 98 9B E4 1C DA 1F 9D CE 88 0C
 D0 06 A5 57 A8 28 DB D4 C5 ED 5F C7 17 65 43 6E
 1F 32 17 2C 05 36 81 47 26 5A 22 02 6D A8 07 43
 A8 63 CD 12 EB 4D 50 E8 D0 74 B3 EE 02 C9 BF 81
 11 98 D9 D5 CC 23 0E 01 A3 FE D7 55 93 48 5F 6E
 69 76 26 A0 CB C6 6F 12 F9 2C 37 07 D5 89 E9 E2
 76 79 AB 04 29 01 1A 1C E0 40 3F 02 A7 4C 58 2D
 B5 EB 0E 8F 83 C9 88 F3 EC 28 39 4F 63 5E A7 4D
 CA 0E 1C 8B ED C0 11 37 B0 32 5F CD B1 66 01 08
 42 85 B9 A9 CC 8C FC 8D 2C 24 86 76 F1 D5 D6 3C
 5B 19 B6 79 3B 1B 9B 11 EB F2 E8 55 64 3E 5E EB
 E3 CE DC A5 C6 19 7C 78 8F C1 99 D8 8B 9D 26 AB
 9F AF 5C 9D 3C 8D FB 16 D6 ED CC 31 54 5C E3 AE
 2C 35 97 CB C3 5B F5 6F AA 75 B8 95 11 7F 6E D8
 52 2A C5 33 97 23 EF F5 DF 5E AA 84 1D D5 21 1F
 C0 90 F1 53 76 CE 8D F5 EB 07 C1 3C B6 C4 48 9B
 5F 8C 93 BD 12 D4 B4 44 2A 0E B4 6E 20 2D A0 7A
 C9 C9 A8 25 31 6F A0 8F 06 6C B8 88 4F D0 F0 6F
 8B 45 F8 5B D3 DC 29 6E C1 47 73 B5 CE 8D 31 51
 2B 39 03 41 BD FD 37 8C 78 27 20 EE 2C BE 39 3E
 B9 7E 94 84 84 52 CB 6C 24 90 A1 79 02 FA 31 85
 19 32 0F A0 19 A1 B5 54 0E A0 B9 73 9C 42 70 3C
 38 E2 63 17 F2 DE 11 B8 15 68 A5 4E 66 A5 38 BC
 65 0A D7 7C 1D CF AD 4E 24 57 91 6C 02 A5 90 DA
 19 5C E6 14 05 ED D3 9B 90 8C 58 6B 74 C9 09 F1
 33 DD F5 C9 CB FD 19 77 E0 8D 99 2B B5 9E C8 2E
 DE D2 47 E4 BE AB 66 9F D5 27 5D 55 31 15 27 B4
 C7 35 0C 69 56 22 15 28 8A 2D 59 5A B2 58 6B 9D
 4F 4C 73 03 FB 6F 41 45 08 18 95 B3 7D 9E 6D 74
 AE 0E 27 A4 A8 6D 96 95 7C 6E 4E C4 3F E9 58 DB
 A9 31 05 37 29 43 5E 10 22 9E D9 7F E7 58 80 0F
 79 77 8F C9 2A 8B EF CC 94 76 92 8A AA 2F DD EE
 86 D1 6E AF 76 EC 62 43 CB 7B 77 14 AF 8E 7E 6A
 C9 55 7F 19 B1 FB 9A E9 E7 2E 05 58 1B 49 B1 6F
 CC F2 EE 37 0C 97 D3 15 CE 15 1A 67 9C 73 B2 6D
 B5 D3 D3 7F 21 D1 6B 12 10 2F 3C 8C A6 DC 9C 28
 A0 09 B6 83 7A D3 77 32 FB 60 FA FB 93 E6 E8 DD
 CC 27 E6 37 3B 63 ED 98 21 FA B0 9F E4 23 C2 B2
 15 A8 07 D8 86 D8 BC 7B 01 90 01 C7 2F 3B BF 3B
 28 9B D3 59 13 B2 B8 9D 99 27 D2 20 24 31 F7 12
 D1 6F 91 02 4D 8E ED E1 CF 4B 38 C6 AF A4 0A 7B
 96 CE B8 96 E5 53 F4 59 6A 9F 0F 76 33 89 6D E0
 C9 66 60 79 E1 F1 F3 DC 41 D5 14 83 6E 80 97 60
 64 8B C4 FF 3D E3 75 A2 29 6D 4F B6 7A A1 58 1F
 3E 5D 07 9F 37 A0 4D 30 CF 62 92 62 86 CC D6 8D
 2D 18 24 BF 4D C5 E7 64 08 5F ED 5D 3E E3 1E 9A
 07 E7 75 E6 2A A3 4C 92 9E 6E 0B 07 E6 72 EC B4
 AB 16 0E 58 30 F1 C9 DF DA 36 13 4A 4F BC A6 7B
 F1 96 84 D3 66 36 81 F7 85 A4 38 EE EB D4 A4 81
 CA CF B1 B1 C1 32 AD 2A C9 FE CE A1 D5 7D 55 EE
 4C 7C A1 8F FF 3C D3 BF 66 D5 A4 5A 2D 61 2C D9
 48 78 F9 BA E7 17 5C 75 70 E2 C8 96 27 75 66 D9
 C7 EC 4A 4C CC D7 A2 AB B2 C2 9D C0 FE 44 A6 B1
 94 96 DC 55 56 7E DB FD 40 89 1C 4A D4 FA D6 53
 AD B0 D0 C9 62 6E FE DD C5 A4 5E 6F DB 86 99 39
 4B B5 67 E1 8A 2C 93 3E 43 5D 7C 13 4B 9F E7 D8
 7C C5 8A E2 2F 25 CC 1C 6E 68 54 07 5D 84 03 A8
 01 A0 16 D1 B2 12 9D 3B 4C 9E B0 97 24 62 9D D0
 DF F3 45 CB 44 7B 59 AF DF 87 AA 6D 5E E6 15 30
 6B 11 0F 33 75 E5 94 B4 79 3A C2 35 11 44 46 38
 CF 05 DB 7F 7D A7 F8 55 00 F6 8D 76 97 4C A3 49
 99 1D 34 E7 93 10 85 82 4D 57 17 86 83 4E F1 2E
 8B 8D CD BE C1 1A 2D 1A B6 35 69 F2 39 D6 74 6B
 F5 1E B4 B4 9F D9 6A 7E CF B3 48 D7 D2 E7 F7 B2
 BC FD 1B 1B 97 6C 74 63 82 2F 3A BC DC 21 A5 0D
 2E 07 5B 13 D3 84 C3 27 56 43 74 BF CD C9 89 B3
 1B 05 6E 11 6D 63 EF A8 0E 02 C5 16 71 60 DB F3
 52 A1 07 80 46 81 AD E3 74 96 F0 72 B9 57 57 F9
 78 42 F1 59 0E 1F 78 67 11 2E 6C DD FE 0F C5 D2
 AA 64 4C 93 A3 D8 C4 9D 7B 92 CC 3F 27 48 85 74
 49 95 06 B4 BA 73 BE CB A2 F6 43 51 BB 18 EF EE
 A9 6D 5B A8 84 9F AA F4 C5 F5 84 B1 E9 85 BB 4F
 0E 40 58 EC 00 2B 3A FF 7E 78 AD 2F EF EB 35 0E
 7D D7 E5 47 BE 46 59 88 26 37 3A CC D7 95 8A 0C
 41 96 3D 99 FE C4 EF DD D9 6B DB 06 AB AE 5F 3C
 31 E0 80 D2 6B 8D D2 9A 37 89 13 2F 5A 06 F2 08
 2C 59 70 12 19 1A A9 05 EA 2E 90 52 2E 63 7E F5
 98 EE 7C 2F 78 03 F8 23 94 A1 76 45 8B C3 4F 2C
 5A 9C 37 CA 20 B8 18 B5 D8 FF 6D E4 3A 9E F7 65
 66 E0 AB 9C 37 E0 80 BD 31 2B 37 9B E1 7C 56 4E
 BB BE 36 FB 3C 56 69 04 66 F3 7A 0D 65 4B 21 7F
 3D 71 55 B9 70 54 EF 6C 55 D3 EF 5A 72 2F 72 BA
 81 ED 7D 72 F3 7A 64 CF E6 38 BE 88 6E F6 B8 16
 42 51 7C B6 A7 7E 41 43 C1 25 16 50 E0 62 8D 27
 3A 95 52 E5 EB 7A 0C 9F C9 BC 6B 3D 23 FD CD CE
 D4 6A E1 96 67 8F 6B F4 4F DE 3B 05 EE F3 DB 47
 E2 B2 F6 1A 8B 37 81 B7 23 5E 89 4E 3C 87 60 FD
 13 01 B3 42 47 FE 9E BF BF 21 FE 65 29 4B D2 FF
 EB 90 EE 44 CA 70 0E D9 EE 66 68 6E D3 14 CB 66
 C8 83 EF A7 A8 CB DC 77 D7 93 09 D0 A8 DB DD CA
 A8 75 97 1E 79 21 98 4D 2E 8E 86 79 6E CB 9E 7B
 B0 3E 97 38 F9 D2 BD CD 4B D2 7F DB E5 E3 CC 9B
 30 4D 5A 56 8C 60 4D 81 23 24 07 E2 3E EC 1E BA
 11 80 0B CF EC EE 5B 42 C4 C6 BD 59 08 6B D0 E7
 4C 69 E1 F2 05 1D 4B D8 68 AB 8E B7 2D E3 67 F9
 B2 35 59 9A 58 3E D0 73 FC 74 C4 59 12 A3 B1 A8
 05 79 5E F8 4F 36 2C 2A B7 91 11 33 56 CF 09 16
 DB 6B 5E 4F DF 2E A4 52 65 79 CC B1 38 8C 00 71
 1C 81 84 58 58 03 E7 DE E1 31 EF 20 A9 8C 70 86
 44 53 63 2C 8A C2 E0 FE B4 8A 26 62 7D 60 E1 EF
 88 40 E4 91 5F F7 FB BE 42 9C 1C 56 BF 69 51 38
 05 77 1A 2D B0 5C DB 11 68 87 6C 3A 62 BB CD FC
 83 8A 22 BB 82 8F 22 50 AC C8 2D E9 58 73 4A 81
 40 E1 CF F1 54 C2 A1 FE D4 CE C2 F6 C6 9C 92 A7
 73 F1 80 0D 63 7E 93 53 7F 19 74 49 A6 49 44 EA
 E6 8A 1E 63 00 C6 7D 3A 39 AF C9 A9 F1 2D A7 2C
 DE 2A C0 D1 D5 FF A0 5F D0 E6 BF 99 35 13 A3 BD
 ED D3 C9 28 49 39 07 87 A4 5C ED AF 06 0E 44 D6
 0A B4 6A 95 44 6E D4 B6 68 E0 AB 72 8F EB F4 7F
 C5 B7 95 00 88 65 C5 71 A4 70 BB DC 1B 3A 79 05
 C0 CC AD 26 94 D2 E6 30 BE 65 2B 4D 0D AB 11 6B
 9B E4 A3 A7 C3 20 EE A7 9C 7D A7 10 6C D8 D8 19
 6E EA 5C EC F9 5C 44 D1 4E C4 D7 7D B4 50 BB 10
 1F 4C 01 C8 7D D5 06 D5 23 D5 EC 8D 58 F1 A5 09
 EB DF 96 31 50 D5 C6 86 92 35 4F CE FC DB AB D6
 93 EC AE C5 43 72 42 57 1C 02 4F 6F 37 FD 4D E0
 B4 45 14 EB AA EB 24 F9 7A 91 34 0C AA B4 E0 1A
 21 F1 6A 49 D7 B1 D5 17 9A 0A 8B C4 B1 E3 12 C3
 3C 29 10 25 41 BF 3B 13 96 7F 36 04 14 98 AF CA
 30 C2 5C 65 01 87 D8 C0 76 8D 7A 32 08 14 EE 1E
 FC 26 2E 20 61 C1 9A 5B 2D DC 22 0D 79 1E 88 44
 28 FC 65 0B B9 6C A4 83 DF 13 42 0B D4 7A FC BB
 BD B5 57 5D 4F 4D 0E 15 F9 94 34 30 13 21 55 9E
 59 D5 AA 9D 8E 4E 0A EF 93 39 4B CB 0E 68 2E 2D
 19 EE 1E C5 99 4E 61 BE DE 35 FC A2 4A DE 45 C8
 EA B2 40 72 C7 08 EF B9 01 CE F7 6C 46 8F 5B C9
 EC 94 FC 05 92 64 B4 BB CB 0B 1B 09 F6 63 2E BF
 FC 27 7A 6B B0 9F 18 4E F3 AD AA 31 20 AC E0 2F
 27 31 27 8A 63 0F AA 82 8F A9 E9 79 89 5E EA 5B
 AA 81 AA 56 75 33 C0 1B 70 68 B3 A9 87 4F 85 63
 22 F9 04 01 81 4E 6F 19 12 03 83 57 D7 C8 A5 64
 AD 58 B2 2D 8E 38 5F E4 D8 86 E7 3A 36 7E 74 FD
 95 CB 3F 99 58 71 8B 7B BD 66 FF 3E 8D 56 BD F4
 58 47 0A 82 4F 14 22 31 39 68 65 1E DD FD 4E 82
 F8 CF AF D2 EC 2E 04 BF F7 B2 1C C1 06 EA 86 C1
 AD E0 DA DF D7 69 C1 C7 8F AA A8 DB DD AE 6B 85
 E8 2B 05 B6 D6 D1 90 9F DE 9B AB 43 98 9C D6 F4
 87 3A 4B 57 81 9F A4 00 F6 5A 7F F1 B2 08 25 EE
 5C 00 4E 91 CF C2 F4 BC 94 3B CF C6 53 69 6C 7B
 3E 69 DB 4D 51 2A E2 48 98 E2 A9 42 69 7F BB 98
 04 B8 D3 1D 1E 63 38 21 9C BE EB 90 89 EB 50 E3
 A2 82 71 1A DC 2D E6 A8 C2 2F 95 79 A3 14 A4 C3
 10 69 6D 09 E3 61 35 E8 AE ED 44 D8 47 B7 0B 1A
 E3 61 4F 5E 55 52 78 9B 06 73 EE 48 BC 9C 1C AA
 A1 A9 F9 45 69 4F B2 A9 2B 0D 9A 9F 02 7B F1 5C
 A4 3B 1D 3E C5 25 C3 5B 63 65 48 56 A0 89 32 AC
 0C E5 ED 6E 5B DA 0F 43 2D 0D FB 6C 05 0F E2 65
 F8 58 15 CC BE F7 39 9F A5 14 C2 A0 BF 31 80 32
 FC 58 33 65 3C 0A 41 E1 B8 55 F4 70 C1 6F 85 5C
 8F 1B CD 9F F9 7F AB 4D 7A E7 81 EC A5 68 B1 7B
 8D 14 33 57 E8 52 02 CB 3F 56 B0 EF AF 08 F8 D8
 C8 AF 57 56 07 C7 FC FE 5E C6 6E B0 63 41 53 B8
 99 C0 BC F8 52 76 51 0D 77 A4 53 54 F8 D8 BA 36
 36 E8 9E C4 5D 7E 7D 0E 1F 06 1C 48 B0 78 1F 6E
 63 9D 09 8C 0C 6E A5 2C 87 C7 97 D3 FD 77 E7 0A
 0B 7D DD 59 93 17 27 CE DE C7 AC BE 0F 6D 7A 17
 5A 0F 8C 61 B1 A6 D4 78 B7 46 2B 1A C8 7B 5A BF
 C9 24 95 57 20 B6 80 38 52 C9 DE A5 CF 39 B6 40
 3A 63 37 05 6B 68 E6 05 92 68 4C D6 26 C1 25 9C
 DD F7 8D F9 66 02 93 3E EB 5E C8 78 FE 3B 1D 05
 C5 39 58 69 21 EC 22 56 AA 40 DF CD AB 37 41 5A
 58 E7 04 C0 E3 E5 93 B4 69 34 6B A6 DE D9 3D 9F
 5F DC 60 0D 73 39 47 B1 A4 36 05 A2 90 B6 D0 D2
 39 6C 20 ED 8C C3 45 18 AE C5 5A 9F 23 8A 33 7A
 66 3E D9 D7 D6 2F CD 8E 05 2B 80 47 0B C1 9D B0
 20 36 01 30 90 B6 DC 46 E2 1F C1 97 96 90 22 55
 86 35 88 21 59 FF 9B B5 B2 53 1C 07 D8 EB 5D 2D
 19 E4 C3 F8 55 CA 3C 8D F1 EA 69 8D 4A 55 06 0D
 4D A6 AC D4 AA D3 EE 74 4C F5 41 78 46 20 14 0D
 9A 0F 3D CC 75 45 0B F8 5A F7 2D 7B 5E C3 05 33
 A8 26 D0 FF 0D 18 A1 A2 B0 49 74 28 99 F9 E3 88
 C0 33 AD 2E F4 52 21 A3 37 38 22 C5 D6 F8 65 85
 5D CC 38 96 D0 78 B0 F3 3F 35 73 03 62 CC 39 F7
 32 68 23 15 1B D3 90 0A 02 02 76 FD 55 B7 06 AA
 0B CE A8 25 45 84 39 F5 46 17 8C 18 C6 E8 30 5E
 59 4A 67 FC 16 B6 13 98 0C 5B DD 55 F4 0A 53 B6
 9B 81 87 C9 A3 20 7E AF F7 4D CD B1 C5 CA 27 B4
 C1 BE 56 FC 86 43 5D BC 36 4B CD 52 32 DF 81 0F
 07 00 3E 3B 13 13 ED 87 56 1F F3 AE 97 D5 1A 7B
 1F E3 2D D4 E1 6E 8C 1F 11 01 89 F8 23 80 3B 4C
 38 4B AD 55 B0 2D B1 2B 1C 3B 43 75 E3 84 89 00
 A7 55 73 33 46 75 B0 48 26 A1 E1 D7 EF 8D FF 19
 0C FE 26 51 4C 3A 06 80 BD 54 A9 21 07 C6 B0 E0
 D3 67 99 DD 34 38 D2 5F E4 3E B7 45 F7 C6 AF 0C
 F1 E1 8D 62 BF 4F D9 AE 10 2A 32 83 E6 80 7E 7E
 39 B2 2A 80 A4 21 0E BD 69 92 A6 90 ED 21 0F BC
 7D 0C C9 AC E5 04 09 96 E3 7C 15 A1 A7 17 99 A4
 87 5E 5C 4B 90 A1 2D 2C 55 BF 15 1E B1 53 07 30
 EE BD E2 7F 41 1B A3 F4 10 13 D2 5F 25 5C BC A6
 51 18 48 25 97 3E 84 49 7B 34 6B 9A 43 F5 6B 34
 39 35 6E E3 32 A4 0D 41 1B 51 04 AB 95 E7 4D 07
 94 13 C1 3F 7B 45 F2 18 1B E6 91 D2 86 56 B3 0A
 EB 49 18 EC EC FB 9A BB 22 CC 24 8B 32 08 09 6A
 6B B7 37 86 14 9E 6B F2 32 A4 33 FD B3 33 89 FF
 E2 27 BC DA 5C 0D 86 F2 98 86 5B 06 AE 61 97 1D
 37 E7 68 FF A4 E3 93 95 FD 58 B5 89 7F 1F 18 A8
 0A CB 21 B3 B3 C9 45 01 90 42 BB 84 96 82 91 06
 86 1F B1 7B 9E CE 2F 2E E3 E1 4F B3 A6 02 88 61
 6D 33 7A CE 0B 95 77 A2 D5 0D F9 26 55 56 22 DE
 45 57 41 03 E4 13 02 E8 5C 9B 92 2D B6 69 2B 8F
 62 9C 1E D3 6D 0D A8 8B A1 B4 56 F6 2C 3C 90 D0
 2B 6D D6 AF D7 F5 9D 42 AD A8 52 0B EB 58 40 7A
 78 4B EA 97 AF 56 87 30 D8 41 9D C8 92 4A 90 6F
 95 1B D6 16 A7 22 2A 15 F3 8F 92 3C 95 5E E1 2A
 49 90 27 D2 F7 6C 18 18 63 75 73 E2 D5 BB 70 1B
 10 BA 0E 09 C4 A7 9A 72 E0 D0 95 AC D9 AC 3D 6A
 EE 5D 34 FA 27 84 71 BC 9A DE AC 4B 10 25 3D C8
 72 28 42 99 08 94 D3 23 E8 74 8F C3 49 14 E1 3D
 14 6F 79 1A 20 B8 53 6C 03 B5 D1 2C 93 31 7C D1
 46 5F 78 E3 D6 E9 A2 EB E8 05 21 CD 36 F9 C3 8D
 29 7B D9 23 27 1B AA CB D7 6B 2A DA E5 8D E1 BD
 B2 06 11 B8 F1 6E 3C 69 5C DD 07 7E 27 50 B3 C5
 8A 76 D5 9F 5A 9C 91 F3 2D 9A A1 44 AC 21 F5 FE
 CD 19 4F 96 95 8D E6 76 24 7D 33 D2 32 40 05 2E
 3F 86 A2 C8 20 7F 91 29 B6 13 10 25 48 D0 5B CB
 E7 9F 95 95 6B D9 52 A7 2E FB DD 56 85 B1 71 A1
 94 FB 9A 2A D9 05 A0 58 33 84 4E 7D 4D EA 69 EA
 30 31 52 B5 01 00 44 AE 73 AA 60 91 82 67 C7 A3
 E9 C0 E5 13 B3 2F 87 3E E5 F3 5B FD AB A6 F1 F5
 7D 3C EE 5E D7 23 63 09 16 0B 81 8A 1E 98 D2 D0
 98 D5 2E 4E 3E DD 74 D1 AE 89 92 64 0F DA F8 12
 C3 0F 6A 92 8D 13 22 63 F8 F7 B0 52 77 A6 77 B9
 E9 65 A9 50 7B F3 D4 86 6C 59 D6 7D E2 E6 31 6F
 70 52 3B 1C B2 E6 72 3B DD DD 2B FD DC 8D 04 84
 9A 24 3F 42 B1 8C FC 72 5F 8E BF E7 37 20 61 6A
 40 8F FF E5 92 9C 90 5D AA 3C 50 5B 86 E3 8A 73
 92 26 23 A2 4A 3C 07 93 B7 3E 86 33 4A A6 13 C4
 95 C5 F6 80 C8 2B 59 A5 EB AF 39 5D 8F 35 53 4A
 35 65 E2 88 64 1C 09 BF 60 51 11 51 22 D8 71 FC
 26 09 BD 26 98 F4 51 3B 0F C1 CE 0F 8E D5 05 75
 38 5E 7A 22 F5 25 DA 2D EE AA 0B CC 7E 9D 51 EA
 7B 49 5C 85 2D 4A A6 AA 82 D2 8C C2 90 58 16 85
 5A DB AC C2 57 05 66 06 A2 91 C3 CF 13 9D FF F4
 80 D7 D1 6D B9 48 EC 14 D9 38 61 38 20 90 AE 89
 8E 92 20 21 74 4D 4D 36 55 38 C1 1B B5 99 4F DD
 A7 5C 4A 04 48 85 B3 D7 30 3B 49 53 68 8E 46 79
 43 1A A8 B8 79 24 9E C6 74 71 1B 32 97 B1 5C 0F
 66 C4 FA C0 8D B2 88 D7 70 35 3C 85 85 83 E0 D7
 BF 66 97 25 AC 8A DE 64 F8 A5 B1 8A 16 EC 85 08
 AF 97 6D B7 B5 FF 12 63 FD 55 23 B3 F6 CF F9 3C
 A8 E0 D9 A8 85 BF BC FD 13 F7 09 C6 FB 32 90 80
 53 D2 BE 6A 1F 01 49 EC 66 BC 94 4C 71 05 E9 39
 3D 6E 1E DA 42 1F 53 89 AA 29 1E 2A 36 B8 E5 C5
 E4 6F CC 53 53 95 AF FD C5 9B 68 F9 92 BF 9B CE
 67 3F DC 7B DA C8 6F AB D9 81 85 A5 A6 AD BD A0
 0E F5 FF D4 BD EB 1B 9C 71 D5 17 10 89 BA 02 79
 F2 EE A7 7B B3 91 D1 A5 CA 23 37 B4 90 84 4D 20
 5E 54 98 14 7B FF 50 C0 85 20 6B 01 62 6C 84 90
 E7 1E CF 15 65 9C 1A 92 8C A6 E8 3C 1E C1 5B 2B
 68 D4 27 FF A7 EE B1 0E 83 3F 25 F6 4F 33 2B F4
 73 A8 7A 58 F5 CF CA B4 AE 77 6F B0 52 49 D0 41
 2A 08 7D 46 81 C7 6F FA BC 35 A8 22 23 C6 BB 27
 87 72 E1 B0 9E 82 E5 DE 45 79 50 AE D7 F7 A0 CA
 1C 08 1A 49 21 16 3E 17 76 52 41 7A 43 74 03 0E
 11 89 E1 73 7B F5 35 B7 9E 7B 4F E6 53 3C E7 D4
 07 48 65 B4 64 D5 C2 CF 06 D2 2F 39 82 E1 78 B3
 D3 F2 4C 44 06 EF 06 39 92 F7 CB 20 12 77 3F D4
 06 2D 3F 19 4C FD 26 55 5D 67 6D BA 4B 61 91 C5
 DF E6 C3 9E EB 35 54 B9 56 3A 30 DA E3 BF F9 A2
 C7 50 AE 13 EE 9D D3 8F 4E A4 A2 0D C4 2F 80 56
 D6 13 F2 BE 5D E9 EA D2 C5 67 E2 B5 E6 B9 56 DB
 D7 AC A2 2B 2F A8 A4 85 8E AA 74 88 49 F9 3F FF
 F9 B4 D2 F9 11 7F F0 EB 53 7D 8D 44 54 08 B4 F3
 25 43 48 0A AC 16 C7 B2 78 8F 0B 1D A7 B8 F6 C9
 23 C2 32 94 A0 D4 F6 C4 01 D8 67 E4 BD 7C D2 55
 40 2E CE A3 AF EF BB 77 52 63 10 52 13 3E A0 73
 DF 57 A8 67 E5 9D 98 F2 55 BC 68 86 81 7A B8 FF
 A3 55 02 37 FD DB D1 D5 05 18 C8 DC A4 8B 93 22
 BC 08 E5 14 14 0E 6C BF 05 BA 09 43 B5 C6 4B D8
 02 83 B6 61 4A C7 90 6E 37 37 A2 E9 37 4C 4A 65
 3C C5 98 5D DC 54 EB 73 83 B9 59 F4 21 1D 8D 57
 88 BE 01 59 80 2F A7 64 11 40 4E 50 BA CD 87 43
 15 B3 C8 7B 27 DE 43 6A BA 56 B6 76 FD 57 81 D2
 E7 90 66 87 3A 30 8C 95 8C 64 2C B0 33 07 A3 73
 A1 E4 E1 93 BA 85 23 91 0B C6 56 86 67 4E E8 3E
 27 50 03 C5 B6 85 6F 64 8C 38 C4 C2 3D 4B 11 66
 11 83 D7 54 9D C4 8D BB A5 D7 60 50 8B 8D AE AE
 D1 A6 D0 DC B4 58 FB 16 19 C0 CD C7 E7 18 74 3A
 C4 7D 01 03 7B B3 84 18 97 A3 1D B3 A8 D5 A4 82
 0F AF 08 5B 84 3F F6 B1 4B A6 A7 38 D3 1A 11 85
 7D 00 D8 8F CE 05 A1 1E EF 60 54 C3 FF 32 0F 48
 23 D7 91 50 F7 BC A2 01 73 8A EF A7 35 C1 5B FB
 BA B9 EA 1F CB 7C 08 E0 E4 90 6D F8 12 2C E4 34
 EB 09 5F 47 A5 2D E1 D1 07 3C 82 42 BE BA 58 C9
 31 7F 0A 46 23 7B 28 AC CC 0E D8 C5 DC 95 20 15
 F2 99 F8 19 0A 02 A6 68 15 0F 09 0A FC C9 A0 89
 6C 44 36 6D B7 1C 72 45 8C 94 F4 DD 72 40 9B F0
 7C CE 1A 38 C8 B7 AE E6 2D E5 2D 57 E6 68 D5 9F
 7F 73 37 66 E5 4D BA C4 40 5F 96 EB 1E 47 FB BC
 49 8D 66 F0 BB 0B 00 B8 3C 79 64 6C 4A D3 69 81
 81 9B 7D 4D 49 A4 45 8A 47 E3 EF 2E 4A 63 1E 6E
 A2 45 34 3E 0F 25 21 67 D4 8C 78 60 EB E0 C3 D9
 51 B1 E6 28 5F F3 94 B5 94 5A 5C 0F DB B3 6B 9C
 B8 6D 9A F0 44 17 43 C6 8B 42 3A 0F EF FD 59 5D
 51 B7 A9 30 72 8F 6B 42 65 16 CE 71 86 44 1F 9F
 6B 73 0E 3C CB FB 2A 57 4D 02 A1 3F 0B 9C 2B D4
 DB 90 BB E9 D2 DD AA DC B0 7D 1E 23 FB 60 0B E7
 11 60 2D 0D C9 02 5B AE 19 4D F2 4B 7B 59 F8 79
 C5 C2 4E 46 35 7D 9A 97 C4 6B 73 36 43 34 48 89
 BD 00 27 C5 90 C8 D7 96 48 E0 93 62 B2 38 62 EC
 12 C3 5B B7 59 DA 23 A6 16 FA 39 C7 1F EF 26 95
 F5 51 6E 5C 5E 87 4D 4E 38 48 85 49 5A D4 05 53
 58 A8 14 35 45 B3 69 B6 25 24 6D 48 F9 83 54 C5
 63 A0 8C B2 86 A8 63 7A ED 02 DA 78 5C A4 B1 E7
 92 C5 55 8A A3 09 39 CA 22 68 AF BE 72 2B 86 65
 60 80 8E 7F 12 FA 65 88 C3 01 EA E6 6F C2 C6 EE
 D2 E5 58 DA 2E 79 FF D1 25 18 00 85 A9 88 1D 0A
 97 50 2F E6 B3 99 35 0F 68 F9 A3 B2 AB A7 AD DF
 58 22 DD CC C2 4C 38 F6 DE 5F 2F 88 13 D6 24 2B
 CC EC 7C 4B 69 3C 2F 18 F8 BA 58 8F F6 D1 EA 7C
 4A 7A 06 EC C6 72 4F D8 E4 2C 7B 40 F0 F6 52 73
 7E 77 A3 29 C7 01 71 EB 8A 37 B5 08 EA D9 F1 3F
 C5 EE CB 49 B7 73 B4 06 CA F3 80 B0 AC F5 80 34
 BE 19 AC 97 46 40 00 8A F5 59 84 86 08 C8 03 6E
 EA F3 FF 87 48 C8 E5 0A D3 01 A0 0F 0F 05 34 F2
 63 2B 96 FE 57 07 6D FC 08 83 7D CE 01 D8 E1 24
 15 8A 99 4F 94 82 79 A5 6D E8 2F 0D 70 B6 FD 12
 D3 F5 91 47 D9 92 1A 19 87 82 23 A4 FC 9C 82 CF
 AE A6 48 77 52 43 3C 25 72 E7 68 E0 16 BE EA C6
 18 EF 53 FA FE 2B 30 BE E0 B0 D9 9E 29 33 E6 F4
 09 B4 D3 EF 0F 5C 3F B0 39 62 96 C3 1D 11 91 64
 21 CA 5D C7 28 C3 9D D3 30 CE 91 3C 05 A3 F7 FD
 E2 EB 78 09 6D BB 70 21 88 0F 1C DA 50 57 D1 D5
 F0 09 8C 9F B2 3D 99 0E BD 21 31 C7 5F CC C7 83
 E5 31 E9 B9 E0 3D 94 F9 DD C4 33 B1 C3 E2 C2 6A
 E7 56 E7 68 03 F2 91 04 97 47 31 DF 8E E0 80 34
 BB 9E CF 55 85 4B 70 F4 13 F1 97 13 79 54 31 54
 87 AA 1A 75 B3 59 04 14 AA D5 D0 E5 3A B2 60 7E
 0C E4 BD EB 9D CD 0F 6F 9F AC 2B 2B 6E 4A F9 82
 8B 64 85 76 8E 3D 62 7A 29 97 DB 0E 15 6B ED 2D
 B4 C9 7F 4E CE 47 A2 47 2B 02 52 D9 78 28 0F 38
 CA 83 A5 7A 21 4F FC 52 34 E8 9E 0D 71 E6 3D CF
 45 2C 13 28 08 26 C0 15 3E 30 0A EC D1 E2 94 52
 E9 82 59 5A 09 8E B4 92 ED C0 81 BD 46 6C 28 EE
 55 4C 1E 3B 07 23 EE A1 46 E2 31 10 97 E1 6F 47
 BE 6F 76 A8 91 42 48 A5 D9 A4 AE F8 67 F5 52 07
 3D 23 FF 49 92 D3 6F 35 B3 74 81 4A 40 F2 CF 17
 79 E9 33 61 9E 3A 7A 6E 6E 80 D5 C5 5C 75 55 3A
 53 49 B2 DC B4 C2 1D E5 1D 01 8E 57 6D 0D 79 1B
 10 8B 64 D3 6C FB E4 AB 0F 54 81 08 2E 74 0B 2F
 0F E5 3C 95 49 27 1D C4 2C 2D 3A 91 A1 89 F7 E9
 AB FC 36 69 36 E7 6D D0 36 A8 27 E4 73 87 E3 C1
 51 98 38 60 4F F9 2C 25 84 CE 38 93 53 E2 E7 17
 3F 1B A7 E9 D8 D7 F6 75 18 34 3A 96 67 BA CA 74
 01 24 63 2E 35 AA 27 DF 50 56 08 45 48 23 CA 64
 2B CF D0 D0 D4 09 95 0D 18 68 72 50 64 EA A0 E5
 D4 F8 E4 DE 5B 43 20 DE 8A 8B 00 98 4D A9 F5 14
 38 93 94 D0 52 C5 0F 2F C0 B0 BC EF 0F F3 C9 10
 0E EE 47 DC E0 9A 88 B9 A4 14 07 B1 47 8D 1C 9D
 5D 78 C8 F2 41 36 AE 04 91 C1 8A E1 6E D9 57 B7
 20 03 F1 86 BE D7 FC 02 F1 87 6B 6A D9 D0 71 AF
 17 35 5B 25 B4 B1 19 28 A0 49 58 5C CE EC E7 25
 17 B4 E8 4F E1 F2 80 D6 25 F7 B1 AC A6 A7 8D CF
 EA 01 9B 6D 4A 4E D9 A2 08 A8 46 93 51 4E 89 2A
 DB E4 C8 A3 0E 17 65 84 BC B2 55 B5 5F 87 C8 BE
 5D F0 E7 39 11 72 64 F8 86 30 57 84 9B BA 9D 0C
 D1 AB 8B 33 35 31 55 91 11 0D 74 E0 8A 4A E2 B3
 CE 2F 77 84 D6 15 84 F3 27 49 38 35 3E 1A 89 72
 38 BC 61 FC 44 6B EB 81 F9 FF BF C9 77 76 57 57
 E6 25 45 D9 0F E6 A1 8C 36 90 98 73 44 C5 6B C1
 23 E5 F8 81 7B 6E C1 0F CD 0F 37 D4 62 BE 21 9E
 76 AD 5E 14 D4 61 5D 0B 9A 44 89 DE 57 5A 0E E7
 1C 7B 5B B3 FE 16 EB F9 E4 9F CD 93 E2 27 D3 27
 69 D1 3E 07 36 5E A2 55 D1 DE 30 CD F9 84 16 C7
 F8 64 26 E4 23 9E 38 2C FB BD 28 47 92 6E 04 53
 85 45 9C 74 B9 80 0E 18 22 E7 D1 12 AD 1A 30 E6
 1C B4 01 73 14 72 2A 44 27 48 55 06 A2 E0 43 0C
 F3 96 6A 58 20 13 B9 A2 76 73 7C 83 81 52 C6 47
 9A B2 31 AD CB EE A0 8B 86 6B 32 3F 85 01 1A F4
 85 35 BB B6 F6 E7 D8 BD 78 92 41 6B F9 1A 38 1E
 C7 21 DC F8 13 F8 19 FB 57 D3 FD E6 B6 1B 94 F4
 5C CD 37 2E 33 6E AD 4F 59 6A 92 C4 B2 59 EB A8
 68 04 6B AB E0 AD 5D A1 BE 4B F7 8B 3B 76 8F AE
 84 0D 16 05 C1 07 D3 B6 58 09 28 50 3C 5B 6E 69
 AA 91 60 D3 AC E1 FB 49 3D B0 9F 0A 30 FE 56 6A
 92 4F B1 B2 17 42 B0 5A FC A1 D1 21 6D B8 AE E7
 9F 93 8E 63 94 9E 74 F5 99 A1 92 22 EA F0 16 63
 E0 3D EA 16 99 CD 8E 76 F6 7F FC 31 51 E9 A3 07
 09 05 AB 0E EE DD 4C BF BF 3A BA 76 8F 96 A7 7A
 01 DC 48 7A 54 B3 91 BE C2 F2 EC 41 C8 60 05 DD
 A5 37 54 58 6D 52 EE DA 7E A9 4C A8 EF 02 00 FD
 0E C7 2A C2 7A 9C 4B F6 42 6F 70 2C 14 13 D3 2E
 1B 6A 96 B1 21 5E 41 FE 7D 92 D6 84 CA 3C 42 24
 A5 DE 40 DD C1 ED E6 52 32 1D 02 8F 78 8F 7B 19
 F5 99 AF C5 E5 B1 F0 67 3A 7F 04 00 01 E5 D5 B0
 54 07 A5 AE CD 1A 3A CE AF 83 D1 E9 CE FD 9E 91
 CA A7 CA F8 3A 8F 20 3E 50 D5 FF A4 B8 88 FE DE
 29 7D 30 51 33 B8 FE B4 23 B1 4A 71 D5 9F 8C 34
 B6 79 E3 DD D7 51 5D 8F 57 7E E3 96 5F 79 E3 75
 1D 3E 89 22 93 18 D5 61 7C 7A 3F B9 98 64 0D 57
 F6 8D 71 C4 42 8F F9 EF 06 23 DC 0E BF 85 AD 8F
 F5 A4 1D AD F7 F9 D4 90 4B C9 7C CA 5C 02 D2 C0
 D5 D0 F0 EF 5D 46 9A E9 3E F4 56 E5 97 CB D0 BB
 6E 58 CB 3B 60 46 E1 31 52 2F FA 8E F7 DE DD 34
 C9 9F A7 2A AA F2 FF 5C ED E8 85 8E 66 F8 08 A6
 2E CB B2 91 8A E0 8F 63 91 30 1E E4 CE 1D D4 B3
 2C 31 A8 A4 0B 33 0D C0 8D D6 AF EC 93 33 5E E5
 49 58 27 74 61 19 DD 66 8A 7E CC 9C 21 C6 61 37
 4B D9 60 ED 8E 02 93 A5 E4 5F 8E 59 A1 96 11 18
 9A 10 17 D2 E4 C7 AD 2B 49 CB D0 63 A4 3A 2A 0F
 4C F2 FE 59 C3 2A F3 38 11 F1 54 62 4A 16 53 D7
 8D 47 5C 91 25 6E BC EC 75 97 AE D0 85 27 14 2E
 5F DA 1B 53 50 22 81 90 8F 91 56 5D 3B 9E 19 A3
 7E D5 9A 64 63 7A C2 97 37 B3 28 00 32 9A E0 D7
 E2 22 2A E3 01 25 A9 6C 72 90 A9 CB 70 E9 4D 27
 16 CC 86 39 D3 8E CB 1A 8F FB E1 56 23 2E 20 FE
 F2 32 F7 06 DF 19 0E 02 94 79 17 7E 7D 97 67 D1
 E5 56 A3 C4 9D D4 A3 2F 69 E9 9E 54 84 B7 32 12
 89 78 F0 05 BF 03 7B 74 A7 20 A4 DF 30 12 86 0E
 36 B4 FD E5 C2 43 62 DD 03 E2 A0 1F F8 10 E5 E3
 D3 B3 82 57 B4 F7 AE 46 6E 29 C5 A1 6F C3 E5 49
 0A 49 91 57 35 AA 39 02 2E 09 5A 4E 9C F3 A2 29
 64 3D 90 FD 79 C0 81 10 B5 A0 A1 51 0D 83 E4 47
 EF 6A 92 F9 D9 E9 0E FA C7 DE EE 50 8C F1 A8 CB
 E7 DD 8D 15 4A 42 38 8D F6 F9 D3 29 B3 27 38 B2
 63 46 5C BB 9B 89 34 71 93 A7 79 00 D7 A8 77 67
 A3 B7 CB 94 2C C7 2D 88 F3 FB EE 1F 5B 56 76 86
 3B 09 6A D6 FD 63 E4 84 79 0D 62 05 B5 10 F0 88
 29 62 F7 E8 78 F5 9E E2 49 95 1B 62 E9 02 7D 97
 DE 56 A9 34 9C 30 06 59 31 FC 1B 5E F1 3C 90 9F
 62 26 C5 B3 BD C4 36 7F BF 8D 39 BF 74 E5 22 A8
 7A 1F 15 39 8C FC AE F9 61 CA 78 60 E1 27 AA 1F
 93 B5 1E B6 48 0E D0 A2 8C 2D 89 17 E8 58 1F 78
 80 23 C4 E7 CC 1E 5D 01 08 FE 53 54 B2 AE D4 E6
 7B E4 D5 F8 EA 1B 1F 22 F2 D9 E3 4A A9 B1 42 12
 B4 49 81 69 42 76 B9 FE FF C5 62 18 E1 20 0F CD
 6B 98 3B C6 C0 59 F0 45 02 DD 0E 4E 4B 78 14 B6
 A6 5F 0C 35 AB 41 82 17 04 22 CF 00 19 1A 40 42
 4A 0F 05 89 7F 2B EF 48 70 2B F6 FD 38 5A B9 9F
 59 BD A1 6C 61 4E 4C 82 A3 16 E3 6C 0C BD 6C 58
 AE 2C 5B 32 86 89 A0 38 D2 78 D3 1D 1C 5E 6E BD
 1F D8 A3 7B A9 AB 26 9C 91 B5 F5 B2 0F D5 59 8D
 DD 35 E9 95 E1 C6 2B 88 4F 8E A7 30 F0 89 47 9A
 D1 A7 41 D0 0E 9D 74 33 6D 67 10 68 CA 43 FA 85
 59 51 AD E5 C0 7A 46 CE 9D 49 FB 0B 93 64 DE 0A
 3D 52 D5 29 75 BB 02 17 00 91 F4 B4 23 EB 62 5B
 1A CC A7 5E 38 1A 61 7C B3 97 B3 0A 3D DB BA 15
 22 CD 3E 54 2C CB 5E 65 5B 4E 32 13 34 BE AE 94
 7C 70 D0 0E BC B1 E7 95 BA E7 55 BA 7D 97 06 44
 91 5C 37 8C D4 28 0F 09 AB 69 1E 9C 8C 08 FA C7
 E4 5F 1A 86 2D C6 D9 F9 CB 5C 56 E4 0A 52 C6 C3
 19 9D 92 6D A5 0D F1 6E 3C 13 FC 00 7B C8 E1 E2
 49 47 47 51 BF 99 7E 21 AC 1B 6C 1E D2 C6 E0 E4
 82 EB A2 9E A7 74 E0 18 EE 6E F4 41 46 36 8B C8
 A8 D8 3B BA 98 97 03 26 92 A6 A1 80 0C C8 0E 0C
 7C C9 28 34 DA 44 2C FE FD AD BC 2E EF E5 A3 55
 4E 73 35 49 FF 75 04 19 51 8C 85 CB B3 0D E9 2D
 D2 B7 8F B1 8D 18 15 A6 56 1A CA 63 3C 2B 3C 39
 67 94 38 D0 19 70 60 55 1D 0B B9 55 D1 55 F0 56
 45 9B 57 39 9C 63 B1 42 CC 05 15 20 D1 2A 04 77
 5C CE D4 40 80 1D 22 D2 33 9C B1 EA CB A0 42 67
 B6 AE 7C 84 64 9A 30 EC 7E 7E 05 86 E7 CB DA 22
 A5 A7 F5 D2 E9 21 33 58 70 76 F3 76 C4 C9 99 0D
 D3 6D 41 B6 05 AC 18 48 5D 27 0F 7D 07 C3 BA A6
 BF 68 D5 F1 4A C6 74 07 41 EA 8E 4E 6A EF 35 69
 CB A0 76 23 37 65 65 E8 CE 5C FF C3 41 37 CB 88
 69 46 F0 40 AF AA BD F2 73 D5 CF 97 8B 94 42 49
 20 C3 CE 50 DE A2 13 9D 01 56 91 81 4C 0C C7 6F
 36 CC 59 8A D1 AA CC 78 AE 63 D9 AA 0E 41 63 38
 20 E9 30 40 45 47 7B B9 43 F6 54 40 0E 82 30 25
 DB 67 EF 25 73 14 63 1D 24 7B F7 BF E9 6E 3A 36
 C5 3D 08 A8 54 1C D7 B5 5C AF 65 B3 BC 96 53 F5
 96 8B 99 2E 36 03 F2 8F 14 80 E8 2F E1 D9 B0 4F
 81 05 41 BE E6 3C 1F 78 91 24 A6 85 BE 5D 82 EC
 4F 97 43 DC EB F0 65 0B D0 01 5F C9 E1 DD B5 32
 A5 2A 85 DE 66 D0 4D 22 BC 74 59 7A E6 29 00 99
 42 F9 D1 9A 38 CF D0 65 91 EE 05 E0 60 7F 97 C9
 A8 29 69 C5 09 CE 1C 1B 99 DF 35 77 70 4C B6 72
 DF 7B E8 31 D6 E0 3C E4 DE C7 49 B7 D8 A9 04 CB
 05 6E 2C 49 F4 58 A5 B5 DE B4 F6 B1 7F DF 0B 92
 3A 15 69 05 F0 6E AF F6 3C 60 44 A0 AC E6 07 43
 93 B5 49 69 22 5F BE 08 AB A2 8D 9F 16 A9 F0 90
 CA 38 3E E4 A3 A6 50 C6 9E 88 C8 27 61 52 67 BA
 69 41 B4 CC 4E 58 53 2B F0 C3 51 A3 0A 0D AB D2
 3A B3 33 3D 61 AE 34 C1 77 4D 0D 44 8C 80 C8 80
 ED 02 97 85 15 C6 94 D8 6F 31 7B F2 57 29 AA 29
 FE 45 CC AC F7 F0 A5 04 3A 70 43 8A 38 C8 E8 00
 3D BB E8 95 EA A1 4F A2 FB 6F 64 15 A5 15 AB 6D
 AD 47 AD A3 69 57 C3 33 FE CA 5F 9B A3 74 4B 9F
 AF B9 57 F3 A3 FA 7A 06 0B 8D E5 10 25 F1 35 B2
 62 9F 92 04 44 E9 84 2A BE 06 20 42 35 0F 19 F2
 6B A1 2A 03 83 31 EA 4D E9 98 81 94 D4 AA E5 22
 7C AD 26 3F B1 8E AE 17 EA D6 F5 7A 02 21 0D 8C
 1E 88 EE 19 57 D0 EE 89 D9 A6 4E AE C0 3C 63 40
 F9 23 09 FC 20 92 DD 66 2D B4 0A B7 49 85 C6 85
 75 84 7E F5 06 67 0E B9 1B 36 72 3A D4 C0 6E F6
 81 EE DA 72 35 87 43 CD 86 24 7D 12 C4 4B 31 A4
 58 0E E0 60 80 53 AE B2 B5 20 5F C1 42 EE EE E3
 33 78 A3 8C 2C 94 47 76 4B 4D 04 E0 FD 26 15 E2
 8D F4 87 5C 7E 28 F2 49 E8 0C 38 BB A2 16 18 06
 A4 3F CC 71 22 1A 27 89 E9 83 D3 5E BD 01 1E 59
 F0 EB 9F C0 37 49 67 DD D6 1B C8 A8 00 F9 8E 56
 AC DE 25 04 AD BD 64 6C 14 7D 86 D7 60 21 E4 E0
 0E 1D 36 51 8B 2D 28 06 D3 84 DD 43 9D 07 CA 01
 92 2B 1F F4 76 73 D4 25 FD E3 37 F2 9C 1B 79 CA
 72 69 B1 1D FA F6 85 0E 26 9D 12 E3 61 4A E8 CE
 36 CE 04 18 93 BD 96 46 73 AF 6C 56 40 9E 0E 9D
 C6 D9 D5 2B B5 3B 62 C7 22 2E BE 5B FC 81 D2 22
 83 C5 3F 70 2B A5 18 70 26 41 C6 B0 FD 34 B3 02
 42 B9 78 C7 87 E7 14 2B 7A 44 FD BB E6 E9 84 50
 86 24 8B 8E 69 54 BF 21 CF FF B6 45 AD 6B E4 65
 2B FB 04 A4 30 37 A7 E6 B6 45 2B B3 4D CF 3F 1F
 67 7C 80 F1 3E 6B 08 D6 3E 97 EB CD FA DF 91 1F
 45 C8 65 28 6C E1 05 17 2A D5 69 28 C3 C0 06 FD
 85 22 CD 1F F2 F3 6D 4B 77 F6 16 E1 DB 00 D5 BC
 C6 91 B6 28 38 F8 6C 6C F3 B3 CA 5E 27 CF 0A AA
 41 FA D8 FB 99 C1 71 C7 A8 18 1D EA 21 E6 BF 43
 C1 F7 51 CF 2C B0 AC D1 EA 06 32 72 64 B3 5D D5
 EA 41 F7 EC C6 53 80 F5 29 A5 8E E9 22 1D A4 51
 96 63 B1 C8 6C 3B 72 F3 C4 85 CC 3C 61 C2 9D 18
 66 23 D8 80 3B CE BA D6 91 63 CC 05 E4 6B 53 86
 31 E8 39 D9 E3 D5 A7 73 EF 14 CF 32 DB 0D 17 5E
 54 A7 BD E1 4D 4D DD 73 E3 D0 2C BD 0E 5B FB A1
 12 9E B4 19 FF 42 AB 63 9F D5 4D 55 AE EE A6 7C
 F0 54 8A 8D 0C D8 78 51 C5 3E F5 FD BE 1E 70 FA
 CB 67 CF 0C 7C 0C BE 3A EA 98 A4 52 35 BA F3 FF
 55 B1 18 A9 E1 F4 B3 46 2F D0 3F D9 8C 02 CA 9D
 54 76 90 05 E1 92 F9 80 65 E9 8F 2D E3 8E D9 C7
 A6 3E 35 DF 28 AE 66 E0 32 42 11 8C E1 0B 89 1F
 86 F5 71 B9 EE 72 20 37 61 78 2B 88 48 34 70 90
 44 A9 67 A0 CB BB 3B F8 3D 63 E9 D8 53 50 6F 19
 84 56 57 C0 6D B0 2A CA 99 D1 30 78 C0 04 DD 24
 7F 8B 99 0C 7F 6C 4B 05 57 89 CE 57 65 F8 55 00
 6C F2 4A EF F7 D8 0B FA A8 CE 8B 0A 62 91 89 85
 B1 D3 5F 2F 51 C4 D9 48 2B 98 31 B6 AB 2F A7 50
 71 66 92 7C 8E 33 2F 35 6E 33 E4 0C 9A 4C DF 93
 E7 70 E6 F9 9D F6 50 D6 5A FB 7F 19 CF CB F3 80
 13 ED C2 FA 45 96 E8 13 8F 53 EA DF 51 C0 B6 EC
 00 16 47 08 3F 71 63 29 11 23 A5 7A 78 B4 B5 C7
 0B 47 B3 C6 B0 E3 D2 54 A4 C3 DC E9 F2 06 27 01
 FB 49 FD 28 0B AC CD 35 FA 5A 25 A1 F6 65 30 52
 62 2A A1 4E 85 BD E4 EB CE FA F0 75 D2 3A 96 18
 AA 8B 52 E2 6A 39 28 2E 8A F1 8C 51 CA C9 9B E3
 CB C6 BD CA 4B AE B1 04 3A 77 DB C4 97 FA BC 1A
 2E C1 F2 F1 0D 53 F9 71 A7 8C 29 95 66 52 D1 B9
 50 54 3C AB 71 31 E4 A8 D7 70 A2 DD 4A 4B C8 91
 D7 F3 3E 87 6E BB EE 88 7D 2B C4 D9 40 29 03 7E
 BE 87 0B 2D 59 5C 03 91 B2 84 C4 13 76 70 D2 C7
 B2 2A A0 B1 93 BE 14 35 C3 85 45 DA 37 55 FD FB
 39 67 E4 D9 50 58 EA 19 4B 23 D8 CC DB E8 02 69
 A5 8D BD 1D 63 9E 88 72 4D E9 62 A1 C9 9A 7B 09
 27 5E BF 45 9D FF 37 6F 0F 8E 15 44 C1 7C F8 4F
 8C 25 2D 98 AA 1C 97 2F 4C 8C D0 39 EC D9 D9 F8
 1E 8F D4 40 3C A2 9F 5B CE CA 1E A0 71 9C D6 06
 6F 71 59 73 A3 85 E1 6C AD 7E 70 91 CD 4F B1 57
 AA 08 5F 4E B9 8A 60 A0 FB 68 30 93 21 E4 68 94
 7A A3 C2 69 BB 7E CE 15 EA B2 78 24 21 3C 12 61
 39 C9 CC 0D 11 4E 3D B9 99 1A 4D A4 47 7C 6A 5E
 EB E2 F2 5B 75 94 21 E5 B0 18 3B C0 E5 74 75 0E
 E3 49 98 A6 C6 0D 4B 87 0F 69 4B D9 A5 EE D0 80
 1B 8D CC FD D9 38 CE 82 5F D9 13 03 9D 2E 93 15
 B7 28 54 BF 23 29 D1 BE 07 9A 0F 6E FA E8 62 CF
 C4 C3 15 27 F6 0E 18 FB 10 6C 24 43 62 DF BB 54
 A5 B7 AD 79 39 B2 AF 42 0E 57 55 A9 03 CF 78 28
 80 29 6D BB 10 72 9D 90 3E 63 65 9E 3B 7E 91 DA
 3A 34 D5 29 E4 6C 5D 99 E4 C1 65 01 96 07 77 CE
 11 B7 29 47 C4 66 12 0F 08 CA 94 8A 1D 50 FA DF
 C0 7C 9C 1D DC F0 6B 4E B7 B6 0F 11 26 75 EC EB
 69 E4 B3 31 6E 51 36 B7 11 C0 AA 38 BE 56 B4 4A
 6B CA CA 6E FE 27 C4 08 DD AD D5 80 3C FF 84 AF
 61 E1 26 56 93 76 C0 25 2A 26 72 F9 7B B9 92 0F
 E7 ED 3D 2D F0 76 4A 40 D0 89 37 8E 81 5F B5 DC
 97 D8 62 C0 D9 32 34 8A D5 22 5D 4D 07 46 83 21
 70 5C 91 8C EE 3F AE 26 D4 E9 20 CE 63 D2 60 42
 A2 80 FF 8F BB 49 46 F3 DF 71 49 D3 AD 82 98 5B
 60 F9 52 44 C1 DB 39 9C B4 72 CB 2F 58 71 D4 C8
 FF 93 71 01 D0 B0 D0 72 9E 19 0C F7 51 32 B8 F5
 39 7D 8C 78 E1 B2 F1 77 B4 1A F1 03 30 AE 9C C6
 1A 5B 56 5B 3D 79 01 02 B8 BC 2D 9A 68 B9 33 FB
 DE A9 30 C4 B1 30 0F 91 AF B1 5B D5 3C 24 7A 71
 06 F7 45 AD 28 ED 5C E8 64 B2 B5 9A 22 10 FF 81
 D0 D5 55 58 96 B0 02 F2 15 06 83 FB F3 80 68 E6
 EC C0 2E BD 23 C1 AA 40 FD 56 D4 A6 2C 67 13 FC
 0B 6F 97 C2 2B 18 2D 69 17 B8 AA B8 18 FE F4 3B
 9D FB C1 DC A0 69 AB 3C B4 D4 A6 61 63 0E 53 49
 1C 23 6D 4B AC 35 F3 63 B4 CF 6F 77 FF D4 CB 87
 5C 82 20 FF 67 0C 20 B1 EF 77 C1 DD 6F 30 E9 3F
 E7 17 E7 33 35 1B 06 1D 8A 40 F5 FA 0C 14 8F 04
 30 4E 61 75 CA FE E4 98 22 9F 06 84 58 09 B8 3C
 95 9E EC 00 B4 43 27 F3 0A B1 31 4D 8C 8F 6B 4C
 71 CE 95 15 AF FA E9 50 5F 51 2C DA 1F 3F 85 92
 D5 44 AE 99 E4 38 31 D6 2D BC F7 CF 66 F8 E2 D9
 52 F2 10 D2 A8 14 A7 BD 7B 7D 41 0C 0A 00 D5 0B
 8B 58 AD 6A 33 2A 6C FD 7A 9E 6F C9 C0 05 F2 14
 22 89 BF C4 93 0E EE 0D 5D F6 B5 5D 72 F6 BA 74
 71 5C 82 A6 80 54 EA D2 D6 D6 4A DC 82 26 F5 C7
 B8 BA A8 97 BB 11 E2 34 76 06 F5 89 E3 8A FA A4
 24 5B 29 59 FC 0E D5 E5 D7 21 B0 D2 51 2A 83 68
 05 08 59 2D 22 CD 40 31 9D 29 E4 3A 41 E6 BA C7
 D8 5A 21 08 D6 A0 A7 C6 CE 65 80 7E E3 13 EA 08
 69 D4 95 AE 93 FF 89 7E AC 63 2F BD F2 1B F3 E3
 63 B5 15 39 75 C1 07 B8 41 CD CB 54 FA 2F 7F 04
 03 09 51 62 5B F0 84 E6 7D 1C 8B 69 BD CA 45 B2
 1E 62 A5 07 99 DD 88 40 80 B1 AC EE 48 D8 93 9C
 43 E1 5E BC AD 54 A3 00 8A 15 6F 14 68 82 C0 21
 AC 4D D4 B3 7F E0 6A 40 DB 75 65 C2 11 2A EB FD
 FB 32 D8 EE 71 FE 4B A3 48 6A 2F E7 30 D3 BC 4B
 4A D3 03 A7 11 DF D7 E6 D3 1B 23 30 CD F8 BC 19
 B4 51 F4 05 D1 77 C3 8A BE C9 3C E4 E3 B4 CE 94
 D7 44 5E 43 3B C5 95 82 80 FC D5 1B B4 08 A2 FF
 1F C5 D9 23 DE 2B 28 06 EF FB 7B 8A 4A 3D 8A C8
 B7 69 A3 1E AA 20 FA 8E 16 F0 21 49 54 6F C2 20
 18 84 F9 3F 89 80 CA D9 90 D3 74 69 FA 2A 94 33
 51 8C E8 7D C0 DB 51 D6 E4 96 DA 94 7F 52 14 13
 3E E5 45 AE E3 32 B0 CD 15 C5 DE 73 EC 37 11 97
 6C 20 6F 9B D6 BC 87 65 B9 B9 31 2A C0 33 0E D6
 C3 DE DD 5D FD 98 C8 82 90 C9 8E 2D D8 41 59 20
 95 F6 72 0E 47 ED FB FE C2 9B 1F 65 95 F6 AD B0
 30 6E 01 C6 30 32 5B 0B AA A5 59 54 B1 D3 DC 03
 E4 95 63 CA 7D 62 AD 76 48 68 76 A7 17 E5 DB 40
 C8 FC AC BF 7A D5 7D CF 40 07 C7 01 19 6F 6C ED
 1A 71 58 C5 0B AD 5A 76 93 9E 08 BE 8E 8C 8E FE
 4B 94 1C F5 10 84 C6 F1 91 9D 58 47 C4 83 01 C4
 5D 0C A3 07 60 4C 24 4D A0 30 F7 03 59 56 5D 70
 EC 65 BF 96 AD 06 E5 42 88 E1 B1 A9 A8 EE 9E 03
 BF 19 88 91 B6 61 16 59 71 C1 15 1E C6 20 26 4E
 FE 48 C2 AE DF 62 C1 20 60 A6 06 C1 AC 42 16 7F
 AE F8 5A A4 FC 68 3C CE 95 25 4E 73 DD 1F 28 56
 12 52 24 81 CC 8C 08 C9 4B 86 08 CA 6E CE 43 96
 F7 A2 5D 19 DB 55 BB CF 3A C4 F9 36 1B E1 E6 3B
 BC 7A 2E 96 89 35 8A 71 1A 4C 8C 63 72 F3 9F D6
 7F 97 0B 52 2B E2 F2 B7 8F 46 61 2E 84 3E B3 13
 EF 7A 58 BA D2 0A 36 CE 8E 89 7E 0E AF FA 38 FC
 92 FC 88 E8 87 66 73 07 39 52 32 57 12 17 EC 4E
 B7 A3 8F FE AF 85 44 9F 1E AB D6 15 8A 53 16 F7
 CB E2 88 51 81 15 72 A1 AD 61 1B E0 E2 EB 51 DD
 47 54 83 C3 7E 65 F2 91 21 7D 23 12 43 D1 3E 3D
 42 26 EB B9 7F 06 0C AA CF 37 06 1A 89 FC D9 97
 2E A0 1E B3 38 55 99 50 ED 4D 8B 28 C1 7C E4 F7
 F2 FE F5 B2 2C 6F D4 7F 35 BC B2 64 AF 56 B8 A9
 0C EC 75 93 95 F4 23 BB 84 A2 C0 27 2E 89 DB 15
 C2 DA 0D 76 7B E1 01 BA 5B F7 ED 4D BD 3E CD 15
 F2 CB 98 38 12 81 41 E4 2E F1 B3 31 7D CD 54 07
 89 0D 36 AB 1D 8A C6 F3 8F C3 61 15 A8 90 06 38
 D4 50 89 6B BC A5 C8 F1 E8 26 EA 63 0B 33 25 72
 64 56 16 0C A8 CB 1F 11 F8 B7 27 85 81 1C 15 C3
 6C DC 39 90 7E A1 57 3C B9 44 85 9E 91 77 5B E6
 7C E5 64 B0 62 34 CA 4C ED A4 7E 49 A9 DE 94 04
 9A 22 B8 1A A9 D3 54 67 4F C4 C7 0A E7 C6 09 E6
 F9 57 2D 75 AD 65 32 28 30 74 E3 B1 3A 6F FD D2
 1E DB 51 13 1E C3 40 52 83 BA E6 AD F7 61 F5 07
 BB D2 F0 76 AE D5 5D EB 1E 2D 9E 7F D8 AC 3C 95
 F5 37 75 D3 EC 2B 09 F8 EA 25 B2 14 0D 3B 08 0C
 E0 D6 36 85 16 9A C4 29 66 77 D9 C1 AA 6D F2 7F
 7E 22 5E 98 F8 9A A5 02 BB F9 37 98 02 EA 6E B9
 60 DC C2 B9 56 A6 45 A3 1B 05 1C B2 B5 C4 E1 79
 24 26 A8 9B 4C D0 CE 77 AA 4D E9 62 6A F9 44 ED
 F5 D2 9D F6 7F 13 01 39 DF 29 D3 FC D0 A1 C4 1E
 26 C4 9D 7D 96 DB CE 1F DC D8 7D 8D AD 83 8F 33
 A2 82 BF 3A 19 5D E1 01 77 98 72 7D 95 74 3C D0
 11 12 56 83 2E DD 21 D6 2D 92 ED 63 E1 F6 47 2F
 09 59 25 F1 97 0D 84 DA 44 06 B4 0F CD 51 F2 11
 2C 9E 46 F8 9F 96 08 64 E3 7A 20 09 67 67 33 7A
 27 39 35 C6 C1 35 12 D9 15 6D 07 9D 85 30 4C F5
 C9 39 B0 A7 FB F5 4B F9 3D 60 AF 34 3B B1 CC 44
 BF 81 CD 98 23 90 17 16 47 47 10 5E FB 00 A8 B8
 21 00 68 72 D2 A5 E8 E6 45 62 8E 07 A3 A3 93 68
 69 74 84 EC 8D 37 E2 10 61 CB FA 4A 1A CF F5 DB
 51 53 91 05 72 89 87 E7 35 5A 5A 89 7D B3 E4 A4
 63 76 88 1F 56 D7 5D 76 0D 2C 8A 17 9B 30 69 7B
 68 DA 50 10 2D 27 27 78 B4 C1 1C FA 0B B7 C4 1D
 D9 D5 BF 75 77 BD 3A 26 90 4E C2 60 94 0E 49 30
 68 F7 9E DC 45 3A 86 36 C4 5C 59 3E C2 16 E1 F6
 3C 59 96 75 E6 47 17 10 CC 73 93 0A 72 32 9D 1C
 66 04 42 F4 8A 00 B7 6C A6 BD EE E0 30 A4 DF 41
 01 F4 AF DE 3D 47 D2 44 B2 81 0D 6F 7B 89 2A 90
 73 5D BC 67 2E BD C7 9E 1F D5 7F 1A 70 3F 63 13
 5D A0 FB F1 F4 B8 7F 50 23 62 4F 3E 80 3B 48 01
 93 EB 72 51 BC F9 89 E8 5B 58 03 BF 4C E5 61 40
 34 82 40 B4 1B 2A 68 46 E7 6E 53 F4 85 96 09 5B
 74 87 51 93 E3 6D 6D C6 CC A5 00 D2 E1 DE 89 5D
 B7 BB 14 D6 37 53 9A D6 F0 77 07 2C 5A 09 AF 0C
 85 59 9A B7 26 5C 46 D1 29 3D C4 4B E5 A8 54 BD
 E5 19 E0 25 1D E4 D0 5E 24 B7 5C AA C5 18 27 6A
 75 80 27 7B 19 CA E9 86 B7 A7 75 F8 37 95 B7 EB
 EA 59 F1 F7 1D AD BC 50 EC 86 E9 87 A5 75 1B 0F
 F3 59 2D 1D 2B 13 E7 8A 32 AC A4 9D 07 D9 5B 45
 A6 81 35 4E 2C 02 1D 9A E9 55 60 E3 A4 BF B2 0F
 F3 51 ED 51 6B D5 33 CA 4D 30 97 B1 FC A9 37 AA
 A4 CA 6D CE 28 C0 13 29 F7 27 CE B3 3C D5 2C E4
 C5 5D C7 9D 12 5D 37 AA 0C 1E 49 25 78 90 1B F7
 73 79 C7 83 47 59 FB 6A CA 31 DF 3E 34 1D 4F 1F
 C1 28 3E 78 08 49 E6 E3 53 BB FC 01 70 05 78 92
 27 67 33 7E E0 D1 88 10 91 DF 2F 1D 1B 7A 5E 84
 77 54 ED A5 75 80 1D F6 6C 07 83 50 20 E9 0F DE
 10 7B B0 9E CF D8 EF D5 80 5E DA DD 8F 2E E2 6F
 C5 04 96 DF 4F 84 32 2D DE A0 3A ED 03 AB EB FE
 57 6B 4B 1F D2 EE 70 11 D6 C2 E3 A5 04 9E 4B 22
 56 1B B0 C8 C0 5E 45 8E 88 B8 CC 5B 0C 68 AE 1E
 3F F7 8B 3B 2E DA CB ED E2 1B 07 D1 DD 9B DA 80
 59 31 33 CA 3A 71 71 43 27 28 94 CF D8 64 D6 57
 C5 89 ED 5A 53 1C E8 DA E0 5D 81 93 12 E8 90 BA
 81 D0 7E 25 3D F0 AC 8A 36 FF 6C C1 B1 7C F0 24
 2E 56 B2 A6 0E EF 52 75 E0 75 F8 EB 8A A8 BE 71
 45 A1 6A 8D 20 C9 92 11 E0 CA 92 55 BB 34 DA B2
 29 BF 9D B5 AE D6 F8 9A EC 50 9A 78 9C AD E6 24
 8D C7 10 C2 2C D5 ED C2 0B DA F3 BC 88 DA 20 56
 6D B6 78 DC 86 61 00 79 A9 C0 CA 89 E7 F8 AC 03
 3B 71 34 B6 E9 7C C4 E1 EF 40 0D 5C E2 F0 A4 87
 E6 2A B0 D8 68 C4 2B D5 7C C6 6C C7 97 7A 4C A5
 9A 72 B0 15 D7 26 CC D4 3E DE A1 F8 9C A9 37 6A
 45 A5 74 00 3B C4 4A 9F F8 38 0B 52 53 40 62 0E
 D6 9E 03 11 FF 79 7C A9 DA 74 AC D3 28 8E 93 6B
 3E C9 18 D9 19 B2 72 1F 9C 76 58 AB D5 6E EC 20
 E2 87 71 87 81 61 71 72 18 F1 68 84 47 3C EC A3
 CF AC 06 55 FF 8B 55 DF ED 7E 08 EA 8D E4 02 B9
 44 3F 93 2F F4 F4 AD 1A BC 88 4E 91 59 35 3D E8
 58 EB BC 16 76 C3 C4 CE 08 22 32 3E 17 A1 EA C1
 E2 B6 F3 BC 6F 1D 22 87 AE D9 FD AB 72 00 DE 4F
 C4 2C 19 30 FA 23 BD 51 67 4E 34 02 CA 63 04 F4
 25 39 4D FB 51 E9 3C BB A2 03 67 00 5D 56 5B 32
 4A 3E 63 8B 1D EF 20 71 02 28 F9 B2 81 9E 13 02
 42 D7 EC F8 04 B2 29 9C A7 DC 9D 59 CC 4F B8 FC
 47 FB 2D EB 7D 5E B4 33 74 68 CF B0 96 D7 FD 14
 04 24 25 4D DD 2F 12 EF EC 7C 5D E7 C3 E6 88 16
 35 3D 19 D4 26 02 63 BA 74 62 F1 B6 73 54 59 87
 78 3E A0 55 70 59 D9 3B 60 90 59 30 0E D6 DD B6
 A2 6E 63 7B BE 7A E9 3A 35 74 F9 E4 7E 25 E4 AC
 B6 45 40 84 41 A2 53 11 80 DC 58 BB BD D7 3D 38
 1C BE 51 21 C7 58 BA E6 A2 F3 1C 65 A7 42 0A 4C
 82 9E 2B 5E 6C AF 12 41 BC B7 93 01 B0 C3 F0 AC
 F2 D1 7A 42 AE 49 8D B4 21 A3 8F F6 74 12 FF 29
 BF 60 62 56 6B 14 1F F8 AB A9 7D 1F 91 4A 62 CE
 EB 00 A5 F2 49 6C 89 64 46 12 DF B2 A2 59 E0 6B
 3C 17 F0 D6 C4 41 06 44 92 A2 14 08 E3 B0 1F F1
 2E A3 8D 96 20 17 D7 30 21 26 B1 92 3C 72 5A 01
 B1 31 89 B8 1D 6F 6F 39 12 2F 6B 22 DE 78 D8 86
 7F 5B 5F 31 E9 5B 95 62 16 00 26 AB 42 07 A8 25
 E6 5A 8F E3 E3 03 DA D1 DB CE 94 89 F8 FF C2 83
 E0 A6 53 3D 33 3D A7 6C D4 21 25 5A F3 B6 A4 B0
 CB F3 29 89 56 72 C2 15 2A 1C C6 A3 0A 9E 93 AF
 55 4C 2C 40 57 27 FC 09 91 D8 A3 27 35 F2 82 B3
 93 9F 46 BB 5C FE 23 32 94 71 5B 58 7B 96 91 0B
 ED 6A 1B 00 9C CE 81 27 8F C8 C7 B8 8C FC A1 19
 5A D1 F8 D4 1E A5 58 D7 5A 8C 4D 89 DA 9D 5A 24
 2A 28 35 32 C9 15 93 B9 62 FE 3E 07 80 71 2B 93
 08 B5 0D FF 63 16 87 56 DD A1 FC 01 54 9C 2A 0B
 F3 D4 2B 10 8D CC 0F 3F ED A0 78 DF 68 A3 EA 98
 4A 19 05 B2 45 4C 6C 47 20 00 A3 86 68 49 69 71
 C9 E5 32 1B 9B 9E 39 4B AF 5A 50 DF 95 4A B7 EA
 9F 2A 70 3B 0F 97 6B 94 CD 6E B2 A6 07 B9 5B E0
 6E CB 47 F4 84 71 45 29 2E 50 85 F3 81 BA 12 F6
 57 29 40 E9 EE D2 30 6B 64 86 D8 53 72 6B 10 2A
 03 4C 67 1A C0 32 FA 33 67 02 F4 88 49 7F 20 3D
 B4 F0 63 92 20 33 50 02 E1 41 3D CD 08 B2 5E 34
 B0 99 C6 CD C1 0A 28 43 74 39 99 C9 F1 83 23 37
 3F 64 13 BF C0 0B 4B C3 66 11 69 78 0C F7 72 4E
 25 7D 40 39 78 F3 B4 5A C0 3D CB 62 41 60 8D CD
 8E 9A 6E 21 31 16 E5 E0 13 AF 49 92 0C 1A EB F2
 05 84 5C F1 16 8D 98 62 11 5D F0 0D 03 E8 9B F0
 52 9E 82 BF 70 42 23 7F E1 D9 81 0A CF D4 B7 81
 36 E8 BC 2A D5 BE 08 F0 E0 C6 BC C5 24 46 60 93
 2B 2E DC FE C2 1F 2F 69 68 02 58 6D 9E FC FE 2D
 E0 A2 05 6D 3F FA 58 1F 1B 3A 19 CB 5E 40 49 A9
 C6 74 AC 1F BD 2E FC FA A0 33 84 DA 19 60 6D B2
 C1 E9 25 35 0F 29 34 82 9E D2 64 F5 88 C5 38 43
 ED 9E CE 83 B7 B2 A0 4F 93 B1 BB 6F BE 6C 82 D9
 97 D5 F5 05 C1 E2 B5 F3 B5 31 9F 2B BE E1 E8 9F
 B4 C1 55 62 80 9A AB 5C 62 F9 B6 80 6E 5C C5 15
 2B 2A C3 5A ED 1C EA F0 90 21 52 61 BA 4A 5D 12
 8C 5F 94 0A BC D9 D0 59 77 10 6F 0F 1F C7 1C 36
 6C EA AC D8 9F 31 F6 01 91 F0 4F 3E 1E 49 B3 0C
 42 5C 1A BA 6F 21 28 EC D9 F7 51 76 6F C5 AE 3F
 62 24 33 B3 41 F4 DF D4 F5 2B 81 C1 DF 0F 4D EA
 5B 26 D8 96 4A 99 D4 08 34 DB 16 79 F2 0B B0 56
 90 84 CD 99 F1 BC 33 48 6D A7 DE B3 0E 84 ED 56
 E3 E9 A2 75 BA 21 E8 30 63 E4 55 3D FB EE 46 31
 B5 29 9E 29 AD 21 E4 23 93 2B 68 66 45 D8 76 A6
 B7 58 4F D5 EC D0 6C C3 E6 CE 5C F4 6C 92 6B 12
 FE B3 99 CF FE E2 37 53 77 F0 6F B3 62 63 C8 13
 6D A2 65 C7 A1 72 FC D5 39 DF 5D BD BA 2E D2 80
 F0 24 28 27 0E 76 31 D2 EB 29 AD 58 A3 9E AA C4
 26 42 BE 2F 4A FE 33 3F C8 E9 9D 44 7B 76 07 E3
 F8 3C F6 F3 E7 68 CA BC DA 53 67 C0 67 55 B7 C9
 F1 62 CE 48 B7 1C D3 B6 9F F6 A1 7E F9 89 C4 D7
 8A A2 9B 11 9A FC F0 A5 75 E8 C3 DB BD FE AC 96
 10 AE 8F 99 75 81 47 AF 52 F2 58 4E F7 27 0B 53
 92 ED B9 8B 59 BC 31 EC 7E 11 17 AB 6A 83 5C CF
 27 7D 3E 3B 6D 65 03 1B 46 DC 1C 97 7C 83 44 82
 D7 C3 F5 BB 44 3D 87 7D 22 83 BA 57 B7 35 68 FD
 AF 01 3E D2 98 8A 26 7D 85 39 8B FE DE 72 3C C0
 0E ED 0D 40 59 3B 9D 9B BC 84 36 03 27 B6 D5 48
 AB DB FB C5 D4 6B C0 FD 03 64 F5 D3 13 BE 13 50
 C8 AC 59 B4 C3 D9 09 B0 6F E9 A8 13 54 9F 4C 14
 AC E2 E6 BD 15 DC AC EF F7 D7 50 37 4B B8 06 7D
 1A 90 63 DD 9F 12 BD 41 70 B4 33 E0 11 18 5F 9E
 66 E0 AD A5 BE F5 C0 05 DE 55 AE 75 AF B2 39 BA
 16 0C B8 36 6D 03 5F 54 F5 D0 CA 2B B4 94 15 D4
 82 CA AA 84 E7 E1 5C 7F C4 AB F9 7B 22 BE F9 67
 61 73 34 4E 63 DA 9E 7B ED C9 8B 98 97 32 4C 8F
 9C ED 82 67 B3 2D 15 A5 1A 0D 5B 1F 91 C5 70 B1
 A3 99 AB E2 60 BC D9 4F 16 C7 53 41 1E BF 52 D5
 E2 49 AB 8B 52 C0 A5 F4 FF 56 12 76 78 81 D7 FA
 DD 60 6A 16 21 91 46 A0 FE DE 6B BB C8 B7 D5 EA
 72 30 E6 9F A9 F6 B4 AA 23 E6 1C BE 3B EA BC 08
 0C 1A C2 C6 6F 76 08 5F 8D DC 16 3F DA 6B 00 36
 E2 47 F0 A0 B9 C3 A3 39 B5 61 58 1F CA DC DE 6F
 2D 61 CC 20 87 B6 38 78 2A ED B5 53 72 31 89 6C
 2D 7C ED 02 7D 05 49 BB 43 BC F0 6F 7A E4 E2 FE
 3F 26 62 62 B9 91 46 22 5C 60 9C 67 1E C6 C2 31
 A3 01 E6 E5 CA 26 A1 8D 1D 47 C3 39 F2 3B FD F5
 E5 40 1E 87 80 38 BE 68 F7 28 29 C7 62 6A D7 9B
 0E C7 EF 87 61 C8 CD 66 A9 AA 57 E1 CB 24 6D 18
 78 9F 17 8B AD 14 57 2A 00 0C 25 B9 B7 C7 2E 1D
 8C 4A 08 B9 D7 FB 8E 6C ED 26 20 F8 4B A0 E1 CD
 68 CB 39 C1 F1 5E EA 37 C7 15 94 2D 9D 9C DB C9
 EB BF D5 D4 0C B2 E9 A5 69 48 40 4B 1D 70 DD 68
 52 BA 96 FF 04 10 5D 67 4E 1C 2E 5E DD B6 5E BD
 52 7A 8E B8 A9 2C 1C 24 DD 48 7E 1A C9 68 EE 2D
 E2 89 A2 5F 02 5A 19 04 CE D4 54 AD E1 5B FA 78
 45 2D 8A 4A 06 B0 FB 70 62 81 57 B1 E8 87 E1 36
 08 5A BC C3 58 AC 25 95 67 D4 A5 A9 71 21 35 62
 6F B5 F7 F7 3F 00 EC 48 F9 15 3D 0A 12 FF 5F CF
 6E F4 C7 53 1C 9F 96 09 70 FF 97 1F 8B 80 02 82
 95 3D D3 A2 31 8B E3 2A EA 4E E0 32 93 34 19 E6
 82 D1 DF 7D FB 52 3B 15 18 C6 3F C9 BC 0C 54 39
 85 11 24 FB 5A C9 57 1E E0 E1 D4 72 AA 7A 1C 7F
 00 D2 56 13 9B 63 42 D4 64 30 06 DA 95 08 A8 7C
 70 28 C4 03 1E 78 75 D0 34 47 8D 9D A8 2E DF 2D
 83 11 6E DD D4 1E D9 CC 79 75 74 31 7B 96 6F 57
 C3 06 58 80 BD 77 75 A1 A0 08 0A 83 21 79 DB 0A
 A1 97 A9 FC 2A 41 01 4A 81 CB 5B 08 F7 3F 3C 9E
 65 1F 96 E4 42 E4 F0 5B 14 F9 0D 8A B9 1A B0 87
 56 62 91 16 82 77 55 C9 E4 7E 6B 9E 58 55 13 BE
 F2 BD 9B 4C 2F E2 FC 59 44 80 38 18 DF F4 A5 91
 6D 45 8F CC 33 2B 17 D5 7D 6A 71 EE 4C EB 1F FD
 76 23 59 26 86 F3 D3 6A 4A 8E 5B 94 EE 90 D6 75
 1E 89 34 9A 0D 12 B1 C3 C2 F9 68 1B 66 0F 6A 3A
 B7 E2 04 BC 27 E8 CF FF 8E E2 17 7B FF 3C 40 EA
 81 84 D6 A4 52 5D 71 34 42 44 CA AE 71 B5 5E AB
 2B 63 EC D3 78 DE 1E CC 12 8D 7A 3B A2 2B CF 91
 A0 41 50 07 4E 75 40 72 1A 7B 09 33 6C 52 46 06
 87 D6 4B F9 BC 3E 5A 08 AB A7 FF 0C 4C 6F 19 29
 93 9B B5 E2 DA 56 E8 65 A8 BC 6E FB 90 55 2D AB
 80 12 0A 1C DF 00 F7 5F 22 6D 14 DE 33 EE 7E 05
 68 AA A7 72 38 48 AF 43 2D 45 3B E8 80 1D B6 9F
 5B 86 83 85 57 C7 CE 5D 29 53 37 99 0F B4 FF 95
 5A 1B F1 6E 6D 54 C5 0E C3 94 96 49 56 55 B9 36
 F6 F9 27 76 5E 9E DA F8 F4 27 AC BD 65 33 74 A5
 85 D9 90 A9 38 1E 40 52 31 59 E4 BC B5 4C 19 E4
 6B 24 17 08 3B 95 B5 62 6C 54 4B C4 B1 6F CA B6
 9C 10 ED DD 3F 74 6B ED B2 5C E6 59 40 D3 A1 38
 24 41 03 64 3F A4 0B DF 58 C4 45 B6 C4 7F FB 86
 7C CD 44 69 FF 90 8C E5 53 3E 2C 73 27 72 E8 FF
 C9 48 2C C1 85 C8 7F 4B 86 93 B5 4C 90 57 12 93
 E6 0A 6E 88 CE 0A 70 5D B7 FD 86 38 13 AE 3A BB
 05 A8 2C F0 55 56 4B 5A 22 82 05 85 54 B2 55 8D
 F5 C5 01 AF 78 4A CA 0E B4 6D 96 DE 75 0A 1E 39
 BD 78 E5 F0 50 05 7E 28 98 AD 6B 14 F9 C9 7B 51
 FB 47 98 FA B6 57 3F 4C FA 8D CD A5 18 E4 75 ED
 49 3F 13 F5 43 FF EA 04 91 D8 05 A6 65 64 55 FB
 06 BF 57 72 7B 52 DF 68 59 C1 C0 17 E7 8B E8 25
 4F 7A 87 8A 75 8A 74 D0 D8 11 A6 21 17 DD 10 3E
 EF 60 32 7B 22 D6 EE 2A F7 19 61 E3 1C AD DA AF
 1F 45 3F D3 AB 55 A2 36 F2 C8 31 82 8A 05 2A 93
 75 F3 EF A8 99 87 64 40 04 8C D5 04 DD B2 13 C9
 64 C9 4F 58 C3 8D 03 28 36 F6 54 C9 63 85 2A 2F
 25 AB E2 83 66 E6 5F 74 5B 7E E5 0B 68 4D BF BB
 45 DC 2D 21 F8 FD 81 11 82 2A 5E DD 96 A8 BB 72
 06 ED 07 13 C0 C3 F1 E6 D4 AD E7 E1 4E A5 0F 09
 2E 11 81 6F CA 75 85 45 00 56 64 FB 5B 04 53 4A
 F9 3C A8 5F F6 DC DC 36 2F 94 E0 95 CC 8C F3 AF
 06 4E D0 EF 8C 9A 00 30 3A 3C EE 0B D1 AE 32 E0
 8C 31 DD E5 F2 2E 76 65 87 AF 17 B3 E2 42 84 82
 74 CB CD A0 22 5C 00 C9 C8 9B 03 5C E0 E3 89 23
 14 D6 BB AA 69 D0 30 F1 E3 18 42 48 88 FB 23 63
 FE A7 1A 40 54 FC 7C 9F 3F 5C 0F 12 67 4A 3E 01
 1B E0 FD 6F 66 80 3A A3 69 52 5A 42 C2 74 EE 34
 C7 A8 2B B7 2D 64 47 5F DD 68 F1 8A AB 07 E9 F9
 5B 7C FE E2 A0 A6 39 95 B3 5E 67 E6 5C 53 22 EA
 08 62 6A 1E D7 0D A2 66 AB E2 DA 58 05 8A 4F 75
 EE 3C DA 4F 91 68 F3 A0 F8 B4 73 7A 54 1F 81 A1
 96 5A BB D0 91 90 D4 5D 15 A2 2A BC 68 B6 29 7A
 32 9F 45 9D FF C3 6E F2 90 15 A9 6D 4F 28 12 8B
 7B C3 43 8E 5A 5C A2 99 59 C2 8F B9 E3 E9 29 36
 64 03 8A C9 4C F8 60 D9 0D E6 D9 84 64 E4 C1 F7
 A3 51 2B FE C9 4D E6 B1 A1 F0 13 2F D8 7A 90 79
 4E 2E 27 2C 0A 82 B8 5F 39 0A 86 61 AD A4 CB BC
 D9 36 7B C4 01 30 F4 6C BC 8B BE 83 2C 15 C8 B1
 2C 14 05 F5 DF D3 6F EA AF 89 B2 B5 7A 3C 65 30
 B5 61 16 C8 09 07 9B FF 8D 28 A6 43 C9 4A 47 74
 06 9E 6D 68 C2 D9 4F F8 5C 28 9E A7 21 10 13 8E
 9D 85 6C 71 C7 A6 0D DA 4C CF 6E 3A B3 8D 37 CF
 EA FA C6 E0 36 8F 53 BC 70 8B BF 5B 82 11 47 52
 02 85 64 A2 21 2E 35 31 FC FD 16 72 71 C3 9C 14
 62 5F 13 DE AB B0 DF 3A F6 89 58 12 F4 4E 96 FA
 B8 A1 C8 52 E0 99 E4 11 34 9A 6D 26 0C 71 4A 2D
 EA E4 BA 76 DB CC C5 3D B0 BC 4E A4 B9 32 51 69
 37 63 AE 86 70 EB 0C E6 9A 64 76 72 AA C1 5F 71
 7E 46 20 8D 70 35 73 27 6E 37 F9 C0 24 5A A4 4C
 B4 30 9E EC 25 D7 DA DF A1 FB D1 ED 16 98 6C 89
 13 EF 73 78 93 45 EB A8 12 A7 87 C9 81 5F B2 F0
 CC 28 30 46 D1 75 ED C6 9E AE F1 FE 12 BE 5B EC
 EC C2 C2 79 F6 BD 5E 91 35 92 8A FD D6 29 71 37
 C7 8B C1 46 66 95 BC 77 93 B8 9E 63 56 27 3F 46
 2D 53 C3 38 30 ED EC 1A E8 35 35 EF 6C 58 70 29
 87 D4 BB 07 1F A3 4C 2C F0 43 45 75 92 55 44 83
 59 81 D0 14 D6 D7 14 9E 94 AC 0A DB E2 84 6C BB
 E5 59 C5 89 2D F7 AC B3 EA 85 1A 91 67 CF 63 0F
 A0 FB 2D C1 FD DE F2 17 B0 68 D3 EE 59 16 EE C8
 98 71 F5 B2 D3 8C 0B 9C D5 F0 0B F2 8F BA 5E C6
 FC 6D 68 77 04 09 79 41 C8 8F 3B D8 BF 3D 51 B5
 51 71 3D CD 5E 1D FE 1C 79 30 BD B3 F7 9C 8D 43
 31 1A AB C5 0E D3 CB 50 BE 1A ED C8 CA 6F D6 71
 AC 09 D7 24 8C E3 B5 4C 9C F5 FF DF FD 0D B1 B8
 31 B4 08 A6 7E 7B 6E 36 4B 7C 77 4B 60 74 9B E8
 0C 29 E8 A9 53 A6 CA 21 BD AE 1D 1D 47 0B A8 64
 CB 09 33 66 5B 14 BE FF 6D EB A9 9F 66 99 3C A1
 F7 04 85 09 5D BF F6 75 EF F7 21 0F 31 3B 26 66
 E8 E4 48 1D 3A 93 D3 E6 07 31 44 2B 5C 95 7B DC
 B5 EA D9 E5 0D 03 D3 37 25 3E AF 40 79 35 A2 9B
 D8 24 E1 FB 3B E3 2E E3 5E 45 90 B3 42 74 E8 96
 87 12 57 19 BD 7D 04 FC 9B 1A 84 F6 AE 7A A7 C7
 FB F7 50 73 D8 2F FB C6 E6 2E 2E C9 2C 86 EE 3E
 5D DF 7F AA BE C7 36 55 A5 6F C9 A4 B3 AA F1 BA
 29 23 D0 C4 8B C7 FA 38 C1 64 45 6C 80 91 33 B9
 94 0B 28 10 4B D8 9A 0D F4 B3 8C 92 5D 0D ED 4C
 50 47 73 95 9D 38 30 21 46 15 0F B7 93 97 2E DA
 B7 F5 2F 1F E0 5B 6D 6F CA A8 5B DC CD 98 D7 EC
 08 87 E6 F3 47 C1 65 A0 01 D8 E2 2A 6C 0D C0 07
 7F 47 09 4F 5B 40 4A 1C 85 3F 5F FC 8F 5C 68 A6
 96 36 4D E7 4D 2A 00 1A 94 95 F8 D5 5D 04 B6 05
 49 FB ED 08 AC C1 6C F5 75 96 98 59 2B 62 19 F5
 0B AA B6 CA 56 01 6A 7C 6F 34 E7 FB 5D 49 1B 56
 D7 5E 8A 36 61 15 52 B4 31 D1 E0 12 90 4C A5 4B
 A5 CB 8F 99 1F 85 4D 1E EF BA B3 93 3B C8 0D 02
 73 75 1D 5F B4 EE 60 F5 3E E9 80 15 76 3D 56 27
 7F BD 0A 32 31 61 B3 9E CC 3F C7 11 94 56 69 11
 3D E8 E9 92 83 07 F9 FD 28 73 F8 3D AF 56 3C 64
 33 EB FD A6 F5 81 8E C4 4E 87 D8 B9 F6 5B FF F6
 D4 21 B3 BA 52 D9 5A E8 D1 D4 79 BE D2 82 05 2F
 32 63 58 95 8C 97 79 AB 29 DE 82 DD C8 7B EA 0A
 9B 89 FC 9C 8E 34 88 13 BC 60 82 76 69 BA 72 1B
 CD F5 B5 69 36 F5 A5 A5 5C 22 48 84 BA 95 65 4E
 5C FA B5 94 52 A4 F8 F5 06 EB 08 39 17 B1 E9 FA
 66 63 B5 79 75 C4 E9 64 AA 97 CD C9 AB 33 16 8F
 23 34 FC 64 97 F0 B7 28 16 5A E0 A5 01 5F 8B 98
 47 36 B2 CC 81 4D 57 00 D6 92 5A C5 92 F7 C5 D4
 CA 5E 04 04 DE E7 79 4D 29 48 55 DE 8D DB 6B 43
 F9 E4 6A 5C 07 A3 EE 82 CA F8 31 E1 22 FD D9 30
 38 EC 6E 11 68 90 58 82 FD 33 19 D6 C8 05 5B C2
 F0 D7 2F 26 74 EB FB C5 1D DE 7A 58 AB 64 A5 32
 FE DE 1A E6 2B 95 ED 9D A6 79 4C 68 0C E6 BF 58
 91 F5 4A 07 84 03 16 97 93 68 5C FA 06 E7 9D 52
 94 23 E1 4C EF 23 68 C9 8C B0 16 80 F8 75 53 95
 05 34 DD 26 54 5D 5D 14 48 22 C9 6C D0 31 7F EB
 0F 8E 93 A3 75 84 7D 34 2B C5 69 CB 54 F8 6E 30
 9A D5 80 F9 76 5F 39 DC F9 DC E3 C5 1B 3A AE F9
 54 4E A4 EF 5F 19 23 74 58 ED 78 FC E0 B3 CC 06
 1E 36 13 DD 3A C0 98 7E 81 BC 62 2B A7 B8 D2 6E
 20 5B C6 8A 5B E8 1A 4A D0 3E DF 27 FD 9C D7 E5
 69 CF 50 A8 37 5C 50 23 7B 89 21 E9 5F 8C F8 F6
 D1 09 45 D9 5A 8F 91 03 BE 6F 4B C1 CD 26 E2 71
 46 F6 D7 13 CE 54 B1 02 10 88 8E 2D 87 84 ED C6
 C3 D9 05 DD 49 35 73 D5 FC 78 C3 20 92 D3 B0 19
 C3 59 CB A3 F5 C7 1E 62 F2 E7 9D 29 D0 D4 B2 F1
 A0 C2 FA 9E F6 4C 29 B5 3C D5 15 35 A1 11 BF 02
 27 68 BB 4D 8B F7 7B 0B 5A A6 19 A0 5D 9B AF 5C
 76 41 1A 70 01 32 00 CA 81 56 DB 72 AE 79 84 63
 C6 AD D3 0A E5 CE BA 07 BD 0A 34 8B B0 50 77 E0
 A8 E1 A4 A2 3C 63 BE 50 6F D6 C0 7A 1B B1 0B 51
 CB A8 AF 4F 3F 56 25 8D 6A 73 5E 67 1A B8 3E 57
 96 E8 74 E4 73 CC 53 E7 D7 3B F9 3D B4 57 5F 6E
 F1 E6 83 2C DE D5 F4 41 58 12 22 C5 D8 98 74 91
 94 0F CE 5F 6B A3 63 A4 DB 26 1F 0D 51 5C 09 78
 E9 94 C8 25 0D C6 AD C6 1D 05 BA 82 2B CE 14 AC
 35 1D 51 0B 61 9E D8 88 79 69 7D 6E 93 71 6C 46
 75 3D F5 57 32 52 67 0B 87 58 80 5A CA 56 DA 1D
 4F C5 28 5C F3 86 53 74 40 92 75 DB DC 9A 19 8E
 36 66 09 89 B6 8E 18 74 6F 24 3D 73 30 7A 61 1A
 FE 3C 7C C5 8C 00 5F B9 A7 C0 4B 93 5F CA B7 3F
 ED 24 D0 52 F3 66 06 2B 41 39 CA 35 EB 18 5B D6
 62 EB 11 E1 8D 3D 56 62 82 7E C4 3E C3 3C 5A 7E
 52 B5 16 FB 36 82 FF 34 29 FC F3 B4 DC 67 91 5E
 46 21 11 B1 54 8D C1 D5 42 94 64 DA 40 9E 70 0A
 42 A6 4F 5E AD D0 0B CD 1F CF 13 4F 79 4E F1 A7
 C9 C1 79 9E 20 49 A6 DD 2A 85 FA F7 9C 03 D4 95
 F8 6E 95 10 97 D7 20 85 20 62 2B 28 1A 08 A8 06
 B1 56 E1 E5 43 91 A8 00 E8 AA 1C 62 D2 0E F9 BB
 70 3B 97 8A 68 70 2C 77 7C E6 51 66 09 FD 65 9B
 C1 1D 2F 10 46 CB 68 10 3C CA 89 FD C2 A2 F3 DC
 D0 ED C4 DE FE 07 FC 01 51 A7 24 CD 0E A2 EC E3
 19 75 4C BE BA CC 6E EE C1 57 96 B7 67 D3 5B 3F
 96 D5 19 9F C9 72 E1 B7 0A BC CF 82 6A 62 A7 2B
 6E 1B D3 D1 89 56 A5 AA 00 F3 91 0A 79 F1 44 5D
 F9 0C 9D D5 D2 3B 28 EC D3 E4 9A 3B C8 E4 7E 96
 24 D7 44 5E CA D0 71 3F E3 11 72 84 63 F4 76 23
 D5 35 ED F4 22 BC B9 A2 94 B2 09 7C DB 57 2C 52
 77 2D 62 E6 B4 F2 79 11 4B 76 0E 8C 1C 6A 0C 39
 1E 48 7C 62 81 49 91 BF 27 3C 01 2C 5A 2C D5 E5
 DD 2F C6 06 D4 E8 89 4D 23 93 66 85 1F E5 6A 55
 2A 15 BF AB BF 38 94 29 EF 7E D0 D1 B5 4D 63 BC
 AF 14 EC 33 1B 45 F1 64 C1 EA 33 D3 00 6E A2 09
 F0 32 BA 3A FB 20 CC 70 60 B0 AE DF 97 50 84 6B
 27 30 08 51 54 15 09 30 4D 8F 99 23 61 EF 62 A4
 BE FE 21 80 78 A9 54 48 51 8A CA AB 75 F6 7B 14
 39 94 BC 09 5E 64 7C CC DB 0A 79 A7 B3 EB 32 20
 CE BF 53 45 4C B9 C0 95 41 C7 AF CA C3 60 FC 9D
 98 11 C5 F8 E4 4A 40 0F 76 D7 34 C8 4B B8 51 FB
 0D E7 8C 56 3A 85 DE 2C C8 D1 F9 DA 9C 68 AB 8A
 FE 10 83 24 2C AB A9 01 A6 DB 3B 64 F8 B4 F5 01
 B2 47 D0 96 39 CB F7 A6 26 0B E5 E0 4A 5F 2F F0
 17 C0 BD 19 39 55 09 B2 F1 7C 5F 02 0B 3F 7B 15
 C5 70 50 45 03 4D 65 06 23 90 CF E3 F6 38 8E A0
 75 17 3E 45 3B C9 54 9D 14 3F 38 25 A5 22 9B 13
 7A 6F 6E 16 62 AA 18 D0 68 5F F5 83 12 54 AD DF
 BB B9 7A B1 D6 88 4B C7 05 36 9A E1 38 66 1C AF
 02 03 2E B1 15 9C AD 3D 85 5B F1 D0 8C 5C 51 55
 11 2E 48 67 FF F9 15 68 40 FC E8 D1 BC EB 93 71
 B4 7F E2 4A A0 E2 A0 8D 00 43 A1 3E 42 FE 7F 9A
 67 85 BE 8D 8D 44 6C 7B B6 A9 6F 11 1D 25 59 D5
 11 D8 42 84 41 D9 0D 28 07 6C 72 69 52 6C BC 2F
 48 46 87 97 DB 30 73 F2 AC 20 A5 AD 4A 31 1A D6
 A1 F2 15 F2 C0 4F 36 AB CF 13 EF 1D F5 6C F7 BB
 07 BA 81 7D 9A 4F 4F DC CC 95 8A 74 F6 A1 AD 78
 CD BA 8A 90 EA 98 83 E2 FA 68 B0 DE 0A 48 E0 A1
 A7 6D E2 53 0D 67 CA 61 C9 AA 0F 09 97 89 C1 ED
 14 E7 BB 93 5A 6F 42 AD 2C 77 69 77 84 96 3A 92
 87 F3 DA 53 8D 65 02 E0 0B B6 90 97 3C BD 54 B9
 6E D6 3B D3 41 0E 00 4D B7 F6 12 8A BD FE 09 33
 33 3F 77 F4 42 E1 2D 0E D0 AD F5 1B 35 A0 52 12
 76 5E CB B4 67 4C B7 3B 11 ED 1D 05 6D 1C 15 16
 BF 70 45 9D 91 F3 E5 D8 78 9E 09 A5 BF 3C EF 3C
 12 63 A7 B3 1F 9A D2 98 79 74 F8 7B F2 7F BF 6F
 E9 C2 E1 11 90 93 51 65 59 4A D9 14 71 0E D3 C5
 C8 B2 94 C8 09 F4 D1 85 EF 2E 4A E7 CC CF 91 B3
 67 FB 58 92 A4 93 AE 52 05 76 E3 C3 87 94 F0 94
 69 52 EA E7 D6 40 89 CB AC F9 4A A0 C4 D5 72 44
 DA 22 AA 11 A1 11 4D DF E1 5C 40 7C C4 52 90 1A
 E6 85 F2 BD 39 03 55 FD 8D A7 46 D1 5B 2B B4 35
 64 EC 45 E2 53 A9 57 A5 1D C2 CA 00 46 B3 E2 7B
 10 DD EF 9D 8F 1D C0 4A A6 E0 18 24 C9 1C A7 A1
 95 12 CE 5E 56 9B C1 F0 AC 53 FE 41 9B EA 0F 46
 DD 3D 7A 6A 19 AB 55 95 E2 E9 C4 CD 69 0F F8 0C
 DE 41 D7 52 F9 42 EB 2C 52 51 64 C6 B5 D3 C1 79
 90 33 45 4B 4D 3E B2 77 9B 8D 52 F9 46 FB B3 E5
 BD 46 A4 FF 8B ED A8 E7 DC A2 00 11 D0 92 3B 79
 11 AC 20 FA 6B 0E CF EB 94 20 8A C2 EF 7B 2E 52
 30 56 1F AD 8C 1E B3 83 61 13 FA 2F F9 76 0A E7
 01 5C 19 28 B8 D4 41 F5 89 C6 5C 29 A0 17 AA 26
 01 30 50 BE 13 14 54 39 CB 5C A3 09 83 04 80 1A
 02 C0 16 7D D0 4A FE BE A2 5E 9C 06 2C 10 A5 49
 A9 C4 CB DC 5C 0F FE 8B 01 38 44 F4 98 6A 3E 50
 12 AC 96 27 B0 5A 06 9E 85 77 E9 C6 3F 01 9F 9D
 0F EB 04 C2 6D BD ED 5E 3B 3D 58 91 37 1A 8D 74
 50 8A 90 20 F6 61 93 0B 3B FC 42 DC 02 B9 BD D3
 0E 71 21 28 F3 EC 8A 80 58 74 65 9F 33 FE 5C 89
 C2 C3 6E D7 47 EC 19 56 43 4B F3 81 16 0D 8E FC
 70 AA 9D AD 3D 93 DB 0E 3C B5 A4 1D 2D BA 8E C3
 78 EE DD 76 EC 0A 55 51 0C A4 AB A1 5F 78 FF 2D
 62 21 65 D4 70 87 AC FA EC 0E 4D 06 AA 9C A0 CC
 9C A2 E5 4C 37 0D 1B 4C 34 46 6D 4A 81 D7 C2 F9
 06 DB 8E 69 0A B8 B5 CC 0A E2 9A 2F 72 8A 3F 27
 48 5A 65 E7 57 53 50 21 B7 67 41 00 7F EC 68 91
 D4 28 FC DE 8C 5C AF 41 38 3D A7 F0 73 25 BB 8D
 03 2B 4A 64 1A 0B 95 5C 68 22 44 05 8B 8F D7 30
 94 E4 15 FE 53 BD BD 9B 4E 9C C2 1C DC 26 10 93
 05 1F 19 60 97 06 E6 23 35 90 18 71 F0 81 55 DA
 A1 E0 F4 00 44 E0 2E D2 44 E4 1D 38 2F 1F 00 E1
 31 68 26 9F 63 82 38 DA 73 6C 15 DF 89 1B 81 35
 91 D6 C5 4C 91 8F 89 45 EC 54 A0 48 D7 D0 1A BF
 51 8C 53 9A 87 BA 7F 05 04 81 DE 9C BE 7A F4 34
 D1 0B 7C B4 58 91 12 D2 22 04 10 47 DD F8 D0 E8
 A1 28 67 0D E5 C3 A0 21 EE 22 6C B4 75 F0 13 87
 61 BA 73 09 58 2B 6A 27 35 2D 59 04 DF 1F 84 79
 41 86 59 20 31 3D 99 65 2A 86 A4 A0 CA 86 12 CE
 E7 DE F4 F4 F7 4A 5B 94 03 EC F0 95 48 83 03 C0
 67 FC 1E BA 6E 5C 04 B5 05 B0 23 CA 80 E7 6C A7
 F8 5E 73 29 E4 EC 4D 35 E5 65 BF 31 EC 45 E5 EF
 33 B3 F5 51 7D 06 B4 A7 B9 DB DA A2 35 83 A0 69
 E7 C8 96 F6 2E C2 FA 62 F7 06 D8 C6 0A 2C 36 AF
 0E 99 45 07 A7 11 D8 30 B8 1F 90 E1 6A 1D C4 A2
 57 C1 5A 57 1A 0A 0C D2 C0 40 63 AB F0 1E 67 CB
 73 94 12 05 D9 25 BA A6 2C D1 0B AE 12 61 0B 98
 0B 29 50 F2 D4 94 43 17 37 3B 4C AF 5B A7 22 A1
 7C 2B 21 E3 83 73 A6 A1 BE 9D 26 4D D3 26 F5 A7
 10 58 E5 6A 6E 10 1E A5 8D B5 92 99 E6 E1 94 07
 04 3A EE 4C E6 1E FD 97 AE 74 DB F2 93 BB B1 02
 7A 5A EA 39 BA 22 38 CF E9 99 E3 1E D4 EA 59 69
 A7 5F A5 04 35 7D 42 A2 F5 A5 6E C1 28 46 6F 83
 E9 D5 8E 81 68 6D 3B 2E E2 98 4C 4A C2 A3 A1 3C
 0C CA A8 96 40 51 B6 B2 B9 4B 5D 5C 01 A5 7C C2
 B8 39 0B D4 11 4D DF E5 89 21 FF E9 79 56 C4 58
 DB D9 3F 2C F1 83 90 14 CD 9D 2C D1 E4 AF D7 C0
 65 DC 5C A3 97 CB F6 E5 31 62 39 AD 86 F8 E4 67
 21 CB 46 6F 18 47 C9 AC 69 F7 27 7C D7 79 89 31
 FF EC 2E 0D E6 3B 05 D1 9C 8D C0 B5 D6 A2 EF 98
 3C BE 20 D7 B2 EE FA 73 41 DB 5D E9 87 53 20 71
 14 09 60 11 E5 4A F3 6B 2B 8F EA 7F 6D D1 14 D3
 16 CE C5 81 DA D6 28 F1 54 CE D9 18 F9 C7 23 2E
 44 13 F3 70 8B 80 D7 02 CF 51 78 20 BF FC 0C 3D
 80 B0 61 05 2C EC 61 14 63 84 A1 55 2F E6 1B EB
 E4 86 B7 B2 6A E9 DE CE 28 C2 6D 46 E3 13 56 AA
 4B C2 3E 1B 90 9D 5A 51 E8 E5 FA 5F F1 40 60 C4
 FF 10 95 6A 69 4B 98 CB C5 15 34 45 6D C0 33 D2
 49 1E 40 D1 A8 AA 57 23 D7 03 7A 33 41 F9 3A F1
 BE C6 BD 78 D0 87 51 68 E0 3F 49 02 C9 CE C1 9D
 21 63 77 BA DE 06 94 F5 FE 83 85 30 09 C2 E2 55
 AC 78 90 34 06 DA 3D AD DF 73 12 02 0B 77 9A CE
 B0 A0 FE 38 F4 08 ED 35 CC 27 9B 4C D0 2D 4A 1C
 3E A3 09 21 AC 36 70 E0 11 78 0E 6B 5D A8 50 47
 F1 E3 B8 FE 7F 08 72 05 96 87 0D ED 2A 74 48 89
 ED C4 8E E4 DC 29 99 18 3D E1 D5 85 E9 C0 5C 1A
 40 5F E7 38 7F E4 64 81 8E 91 3B 76 40 F7 D5 4B
 83 85 6E B1 BD 1E DD E3 5E 45 00 89 42 10 23 4E
 3B 99 C7 73 10 65 90 D3 3E 78 81 24 4D D1 2D 7A
 CE 4D C4 DA A1 74 B1 51 D0 32 D1 AA 42 3C E0 D8
 42 77 31 D8 4C 2A 2E 05 92 83 E6 51 49 5B 4B B7
 04 CD 98 E7 38 01 68 3D 10 27 A5 AF 02 73 58 70
 48 B8 DC 63 92 75 37 32 6F F3 E0 C0 49 62 C0 28
 B5 74 AC DE BB 2F 12 E1 4B 83 FE 36 3B 6F 40 3A
 3C 5B 6C 5E C6 81 EF A2 C8 6B 6B C9 10 86 57 1C
 1E C5 73 F1 D2 DB 43 F2 69 CA CD AE C5 87 03 7E
 F0 85 0B 91 09 70 AE 41 CD 91 A1 DD A4 D0 D7 92
 3B 83 4B CA 17 BE 9C 23 71 1A C4 6F 7F 73 DF BC
 17 C7 23 5A 93 35 49 D1 CC 74 FF 8A D1 1D 50 7E
 6D 5C 62 A3 4F 35 03 21 0E 9E F4 08 E5 75 ED 04
 DA 15 98 BA 3F 3F 2E 41 7B B3 32 25 57 96 44 53
 F2 2C 19 C1 AE AE BB A1 2D 2D 78 8D 08 20 FA E1
 3F 7A 3B 4E 14 04 3B 5E 85 2E DE 6E 95 27 6C 84
 A5 35 2A F4 E3 09 64 44 98 36 65 25 66 5A 1C D1
 8C C8 C2 35 6A EA 87 67 DB 8F 65 5E 12 12 23 E2
 45 57 FD 3B 10 FB 5E 1E 0E 42 B4 A5 06 9D C8 1F
 55 D5 8E A6 D8 1E F0 FD AA 38 67 4B 97 13 62 FB
 DB C6 A7 25 B4 9B 75 68 8F 47 1A 89 2C 1A D2 B9
 5B 33 DA A7 1C 86 2F 1D C5 5E 36 D1 D3 BD B6 9C
 4F 50 A7 7B 12 CD 67 C2 DE 4A E3 77 1B 34 FB 71
 D9 0F 9C 93 09 D9 83 D5 08 97 82 D6 20 D7 B0 96
 1D 55 D6 87 E5 A1 C8 3B E1 A1 3A 1C 7B CD 64 CC
 13 20 02 24 16 7A 73 E5 3F D4 09 BD 50 BC 8F 07
 8F 77 29 EC 66 A7 AF 29 30 4C A0 A5 61 84 89 7A
 D1 C1 63 E3 E2 97 24 E7 15 D2 E6 6A 41 DF 74 B6
 B3 8C 3F 28 1A 11 8C 84 9B E9 C8 BF 50 E1 FC A8
 49 B3 2F A9 DC E4 65 57 68 CF F7 26 72 2C 2F A7
 B7 01 C1 84 B4 D9 67 BF 65 67 2C B1 58 01 0D 7B
 90 6C 87 63 E3 46 BC AF 74 7A DD B0 10 76 C1 A7
 66 4A 32 81 82 B9 BC 24 20 71 9F FF 41 A5 AB F5
 F0 6D 0B 4B 07 13 77 38 4C 84 92 14 A1 61 B5 9B
 0B 8F 5B 3C AE D2 68 7A 9F 62 5B 59 17 6A D7 7C
 78 D7 24 34 A7 9F 96 87 33 B6 57 58 78 7A 74 76
 7C DA 3A 56 77 EB AD 66 6C CD 0A DB 85 F5 F1 EE
 91 97 BF 99 2F A4 F8 EA 87 A1 8D E8 22 84 01 E2
 C6 DB A2 02 49 3B A3 CE 6D DC A5 9E AD 38 13 35
 BF B6 83 4C 22 89 D0 F8 FC 6E 4A 54 47 9E C4 55
 C8 83 B7 75 A6 3F FE DF 7B F2 1F 80 47 B4 86 8F
 AE B7 16 B6 BC 68 01 92 94 5F E0 40 CF 7F 6C F1
 A7 89 B3 22 2B 1D F9 F9 B2 9C 9A 3E 1E 1A A9 A4
 6C 31 E3 FC 95 99 62 6E D9 C5 14 3F A4 9D 2E 85
 6F DA BF AD 69 56 CE 18 17 E3 E2 3E 7C 21 5A CF
 83 B2 13 BE 06 83 9B B0 46 E9 FE 30 C4 CA 72 46
 2E 5B 94 76 1C C4 4E 1E 9E 99 5B 01 AF D7 C2 6F
 FC 87 8C 76 44 AA 74 F9 1D 69 7B 69 19 1B 8D EA
 C4 3E 84 4A B5 39 49 5A 5A 95 4A 92 7E 06 84 FB
 13 E0 A2 8D 15 87 EC 4A F4 0C AB 0C 28 D7 9C 0C
 E3 FA B7 D5 5C 4D 60 69 57 FB 63 E2 EB 5D A0 03
 E6 F7 66 2A 20 91 3A 1E 3D 71 11 A9 BF 58 82 32
 AE BE AF D8 7A 69 2F 8C 2A 75 06 4D EE F6 12 2E
 1A 9F 7F F2 A7 A5 33 A5 6E 03 E7 28 C6 2E C6 19
 E4 32 6E 1D 90 86 91 A8 B6 4A 2C C8 6A 15 AF 56
 A0 30 0C 81 31 09 AC 64 EA 54 65 F6 D3 3C 56 81
 72 10 BA EA B8 AD C3 8C 89 B3 FD 24 78 C6 ED 5F
 2C 07 19 3C 1C BB 48 F8 1D 20 F3 B0 71 90 15 AC
 E7 62 66 8B 05 AF EA 22 86 E5 DB 6D AF 41 C7 5B
 1E 52 FA B0 DD 55 0B 21 E2 97 13 3F F0 D4 F4 8C
 C7 5A B8 E2 D6 EF 1E AB 11 AA E0 A8 59 D7 E4 84
 CB DB 6F D7 35 00 7D F0 B0 BB 32 51 55 9D D1 C1
 DF B2 A3 58 28 54 7D CC C1 73 35 72 62 6F 8D 8E
 94 8D 37 92 D1 3E D7 3E AB 98 0F 00 57 2B DF D4
 41 8A 6F FD AC 0F 92 23 83 E2 EC 50 A6 70 A1 58
 C9 59 C2 96 B8 67 F6 E9 01 E1 F4 79 B1 54 D2 C5
 BB D3 3E AF 09 6C 00 83 F0 F8 63 E8 5F 34 7A C7
 D1 FD AE 80 03 D3 50 76 D6 CB 28 96 2F F2 2F 8E
 4D 2A 4E 66 8B 60 8A 17 B0 3E D5 35 34 18 2D C5
 9D AB ED BA 27 77 F8 D0 C5 95 A6 A2 72 81 A0 81
 CC D3 72 77 48 4E 14 8D 1B 90 DF 01 4D 3A 43 D6
 20 08 B5 DB 91 9E 24 D5 CF 56 4B 1C 53 C1 2F B5
 0C 29 D9 99 94 E8 1D 14 78 35 94 3B FD 61 89 C5
 09 D2 D6 8E 41 D1 35 E1 E5 03 C5 E5 8C C7 43 42
 3A 1E 61 56 3E FB 71 02 65 01 63 4A 2B C9 D3 38
 5E E3 13 41 F2 79 6A 35 0D 06 76 33 67 4A 1A 03
 34 1E F7 AF D3 42 6B 0E 00 AA 56 FD 5B 05 25 13
 E3 F3 83 2D 1B 2D 9A 3C F9 77 59 E3 CC 4B BC EA
 AA E5 30 24 8D 51 C4 B1 7E 0A 8A 79 95 EF A7 4B
 7F 77 8F FB 14 BE E1 BE CC 83 4E 8F FB A4 3E 99
 4E 3B 9D C1 27 05 CA AC 9F CA D5 3B 6C 76 C9 24
 98 E4 3C 7D B2 CD FD 60 E3 60 2F 4E CE 3E D5 69
 03 7D 8F B7 5D E2 81 87 D1 17 1C D4 FD 71 C2 94
 BA 57 C5 09 20 45 97 3A 01 14 93 A8 7E D6 70 34
 14 F2 33 30 E9 E8 BE A9 23 F6 CE E4 AB 9E 68 62
 41 71 95 D7 F9 6E 94 90 6D 7F 74 07 26 37 DE 15
 CC E9 34 8C 48 74 FB 3E 0D 9F 1A 0E 31 72 5E 91
 01 FF 6C 2A C7 53 D6 D7 3D 46 E0 16 9B 3F 20 B9
 7E 19 E8 DE 93 22 6F AC D0 B3 C1 1A 1F CC F3 49
 E4 E0 44 BD EF 9E 54 D9 6B BA EE 91 2A 24 4A 3E
 2B C9 AB 8E 37 FB DA 94 A7 1F 7A EF 67 AF B6 77
 EB CB A3 05 CA 46 83 C8 33 76 9A D1 B1 AD 39 41
 C5 A1 21 4C BA 8A EA B7 F4 E3 7F 25 DA 72 5C D7
 76 F1 5B 8A 78 42 B3 AB 73 EE C7 38 EC DB 2C 21
 6C 7B 0B 46 F2 94 EC F2 29 CE A3 EF 4B D9 3B CD
 1E 5E 00 A9 A1 4C 76 21 59 5B 0C 27 4F E4 20 D2
 39 0D F1 F1 6A B5 A9 C8 2D B8 EF A1 A9 B8 54 B0
 C4 DE 7B 3E 0D 51 0B 98 4E 35 02 48 04 C2 F9 91
 1A 80 2F 73 EC C0 40 3E 89 B7 94 24 D4 10 81 EB
 CA 0A 66 36 03 FA CE 90 21 38 09 08 C5 97 BE F1
 25 25 AF 96 0D 62 C8 EA C2 33 89 46 AC 3F 4A 33
 98 D7 91 B8 B4 38 DD 48 FE BF 2E E4 F9 A5 9A BE
 51 EA 9A A3 D3 67 00 43 A6 6C BE EE 12 E1 C6 53
 40 90 14 0B AA F5 B5 4D D5 9C B0 71 3B A6 D5 96
 B4 68 DB DF 2A 4B 13 D8 B5 33 CF 91 C8 3D FD A0
 9C 6C 14 C2 7A 06 86 E9 FF 66 51 59 B3 7E 2A 1B
 46 94 79 C7 47 67 F1 67 08 9F D0 C9 BB 0E EF 58
 88 EC 7D 8B 21 13 DB CA 71 15 82 84 91 7D A6 D9
 14 83 E1 BA F0 CA B6 FF CF 21 7B C0 60 C0 30 52
 37 B0 7F C8 FF E2 70 5A 06 57 75 01 D9 D7 1C 0D
 40 B4 41 C0 65 EA 3B BE 02 73 6E BF 1B EA DE EE
 95 DE 2A 58 13 19 8C E8 2D 47 9F 0A 75 02 41 5A
 8B 71 0C B0 DC 19 91 EC 7A 88 65 29 2A 87 76 BE
 AA 9A DD EB 63 EC 8C C4 39 BB 20 CA DC 32 80 2D
 3D 40 C6 D2 2A 98 8B BE A4 8F 75 9B 31 9D 35 FF
 DD 96 E1 9E 82 84 73 3B 5E 9A FA 3E 7B 25 F2 0E
 A4 4F A8 80 3C B1 1E 7D 34 75 C7 7D D0 5A 3E 86
 72 DD 1B 05 9C 18 F2 0B CC F2 87 D7 D2 8C F3 99
 51 81 C5 E9 55 2D 1C D7 32 8B D2 78 44 5D D3 72
 7B 6F AE 34 DE E7 E3 F1 0E CA 24 55 A9 38 37 B2
 04 F2 C4 D0 27 AB 14 EB 97 62 CC 52 06 C6 AE F8
 92 EB 4D D2 AB 51 D1 89 37 C7 9A C5 BE 3C 53 71
 7F E5 E5 A2 44 6B 02 E1 69 D2 29 97 DF 09 7A 9A
 CE 3F E2 42 D7 BE B3 FC EC 0F B7 C8 EC B3 73 18
 F7 CD 81 0A FF 56 D6 D8 16 8D D5 09 8A 1A DC AC
 7B AA 71 60 95 20 06 B0 ED 7A E4 17 3B EB F4 79
 29 6D 7C 9E 25 16 CB 5F 90 CE 55 DA A0 4A 30 18
 BB 6F 3C EF 4B B4 EA 3F 4A 0F 49 97 7C C1 7E 1D
 6A 77 97 EC E1 7F 34 7F 33 36 5F A7 2B CB 81 11
 05 53 69 F5 E6 23 DA 67 37 B0 EE 53 72 13 18 20
 75 15 0E 40 5B F1 D0 3D DB 73 95 A9 D6 8E 49 11
 D3 09 5A 83 12 7F C4 34 FD 89 6D CA FF 5B CA C3
 FF 98 A0 22 FD E5 13 BF 73 FD 86 C6 44 83 E1 0E
 A0 0A 4E CD 5C 50 E6 49 2B E9 07 66 54 A6 E0 A6
 21 2A 42 A5 7F AB E0 DA 36 7B 45 94 57 90 62 29
 53 15 1D D3 AD D4 86 0B A5 11 96 63 8C ED DC B4
 E2 41 60 6B E3 7B 71 4E 69 28 1A 52 AE 11 98 D5
 D5 90 D2 DF 54 63 E4 E1 43 67 4B 27 8F 78 CC 65
 46 77 C4 A6 65 01 5D 7C 48 24 9D CD 7C 9C 2E D0
 72 0B 8B 7D C2 BD B1 29 CD 7F 90 3F 12 70 FF 07
 B5 1C 9E D8 77 BF 31 9F 0F 33 C6 74 26 1A 88 1E
 20 73 0D 1E AD 48 95 52 51 29 DD EA BA EF BC 90
 4A AE F1 9A 85 73 6F 7B C8 33 34 DF BB B0 21 64
 7E 83 13 87 EB 37 E2 5B A2 52 98 0A 6C 90 4D 8A
 B4 5E FF DA 34 B8 9D C3 55 F9 20 43 1B F8 E9 3D
 2C 89 8C 07 3B 31 B5 0C 9A 29 F0 CC E0 AC 57 33
 71 4C E9 80 23 EE 28 E1 64 FB 3D F1 C6 8C 29 FA
 BC 51 7B AA 0B 31 F9 0A DC 69 5E 1D FE 9C 8C F4
 23 5F BD 12 FC F8 9D CF 4E 85 6F BD FA D0 48 EA
 69 FD C9 73 6E 5E 11 4F 1A 66 04 5A 14 88 D1 76
 68 9A A5 75 E0 DF 99 29 62 CA C9 7F AF 34 A6 E7
 80 FE 8C 01 A6 2F 55 8D A3 69 DD BF FB 83 AB 7A
 28 82 84 0F 1D 5C 74 77 68 77 9B E2 1B 0E 6F 86
 9F 31 35 64 3B 55 1B 59 F4 D1 23 59 47 E7 ED 97
 D6 E7 1A 40 95 87 2D ED 2C ED 56 41 A1 FA C5 2E
 20 92 D8 AA B9 3C 7A 12 6D 73 4C 3C CE 94 AB 30
 60 5D 32 07 A6 0B 2A 17 39 9B 13 CE A2 C5 D3 59
 8C 83 8A 10 C6 C8 DD 4F 6F D6 6C 8B 0F 50 41 A3
 27 6C A8 5B 1B A7 67 D6 31 34 F2 2F 50 D7 9A 3D
 E5 6B 29 D3 55 F6 08 C2 F3 A7 F6 45 CA B0 FF 53
 42 02 A3 58 F5 DA 27 DB 33 69 5D 9E BB DB F0 84
 B7 EA 27 47 F8 DC 94 49 3A E4 31 5A 69 42 30 7D
 9B C4 46 46 8C A5 C9 88 80 CF 9F 70 ED FA 6A 13
 CC 39 69 08 48 E2 D4 84 C6 C5 5A 64 7A E2 09 D5
 D5 39 D2 AC 81 6D 33 F2 FB AA AF DD 7A E2 B0 DA
 1E 95 3D 0C 0C CD 22 E5 26 A9 51 AE 02 CF 95 EF
 6E 16 BB B5 1E 1D 76 F8 00 3E 19 9B C7 10 44 CD
 0C 48 EF 92 D7 12 5C 23 CD 57 15 E1 50 F2 CD 63
 FE 3F AE F6 C3 59 D2 16 D4 EA 71 7D E9 41 40 F7
 FD C6 B8 C6 F8 11 5F CB 31 28 4A B0 4E 13 79 51
 39 AE 19 8D A5 C6 8B 52 AB 8F F2 F3 AE 39 D9 46
 AC E0 25 26 8E E5 94 97 6A D6 60 C0 E7 7D 12 D2
 57 0A FA FB 84 60 DB 5F FB 7B 6D F1 EB A7 D7 41
 13 14 3B 30 DF C5 27 D7 3D B0 29 23 6D F4 AA 2C
 93 5F AB 2A B3 B8 4F 1E 34 2C CF 6C 9B DA CB AD
 84 DE 1B E1 CB 2A 94 14 88 5C CD 75 C7 6A 2F 8C
 24 6B 4F BA C8 BB 99 C8 31 E5 ED 19 5F D6 34 FD
 22 54 1C F8 31 63 49 18 AA 93 F7 98 45 D7 09 33
 EC 6D 2D D5 D3 41 99 BE E4 89 BC 86 DB 32 E9 9B
 FD DF 33 9A CD 9D 42 0C 68 BD 85 84 25 F9 D5 59
 8B 7A 8E EE 64 18 F3 26 C0 D9 C3 73 F7 CD 83 29
 1D DE B8 2C DD E5 95 65 9A E9 F5 63 D2 56 CF 9B
 65 32 0E D6 4E 07 70 E2 4A EA 07 18 BB C0 AB 9F
 05 EE 88 7D A4 DB 76 80 A0 AB E2 D6 25 0A 09 E3
 83 16 EA A7 9A 82 49 7A 7F 72 C3 15 D8 0C 57 C7
 D3 E5 09 B3 FC FB 7C 6B 19 EE 56 4B C6 3F 46 77
 32 E7 7B 4F 23 DF 73 F3 BB 76 57 08 C4 6D 27 B7
 ED 3B 8E 06 2B 31 22 B6 64 55 0F 6F 31 8F 3D C8
 59 83 A0 B2 99 8C F0 3D 33 39 38 1B 79 2B 89 41
 78 24 8C 25 10 1F 97 CF 4D 8C 98 44 1B FC C6 F9
 59 D3 20 F4 FE CB 55 ED 16 30 C7 11 26 C4 C0 EC
 B4 0F E6 39 A6 96 00 12 7E 45 DC C0 1E 55 77 E4
 94 1A FF 66 07 CA F3 1F 42 7B 61 28 2F C5 78 60
 3F 4C 7F AE 6F AD C5 E6 A1 8C 14 03 21 4E E7 42
 3D A8 BF DE 7A 21 C2 9C 01 44 98 36 27 8C 8E 38
 45 6C 3B E1 3F 5C 9D 18 16 1B F5 58 37 69 22 81
 51 50 09 5C CA C3 93 3B 56 65 3A 2C 2F 5D 26 21
 94 37 63 90 99 45 DF 91 EB 70 78 B7 B9 97 73 DD
 6F 44 38 7A BA FE 66 D5 AE 8A 35 9F A6 52 F2 0F
 39 04 ED 23 17 3C 21 7D D5 DB 7E 8E 36 06 4C FC
 C7 BE 39 8C C0 E1 4D 52 CE 31 C7 03 C2 33 30 43
 5E 52 C0 B8 9A CC 9A BC 3E 46 47 8D 3A 81 16 34
 34 E6 F2 74 B7 0C 25 E1 90 30 8C C2 7F 63 0C D7
 1E 95 D4 50 00 FE 57 4B 2B C0 1E 90 67 B8 19 A9
 6F E1 68 41 BC 46 7C A6 5F BB AD 01 86 71 15 E1
 2F 31 21 1B 81 3C EC C5 87 E4 BC 5F 2D 93 31 DC
 1C 17 54 74 54 55 96 D6 4E 58 77 E5 3E 6C 4D CE
 29 6F A7 86 21 59 41 BE 36 0C BE BD 96 EA C6 2F
 CA 26 2E F3 4D A3 0A 54 26 63 A5 47 CA 73 ED A6
 8E 49 CA 26 69 30 41 83 B2 89 56 41 E4 FA 1C A4
 63 5E 3E E7 7A 24 1A EB 70 14 F1 22 C2 9C 54 74
 FB 89 A5 BE E6 A9 CC 2B BE 00 0A 89 FB 62 BE 9F
 F4 B0 BF 06 79 5A 06 45 6B 33 8E EA D8 50 FA E5
 30 83 DF B5 33 66 BD 1E 00 E1 06 EA BB 1B 32 21
 A7 B1 8F 02 8B 8C A6 E5 B1 95 5B 2E B6 C8 85 53
 80 C6 28 A9 1E B3 D8 59 E5 F7 30 C9 24 DF 98 96
 2D 6F 40 32 2D 4F 74 5E A5 A8 02 4C D5 87 7B 70
 B5 D3 D8 A2 CD 2E C1 AF E8 19 DF 5C 7E 7B 8D 5A
 01 83 08 2F 85 CE 87 4A EA DC BE A4 C2 FC E7 FC
 CA 3F 58 C1 FA 72 EC 1A 62 98 45 DA D0 40 93 38
 A5 34 BA 55 C5 98 45 7B 3B BF C6 33 4B 88 BA F3
 0D 31 AF 78 31 7E F1 4E 0E 29 3C 49 E8 94 88 D5
 14 72 A0 2F 10 17 7A 66 1D FE 59 B5 31 31 41 39
 1F 3D 28 07 91 74 04 5C 1D 97 B9 50 8C 96 C1 F0
 0A 68 EF C8 C4 80 7C FA 01 B1 16 B0 05 9B EB 58
 BF C1 14 12 07 30 4C F6 D8 2A 0B A1 71 07 9A 43
 39 D8 32 FB 61 83 25 34 68 F4 39 48 20 DF 58 A3
 03 05 28 FB A2 DE 13 DC CB AA 60 36 57 56 A1 28
 AE 36 59 0C 29 88 3B FA 5C 39 8F 16 48 35 86 CE
 BD 21 15 EB B8 86 D5 5F 56 DC B0 0A E7 B6 91 1A
 9C C6 CE 45 61 44 99 61 C5 77 30 E0 38 C7 06 6E
 62 04 92 88 42 8D 3B 49 12 0B E7 98 11 E7 C1 C2
 65 0E 03 6F F2 07 5E F7 39 F6 1F C0 06 E1 1A 61
 CD 9D FA 22 A2 E3 8B BE A5 6B E2 DF 4B D7 E5 86
 0C 40 F3 A6 17 CE F6 BD 73 74 82 82 28 1A F1 33
 9A 4E CB 0E 2A A0 BF B0 5D D4 9B 42 48 5B 05 7A
 DF 74 F6 A4 75 73 36 76 BB 47 75 E5 22 FF E5 58
 1A BE 2D F1 3D C8 28 56 97 6B 26 47 FB F9 DE 83
 12 EE 44 15 07 8A 15 4E A6 D2 FA 25 C5 41 DF 25
 5F 20 27 F3 62 F5 5C 09 C2 76 1E DD DE 7B A4 05
 33 67 B5 6C 01 26 1C 98 D1 4F 2E C9 22 CA CF 0E
 68 D8 38 83 C9 FE B5 13 4B DA 42 89 BB 7C 87 83
 93 82 C0 F0 F5 C3 A2 38 27 02 28 03 2F 20 AB 5F
 F2 4B 1B 59 9E D2 91 FE AB F6 F7 43 36 0F 92 5D
 58 CC D5 16 42 E5 D9 F1 74 5C F9 22 D6 A1 35 13
 8B CD 21 5C 0C 22 B9 4D A9 09 4B 6D 12 E1 09 55
 CC 1C 33 47 9C 3C B9 C6 4B 51 E8 2F 76 28 2B 99
 C6 0C D1 81 4C 9B 1F C6 CC 13 1C 38 DF B7 48 05
 7A B6 4A 7C 4D A1 1C 2C 61 D8 84 F3 7C 01 4B 6B
 AA 67 65 81 A8 F5 63 AC C0 44 A1 62 15 D9 3F 3D
 D2 80 7B 52 B2 6E D9 59 C5 42 11 B4 FD 6B E4 71
 EC F1 F5 45 A8 E5 FE 71 4E 18 9A 42 15 1A 19 3F
 29 43 93 AC 8C 6D FB 95 B2 E2 8A 69 AC 1B 1A 88
 4D 5D 0D 14 46 9C 65 4A 8E 83 EC 90 04 5E 96 9A
 E6 9D CF 5C 58 63 DF B9 84 3A 99 56 46 28 35 89
 7C B3 22 C6 DE 8B E3 BF 03 5F 05 34 43 AF A6 32
 31 A5 9E 25 8D A5 99 D9 C1 95 05 65 3A AE 88 C6
 77 44 58 38 4E C3 00 10 8B 2C AD 7D A1 0C 2A A6
 1B D3 76 BD 22 FC AA 77 EC EC B2 A7 22 3D 37 27
 2F 2E A2 47 92 7C A7 2F F5 A8 DA 50 86 5C F2 B0
 65 C0 79 14 EB 6C 29 3B 0E E3 1A 2F 0F 78 D9 C6
 C3 13 AD 2C 9D F3 23 9B B6 E7 EA F4 F6 26 2F D9
 95 E3 29 EA 5D 91 2A AE C0 25 11 13 1C E4 A0 DD
 B3 D7 88 43 5E 64 E8 9D D6 3A 2F 45 82 F2 74 7C
 80 42 75 F9 3E 59 D4 E2 31 E3 96 DF 66 24 19 E5
 1A D2 70 31 DA F2 B8 3A 66 F4 AA F0 79 61 BE 03
 F0 EF AE 65 25 EB DA 3F E9 43 CF AE 3C 56 3D 90
 7B 9D 9F 28 3E 2C AD B7 F6 0F D2 3F 25 D3 ED 09
 96 D1 53 8F 7D 66 B1 16 33 92 09 0C 02 54 86 AB
 39 5B 22 CB EE 68 AF FE 38 50 4E 12 E6 AA 85 C7
 56 BE DA BC C5 1A 31 66 BB EB 60 BF 64 3A 6D BA
 27 8D 9B 3E C1 4C 97 AC F9 7B 16 73 96 57 BB BE
 5F 9E 2A FC F7 25 64 3E 9D 20 84 B7 FE 61 87 A6
 99 E2 4F 91 97 3D 35 B6 46 7D 54 EF 2E 0D 4B D0
 24 A9 40 F7 A2 C9 ED 7D 4E CD 0A 18 58 78 A4 AB
 E9 11 B6 38 D9 97 32 C3 A3 A7 E5 67 50 F6 EB FB
 6A DE 63 F3 CD EA DC 42 68 D9 B1 02 0B C8 31 18
 D7 CA CF 6E 86 69 C3 F3 0B 37 04 6F 97 83 21 40
 2D 1E 15 06 37 F1 7C C9 F9 94 ED BE 28 87 59 EA
 A9 23 96 96 DB 0E 60 FB 5E D0 14 CF A9 96 D6 B9
 61 3D 0A 2B 97 FF 63 BD 56 7F CB 96 67 12 9A 38
 D8 04 40 B5 87 19 B5 AC D4 7D 8A DC 4F 65 8D 53
 D1 A2 95 B1 20 F6 91 F2 22 32 B7 90 4E 2B A8 28
 B0 5C 0A B9 7C 10 72 75 18 8E 7F A0 AD 3B 81 46
 41 94 CA 38 7E EA F6 D6 83 8C 98 AA 11 9A 93 2C
 A3 59 5F E7 CB DF 29 30 27 58 61 7F A9 D4 27 3C
 13 CE 29 B6 A7 19 8F 6E 2A F2 BC C6 AB CA C1 FD
 DA BD AC 55 53 02 EE 38 9C 91 F1 BE D5 D6 24 2F
 A3 CF 14 00 D5 CF F7 DC 98 4C 96 5E 25 60 01 76
 BC D2 14 2A C1 AB 19 A3 28 42 07 90 02 48 99 2F
 6B 82 29 CE C9 D5 D1 B0 F0 ED D9 E1 2C 1D 7F 20
 52 AA 6B 4B A1 95 F7 96 A6 41 47 8D F4 1C BD 3F
 D6 64 D4 C9 E5 06 98 91 29 65 79 C4 7D 49 1D 78
 A5 5C AA 0A C6 4F 0A A5 9D 8D 6E EC 22 47 07 57
 F4 BF 2D C5 C3 E0 CA 83 17 02 99 DB 6F 43 01 4A
 A5 94 A9 39 DC 47 D4 53 7C A8 98 D3 DA F8 F4 93
 AE D7 28 11 24 91 17 A7 A8 1B 03 44 0C 01 C4 3F
 64 56 CC 7B CB 34 96 FA CB 08 0F A8 61 0E 35 FE
 BF 00 97 54 41 20 7D FB 00 04 CE 61 E6 74 A0 FD
 7A 9F FC D9 CB 11 03 7E F2 F8 FA E3 5C 5F 9B 98
 98 48 EB C3 96 31 80 DB 75 4C EC 5E C5 50 6A FD
 B4 A6 55 BE ED 22 6E D0 72 42 E8 8D CB 90 7F 83
 F8 22 B3 98 89 40 23 2E 1F 17 03 F1 C5 DC 87 6B
 6F D2 CC AE 3F 0F 71 8D EC 4B 1A 29 11 92 83 CE
 02 76 5A 47 E3 D0 EA 0D 83 F3 CE 57 4B 6A 43 4E
 B0 A1 CF 87 8C 16 F4 AB 18 F6 CD A4 91 11 6B 86
 B4 D9 44 5C 97 ED 22 25 A4 33 8A CE 19 CA D6 D2
 B9 CE A7 A1 7D 96 B3 D3 D6 B6 1D 6D 08 84 04 D2
 67 79 B5 02 81 E3 56 1B 16 D5 35 98 B7 DA 7F F0
 33 18 9E 6B 15 BC 0F 70 2F 71 27 7D F7 39 14 33
 D2 2F D7 D6 81 06 C8 41 2D 71 EB 3E F5 EB 28 13
 1D 44 A6 25 39 E5 BF 7D B1 D7 6B D4 37 CD 02 78
 67 8F 0A 3F CC 7C F6 87 9A 0F 49 D6 07 A1 5F 52
 DB 4D E5 A4 56 7D FE EB 62 41 B1 F5 F5 4E 9C 42
 34 B3 96 C2 05 E7 10 4B 5C EE 82 FC 36 4E 6E 10
 F9 1A ED BB 3C DC 6B B2 31 F1 14 F8 3F 84 33 22
 A3 41 01 25 2B D9 7D 2F BE 4A 39 0D FE 5C 8F 27
 02 07 B6 24 5B 33 B0 51 D7 F5 03 BA F6 34 B0 C3
 C7 8D 96 A9 04 02 D9 F9 30 40 EA 70 20 F1 2C CF
 03 2B 5F 9F FA 78 91 2B CA 73 B3 0D CC 46 5A A8
 15 AA 70 5A 82 5F 01 9D A7 C7 D6 AB 09 87 9C 43
 9D 96 A0 54 39 50 3C 2C BB 6A C2 47 19 66 C5 79
 7A 92 47 4F DE BC 3B EF 1C 6E DB 92 5B 4A FC DF
 F9 82 FA AF F7 B8 DF FD 1D C2 D1 AD B7 5E D6 66
 FE 63 2A D5 0B 1C 53 B7 EF DA AC 22 53 C0 FF F4
 61 7A FF 16 BA EE 3A BD C5 62 2B F8 DA 4D A9 26
 6E FC 9C 8B E5 F2 21 35 9F FA 77 6D 91 F7 72 AB
 CD D2 37 41 CD D4 59 EC 48 CF 22 2F 60 63 A3 57
 4A 1A EF 97 76 C4 7E 2E 1C CE AA 31 0B F6 C6 64
 A5 9E 5B 1C 05 4A B7 33 34 F4 BC 15 69 7B A1 96
 15 68 29 C7 50 40 5B E4 D3 38 B9 BD 7C E4 D2 D7
 A1 8D 4B 92 D3 B8 B6 AD 22 3C 11 48 93 84 7C 36
 4C 1C D0 F3 10 AE 5B F3 DD D6 CC 91 30 70 37 B0
 54 91 3F B0 88 4E 80 9C 81 AB 69 79 A4 5C 2B BD
 94 73 FA B4 6F 47 4C CF 38 49 E5 08 E4 A0 1A D4
 28 63 E8 24 76 E7 D1 49 D1 80 21 00 F4 62 20 EC
 03 9C 41 4C 3D 95 FC AF DF 00 27 23 BA 68 29 CB
 41 08 3D 96 18 D6 CD 1F A2 53 4F B7 10 6F 03 12
 8F B8 3E 59 30 86 58 63 FE 39 10 AE 72 8A 65 C0
 6E 70 0F 3F 4C EB 05 DD F8 4E B8 AE 64 28 BE E0
 3F 6B F4 E1 84 6D FF 5A CF 4E C9 6D D2 07 9A B1
 2F 6B 5A 12 A2 D6 9E 54 4A AF 3E 27 45 C1 BB D8
 9B 17 0B E2 3C AB FD 55 1F 6A C4 AD A1 A9 7E 8C
 CE 83 92 4B 2B DD D5 5D AF 8A 33 84 25 C9 5A 1E
 E7 DD EA F1 0B 31 8C 2E 25 04 15 6F BF 95 07 40
 13 57 42 B1 F2 27 D6 52 96 C0 37 EA 97 B5 E2 85
 0B 0A 65 70 3B 8D F6 55 45 CE 17 9A 34 76 4E 5F
 55 03 B4 FC EB 1C F6 BA 0A C9 6C E0 15 D2 19 23
 32 09 9E 9C 99 B8 05 71 6C E5 AD 4F 4A CF 5A 6B
 EA 9F 2A 21 35 6A 3B 2A 5D 7F 50 6C C2 06 3C 34
 7C FC 9F 23 BB BF E4 64 04 51 8D 0B CA 47 65 84
 3D 62 D7 A6 F1 EB 31 40 7E 87 94 3C E5 D2 70 EF
 6E C0 52 94 C6 C5 A5 21 41 8D 2D C8 4E FE 8B E0
 5B DC 62 B0 67 37 DA DE 2A 9E 94 C8 2C 01 47 65
 1C E5 7F EA 57 03 C5 33 5C CC C8 ED 61 22 5F 49
 7C 1B D2 2B 19 34 DF 81 87 1D 87 4B E7 0A 66 E5
 4B 78 C7 CE 1B 82 42 D5 01 41 8A E0 8B FC B6 E9
 0E E6 0C AE 1A B3 B7 28 20 48 D1 29 99 0B 69 4E
 91 AF 64 F5 EA 01 33 C5 04 F6 58 52 A0 39 4B D8
 B1 EF E7 CD 01 A2 79 2B C0 7E 5D 94 CA 7C 6D 8D
 13 4F DF E6 F7 BE D4 AE 8B 8F 4E 27 81 A0 A6 59
 75 D4 AA CB 72 2E F8 2C 64 79 43 30 CC 2A 46 F9
 08 F2 C9 C2 15 E6 1C 3F 57 BF 46 C8 F2 5D F2 59
 6C 91 A5 8D 34 7B EA 9B F6 4E 79 63 47 74 E2 85
 D6 27 6F 1F 23 C2 8C A9 66 A3 D0 65 77 61 86 6A
 70 0D 1B F5 94 05 55 4A 4D 37 86 70 53 1D CE 0F
 B7 EE 6A 1B 17 CB 31 F4 22 8E 55 73 BB CA D4 69
 15 9F 43 D8 8A 23 3D A3 1D AC 3B DE 96 C7 16 01
 EA 23 17 F1 3C F4 8D 60 74 5F 77 EF 62 97 52 8A
 6A A0 CC 6B 95 A4 F6 DE CE 92 6C 0E 4A 9D F1 1F
 BB 95 27 09 E4 0E A0 EC 30 E4 92 A2 46 74 93 9B
 B5 F1 F4 79 DE 05 0C A8 7F 3F 51 DE 3E EF 87 76
 98 A8 E4 2E 41 1B E8 21 25 DA AE B9 8C 3E AB 5A
 AC 4F 8C FE 27 78 FE 3D E9 DD 53 E1 FD 77 75 B0
 79 51 6D D8 09 DE DF 31 48 50 54 03 6E 6F 2E 73
 43 31 4A 84 31 3A DC 89 07 F9 E2 E3 8F 26 FA A6
 38 77 B4 76 C3 1A 51 AA EF 4F 8E 69 F1 03 1D B1
 0B 74 5C 5A DE 52 DC 62 86 0A EB 10 AF F5 1A 7A
 0C 23 7E EB 79 52 3E E2 34 C1 92 78 91 7B ED 8F
 A4 E2 F0 36 D1 5F 15 84 B6 F1 11 63 3A 07 DF E3
 27 2A 88 73 59 D4 5C E9 47 47 47 75 E1 A9 48 0C
 B0 AB BE BE FF B0 A6 C0 D6 8E 97 E8 A8 11 3E 1B
 F8 27 AA 73 3C 62 73 24 7E F2 AC E8 38 B8 B1 BF
 40 BD AB 52 0B 17 BE AD 8B CB 72 0E F9 4F 29 D6
 A7 1E 0D 73 FA 62 53 3B 24 A5 8C 30 48 BB 32 3D
 DA 20 50 98 71 21 25 39 6C AB 45 7B 8A 6D 16 24
 87 1A B5 11 AF AE 32 89 DF D5 AF 33 D2 91 CD 4F
 7D E6 2D A5 2F DC C4 1A F1 DA D3 87 F1 CB 42 89
 A1 BD 41 E4 32 8F 8A E7 55 FD 86 79 DE 8D 4C DB
 B7 03 4A A5 DD 59 61 34 F4 30 04 37 BB 70 D7 4F
 8C 99 67 1A 30 47 E3 E6 14 73 4C 4B 5D FC 5E 79
 69 05 8D 5B 10 3F 0B 5F 20 2D BC DE D0 3C 31 27
 C0 CE DB 8D 68 AE BF DB 11 69 FF 2A C7 43 32 CD
 3B AF D6 FF 0F 30 97 4C 37 99 70 B3 70 DA 75 FD
 52 19 11 F4 E7 12 BF 2B F7 EF F3 B5 77 51 A3 F7
 3B 9C 99 64 E5 25 47 5E 8D 2C C8 7E FC 91 84 7B
 09 6A 5E 12 FE F9 89 40 13 D5 0F B0 44 F1 82 30
 68 46 75 02 56 B6 4A 78 E4 CA A9 1B 3C CC 78 A2
 50 DB 15 01 DA 6C 4F 78 96 62 B3 B6 C5 B0 DB D6
 C4 1F 4A A5 0E 4C 76 FD D2 24 10 FB 2D B1 2F 3F
 A0 FC 07 EB D2 30 68 C5 85 FB CC 9B 91 F3 8D A2
 96 91 DE 2B D1 D8 D5 40 4C FC 47 F8 B9 31 A2 9D
 62 29 58 83 EA 61 8B 49 49 63 BF F3 FE 34 EE 96
 DB 6E 3A 33 2D 7A 95 29 9E 7A 3F 5D 14 9B 51 32
 5B 8F FE FD D7 48 FF 42 F1 D3 39 E7 14 B4 6C AF
 85 B2 2B 33 4A 2C CD 33 28 4A 2A D3 16 C0 BA B4
 2E 1B 55 5F D8 A8 95 09 64 EE 00 27 5D E0 7A 8D
 09 98 EF 39 8D 13 CE 71 B0 83 AD 0E E2 05 66 1F
 81 5B FE DE 70 47 40 FD 83 64 E6 FE 6F 3E 97 2A
 A7 83 B3 9B 47 1A FF 79 21 1B 2A AD 68 79 A4 E3
 F1 43 FC 65 EC 2B 35 14 01 12 A3 74 9C 4F 36 31
 F0 81 73 C3 C0 1F 2A 4F 11 16 43 A9 43 E0 43 BA
 79 EA 86 15 BD 90 4E 54 88 68 8F 0B 7C EA 2A 56
 EA A3 4A 57 BC DE C3 3A 86 79 FC 01 E8 65 37 31
 14 2E 0C 96 51 15 01 70 34 F4 B7 9B 3A BD 58 F5
 2B E4 FD 36 A7 E7 28 9B EB EE A4 A1 51 70 A0 C4
 1D B5 59 CF CB D4 9F 76 A9 0D 48 BF 9B 0A B5 EE
 79 55 8D FB 30 B1 A4 15 D0 62 44 59 D0 8E A8 8C
 67 2E 0D 0A D4 D0 D9 C7 1A 98 51 1E 4A CA 76 8D
 34 3D 6C 10 BD 03 FE 04 A3 55 B6 67 EE 55 77 70
 F3 55 FD 6A 5F 03 BE 50 D0 3C 71 F3 D2 EF DD 58
 CA 53 FA 7C 90 FA 88 B4 82 AB C2 22 25 F4 82 39
 2F 57 F8 3A CE 28 93 F6 D9 58 7A FD 60 E5 40 16
 B8 5F D6 89 F4 30 DA F2 A2 06 E9 B4 29 B5 99 7A
 C7 B3 97 A7 EE 5F 68 D4 0A 5F 3D 99 B7 0D 23 51
 6D BF 97 FE CD 32 DA 31 AD 69 25 8D 64 F7 7F 7E
 C2 F2 D1 3A AD 95 99 77 17 23 5B 0E 7D AE 2C 72
 43 F3 4D 6B 1D 8B 85 06 CC 38 A1 10 9A D9 08 DE
 69 93 B4 B7 1E 86 BB A5 DB 6A FC EE E5 31 66 3B
 AC AE 19 78 F6 32 51 AF BD 8E D0 4C A1 E9 46 40
 55 11 69 53 2C 2A 38 F0 4F B4 56 2B 46 15 98 EA
 0E 60 46 8A 9C 13 9C 35 A3 C6 48 26 77 B5 D0 EE
 5B 84 22 BB A3 0F 02 91 8E 61 49 1A F5 C3 BD A6
 18 6E FB 0B 7D 7E 68 83 29 61 39 62 7D F5 BB A9
 64 85 A6 92 A9 E0 E7 3B 20 DD F0 0A 14 E7 8D 7E
 56 04 4D 71 22 57 8E 5D 3B D1 FF 25 A4 63 C0 35
 C4 12 8B 5E 10 2F B8 FA 5E B8 17 89 9C 24 C4 01
 3F 7F 12 82 D5 1B 40 05 54 AA 5E 80 C1 4A 4E D5
 DD 48 02 86 8B 24 D3 49 8F 3A 36 7E D1 84 CD 04
 88 77 9A 31 5F 33 82 47 FA FF 58 9B BF DD 32 5C
 9E 7F CE 2D 40 2F FB 1B B2 5B 3E F7 31 7B 40 FE
 64 2C 42 DB 8C 01 3C 60 51 04 E3 2D BD 21 BC 31
 88 91 74 69 4E EF 43 BF 98 42 64 12 4C 4F 84 35
 10 84 77 20 B4 F1 CE DA E3 A2 81 E2 59 E2 8E 25
 0E D3 4F 3E BE A3 8A 1B 26 55 77 40 AF 73 34 C5
 56 C5 F5 E2 C0 BC 5E 28 53 FE 16 78 91 19 5D DC
 B0 08 99 3D 48 13 51 41 C2 D0 90 20 76 20 DE 26
 59 9B 49 66 CD 14 52 73 41 7A 9A 78 CE 5F F2 BD
 FF 05 30 5C FD DE 0A EA 72 92 DC 7A DC 32 AE EE
 06 5A 3F EB A5 C9 7B F9 60 06 4D 0B 28 9D D5 D7
 52 7E B9 4F 69 85 9E 60 B8 F6 17 A5 DD A9 41 4E
 69 F0 B8 66 FE 29 E7 71 53 63 C1 29 1F B7 1F CC
 D7 E4 B3 13 EF 76 54 5D D0 80 D0 32 AF 6E 5F 57
 32 14 0E E1 3C 1D 70 6E 3B 26 23 85 00 36 65 86
 EC 91 5A E4 94 FF 84 F7 71 78 8A 7A 45 32 12 39
 E3 D5 BD DF 4E 4D 2A 0C 4F 4F BF E6 0C 67 FC 3D
 FD 26 9E 64 31 3D 1C 88 C1 A3 82 E3 00 C9 96 B1
 77 C5 CF 9F 77 7E FF E4 29 73 9A 1A F7 C3 23 F7
 7A 57 8F 90 9A 20 17 B4 E2 3F 3F 55 AE 8D CA 1E
 FE E1 36 86 A5 98 83 41 BB 5D 6D F0 C2 29 DB F6
 58 D3 CD 8A E3 69 27 96 D8 92 C2 9A F5 16 F7 DA
 2F 50 39 79 23 97 13 3F BF ED DA BF 2E 9F 46 99
 86 D9 A7 75 D4 CE 3E 5B 0D 4D 1B 78 DF D3 1A 7A
 54 F6 A8 4E 74 90 98 70 E1 CF F6 9B 4B 4F 7F 44
 AF 5C 06 1A 43 28 B0 22 99 A6 07 08 07 ED F5 FA
 0F 64 B4 63 D4 FB 99 4C 12 B4 9E 51 5B B2 BC 16
 73 2F 32 A1 FD 80 2D B4 2D 89 DD C8 62 57 8C FF
 61 EE C2 1F DE AD 3B DE 25 09 EF EE AB 0E C2 DA
 14 77 16 71 86 DA 6B 40 63 7D 10 A6 2C 6F 7B 67
 CC CD 75 05 75 B8 85 1A B8 06 86 70 62 44 1B 81
 76 08 76 06 DD CF AD B7 5A 3F 10 61 4A 12 11 7B
 C0 5F 4C EF 68 AE 6F 43 9E C3 23 5A 5A 10 8E DD
 8E 8B 88 B8 FD 3A D8 60 99 50 3D 46 13 FB FC F2
 2F 09 76 01 51 06 C7 41 CB 8D 5C 86 32 60 A2 BB
 3E 6F 7C 16 D3 84 0C 16 8B 97 BD F4 3A 3E 51 FA
 F3 1A 2D 2F 8E F2 D4 82 2C AA 7C FA AE 81 F5 32
 B9 45 56 7D DE 0E D8 3B 35 85 8A A9 8C 99 C3 C4
 EA CD 7B 6F FC 35 5E AB 79 DB 66 35 14 A5 95 31
 61 1D F4 C8 E8 3D BC 58 26 71 ED 91 74 B4 65 5D
 0B 44 DE 09 55 16 29 8C AE 49 64 6E C9 89 1B F7
 C4 F7 ED BF 51 D8 7D B7 AF 93 25 8C BD 85 79 C9
 C6 FB A9 00 D7 51 02 4E 99 94 FA F1 3B 4A 01 3A
 67 DB 69 E7 9B FA F7 9F 62 5F 2A ED 15 EA 72 91
 F1 EB 97 FC 0B 3E 36 6A F6 85 32 21 E0 30 DC 4C
 84 25 11 B3 0E 81 D3 93 1F CC 8D D8 73 F2 C5 D2
 22 EE A2 78 75 1D 5F 10 F0 B8 C6 36 73 41 F2 AE
 EB B2 A1 0E 4D EB AA 2E 08 63 A4 87 76 27 69 59
 E8 4C E0 29 63 61 20 BA 39 CD D4 D3 B7 32 C2 58
 31 87 A6 18 2A 6B AA 03 15 F2 D9 65 DC 3D 3E EC
 B6 44 18 91 BD 17 98 A0 74 05 BD CD 7A 93 77 C8
 12 94 E5 24 CB 88 2B 34 8E DB C8 7C 12 F5 A7 56
 E2 1C EF A3 86 4A 77 A6 3C 2F C6 4F 13 C6 19 C7
 A2 7B 81 C2 CA E6 30 24 A2 81 F8 1D A0 8B BA 4A
 C0 CC A4 B5 14 FC D1 C3 BD C3 A4 FF 30 E6 2D D9
 F0 D7 87 17 71 D9 D4 34 6C 75 7D C1 5F D0 49 39
 52 A9 A4 EC 27 B0 A1 F2 4D 80 D9 7C 21 CF 3C A2
 8B FE 1C D3 30 2A 70 5F E6 A4 8F 3E 86 B6 E2 AE
 C2 5F 39 A6 EC 1B 09 C9 2D AC 7F 5D 7C 67 DF 45
 68 F9 F4 0B C2 59 12 FB FD D0 33 85 F9 E4 39 65
 51 9E DE 8E 84 D6 42 19 AA 75 B8 BE C6 C9 E8 84
 FE 36 D9 42 09 E1 89 BB B8 5B 38 9B B8 2A D1 09
 B4 8C 23 27 55 9E 1E D1 4D 6A 57 54 2F D0 E5 5E
 53 98 3B 23 98 0B F7 79 21 11 25 DE 6E 8D B6 7D
 AB 4D DA 77 8D B0 36 25 88 12 2C C6 5B 51 FA C5
 41 B1 BA 9D 20 96 40 22 4B B0 BC A7 5E 2E 29 C5
 E3 3D 1C 7D 89 39 47 95 E1 2F 41 B4 1F 8A 88 3A
 3E B3 B1 83 FE 4E 34 98 81 DD 4A 04 E5 52 7A 57
 53 B3 98 CD AA 29 26 3E 38 B9 E0 59 EA 5A BA F6
 4F 63 4A D9 0F 1E 96 7C 02 05 51 D6 EC 00 73 F4
 CF B8 55 39 21 DC 8F E7 56 30 40 C6 E3 49 F6 9B
 70 2E 59 07 F8 B1 D5 3A D7 D5 F0 C2 ED B2 BD B0
 CD 5E C1 B8 7B 9C 18 A7 7F 6A F3 BF 0E B3 AB 98
 5D AD D4 44 79 C3 02 D3 82 91 AF 73 35 FF E2 1D
 CA 7B 4F A9 98 0C 45 35 D4 C0 C2 6E 71 39 A0 D8
 7A C7 0C EE A7 E7 96 BD 7E 93 2A B0 59 12 27 47
 39 38 C9 57 7E 39 2A E0 1B FB AE C5 E8 BB 7F C0
 0D 72 2B 77 C5 17 A6 D5 D8 68 38 77 2A 01 5F 63
 83 C0 EB 79 E2 05 52 91 D5 4D 78 E3 B8 87 B9 F1
 94 CF 17 82 80 38 A8 A9 43 55 12 4C 4D 4A 51 84
 FF 8A 15 35 E7 CC B3 16 52 D7 52 D9 A6 9B 1E 77
 FB F6 95 AF B0 9A E2 12 F9 8C DC 69 26 DC 37 4B
 9E 54 07 11 E7 43 9B E3 7D 8F 50 7C E0 DF 24 DF
 1E 23 0C 19 35 FA FD 82 BE 7E 66 4B 1F 24 A2 21
 CB 8D E7 F6 9F ED 39 4A B4 AE 8E D6 E5 28 BD 1A
 12 88 F5 BB 4F 59 44 EB CD ED 4E DF 4F C5 1D 05
 E5 50 89 50 85 EC 9B B5 67 EC DF FA 95 81 81 C2
 0D B5 EB 9D CA DA 1C FA 36 7C C4 44 92 D4 DA 04
 13 D4 3B D1 A0 88 63 6D 80 77 92 D2 32 C5 7C CF
 ED A5 E3 01 8A CE 39 C4 08 5E 7C 1E 77 1E 8C A5
 8A B9 41 56 2C 46 29 AF BA DC C7 B0 02 E3 E9 78
 E5 03 A9 3C FC 0D A3 0A 61 1C EA 1F FE CD 66 86
 70 88 6F D3 EF 38 37 F1 24 5B FB 8A CA 27 B2 A3
 A5 7C 79 4E 05 F8 63 6D 51 37 0B 2F A6 50 E3 5F
 C9 0F 67 96 06 9E 72 A6 66 CB 8A BE AE 70 0A 09
 FA BB 85 28 29 D6 D9 FE 81 B2 25 DB 83 35 F6 E9
 41 5E EF 4E 4C 20 36 35 74 2D 37 54 50 11 3A 66
 00 E0 D7 4D 3A 26 47 36 BE 95 35 73 CE 81 7E 6A
 64 14 66 16 ED 1A CB F7 9A 65 57 56 C7 A4 AC 80
 79 D7 DB 69 D4 65 AF 0C 20 24 0D 0D EC D1 C7 61
 B5 2E EC E2 B6 09 24 09 98 0B 10 5B EB D8 A1 04
 DD 3F 1B 38 8A 8B 49 E5 C5 8F 22 D0 04 B7 42 02
 B8 34 86 49 BB 81 D3 B7 41 8F F9 C9 1F CC D0 62
 B4 98 A0 12 E6 85 F5 38 E6 C3 FB EE 14 13 E1 DB
 FD 08 F0 EC 1F FB 28 89 9D A9 18 D9 45 48 F5 22
 33 65 02 C7 7B A8 39 26 C2 97 F6 1D 05 7B 5B 3C
 2D 38 FC 17 2D 3F 83 3E AA F1 52 1C 83 74 22 87
 54 D7 98 86 5E CE 10 48 AB 8F 3C AE D5 F9 D3 A9
 BA 0F 5D 15 0E B3 6D A7 F6 20 E9 60 9A 2C C1 B8
 DC 36 E8 9F 9F 84 BE DA 5A FE C9 FE 09 C6 C5 03
 AA CA BD 5B 32 D4 73 E5 1B 0E 19 9F 7D 6B 77 32
 BA 71 1D 19 F9 12 29 15 9E F2 6C A2 D5 66 49 27
 C2 08 47 EA AA 46 75 CA B8 0C 59 83 69 6A 0D A8
 4D D0 CF C2 E9 1F 1A 31 DB B7 63 A8 CC 3E 59 22
 70 E5 E5 26 50 0E B9 28 D3 F4 9D 44 6A EC 19 4E
 C0 B2 A1 7E 94 1E 72 2B CD 44 3C 5A 1B 74 22 B9
 0E 52 F8 2C 8A C0 9E 41 C1 FC 71 8B C1 B7 E3 4D
 0D 0E EB 39 50 09 1C 01 10 91 10 3D 15 3E 17 FF
 69 9D B6 1A A8 43 19 2F D3 C7 15 5F 74 B9 5C 34
 B0 D8 3E 5B 1D 37 A3 A4 C4 43 E3 40 89 95 87 5D
 63 E6 98 94 5C 0C 07 07 82 F1 47 13 0B 95 26 DD
 53 7C 1D E2 8B DA E3 10 80 A6 8F F1 9A 91 C4 ED
 DD 42 50 6A 60 F7 AC 46 3E 4B F8 E8 54 7F F7 32
 EA 1D 7F 70 4B 4D 55 61 45 86 21 F8 32 3C A6 82
 51 06 55 50 3D A0 77 87 23 CA AD 06 68 20 7C B5
 57 08 23 3E 09 55 93 FD 3C 94 10 AA C2 B9 BA 10
 D8 40 9A EC 7C A6 CE D9 83 9D 8F E1 D9 5A AD DD
 38 0C 87 B5 50 DB 83 7F E0 C2 DB C3 4A D9 F5 24
 49 E8 15 76 B0 63 A2 B8 DF C4 D3 6D 61 20 5A 8F
 AF 00 0B 07 F0 53 A6 3C 0F 16 EC B5 09 1A 68 7C
 94 E8 E1 A6 97 57 0D A0 CA 2A 1C 2A 14 F3 CB 7F
 67 A5 CD 87 BA AD DE 8C B7 CE 49 BB 21 95 09 93
 C2 79 20 42 E9 48 7D CA 14 B9 2B 8F 29 27 81 B6
 53 C7 CB 70 B7 EE 95 AF F9 93 93 65 3C 04 CD F0
 B5 16 8D 63 76 8F 01 23 C0 A5 B3 1A B9 67 EB 2D
 33 E8 51 1C DC 83 C0 F6 1D 74 BB A7 72 FC B6 85
 F0 4D 06 8F 5C F1 80 B5 EB 4D DD 2F 0B DF BE BB
 34 46 B8 B6 0C 27 DB E4 B5 BF 28 36 FF 48 C2 BB
 37 76 5B 3B 72 36 34 72 95 C8 6A 06 63 CB B8 74
 4D 3B 84 BD CB A8 24 3B E0 5A 35 63 02 0F F9 88
 05 A3 6A 2C 23 D7 E6 A2 9D 00 F6 23 8D 7F BD A0
 49 F6 B8 83 1E 6A FF 1C 1E 57 29 57 2A 30 1D 5B
 4A 29 BD 50 15 A2 5A EC 21 4E 74 1C C8 21 46 B4
 78 F9 8F 16 6B F0 76 38 07 CC EA B3 D3 E4 00 F9
 CD DF BF 2F CB 99 9C 33 8C 01 5C B1 58 68 96 CC
 23 3C 4A 8C 3F 05 03 6D 9A 3C 9D AA C9 4D AF 41
 85 F9 3B B9 7E FF A4 2C FE C8 15 8C 4D D1 CE F8
 B2 59 56 2C AA D1 7B 98 38 35 58 C6 3F 54 CC B7
 86 DA C0 72 94 7A 0D A4 2B EB 86 60 0C E6 1F A9
 BB CF C8 C4 9E DE 96 D5 5C 40 DF 1A D0 7E 0B 1D
 04 65 F3 D5 5B AE 5D AB B0 B6 45 15 1D 96 98 FE
 6D 2B D6 B9 B0 6E 3D B1 2D DD 6A 48 21 DF 2A 15
 B1 AB 4D C6 A8 42 0F 0E 12 FF AC E7 B7 21 E4 06
 13 26 25 BB 59 8A 20 B9 80 42 3B 2F 2D 16 7E 63
 2D 43 97 3F BD FC BE 22 C2 AA 01 E1 BF D4 C1 48
 21 29 00 D8 6A CC 83 C0 2F D1 FF BA 5F 9F D9 73
 1C A7 16 55 5F 82 98 4A C8 7C D8 0E B4 F4 EA E6
 18 9E 2F 83 59 99 E2 90 42 08 04 C7 24 C1 3E 6B
 1C 0E 6C 98 06 C7 02 CF 07 74 AD A0 DD 85 BB 9C
 94 24 16 B1 02 52 3E 09 D5 A9 E5 88 5D 43 12 56
 77 91 F7 7D 23 25 E7 84 C1 26 DB 6C A4 A5 93 BA
 A1 26 07 94 9B 40 CE 9D 4F F3 20 F3 6E 35 66 CA
 BA 81 16 4A E1 F5 77 5E E0 6F 2D 74 E3 E2 28 0C
 02 41 3D 49 60 8B C1 43 E8 6A 3D 50 1D FF 01 D2
 11 19 03 60 A2 8F 80 F6 F7 59 83 A1 66 21 C1 EE
 29 9C D6 23 F7 D5 68 EB 23 32 E1 1D FE 0F 80 E5
 9A F3 8B 14 63 15 29 9E 1D 42 CB AE 09 4C CA 8E
 DB 76 A5 5B E9 CD 0B 56 EE E4 8D F7 D5 99 F8 42
 BC 50 68 D5 18 ED CF 37 B5 7B 09 B9 C3 06 CF 76
 E5 4F 6B 98 72 EA F2 B2 E1 3D FA E8 FE D7 2D 25
 16 C4 89 C5 3B FF 99 F0 3C BF CD DA CD 3E 68 49
 DD 7A 1F E2 46 1B 8F E3 40 31 69 D6 E4 E6 1E 9F
 06 6F 59 90 A9 BC 48 BB 2B CC 0C 10 06 B3 AC 15
 15 64 04 80 7C E0 1A 76 13 44 09 7C 03 2F 19 BF
 B6 75 68 7E CD 9B EF 49 58 07 30 78 3E 74 1B D5
 D5 BE 1E 4C 53 D8 2B 49 8F 46 B6 F6 29 E3 C8 E2
 85 E8 8C 37 D5 19 07 BF 40 59 BD BE 45 EE 31 DF
 AC 77 D6 02 12 59 72 54 FC BB AC 99 20 2E C0 7B
 B3 62 7C FF 83 9B 69 60 CA C0 59 B8 4D 60 27 40
 4E D3 45 E8 78 4E 32 05 F6 D4 F2 3B ED 6F BB 20
 55 06 06 00 21 8A 08 96 72 B3 76 E6 B2 75 EC 9B
 C7 12 4E D4 38 E5 63 59 DB 02 CC 4A 87 7D C1 56
 6A 7E 7F 21 B5 8E F9 36 0F D2 D4 26 36 BB 83 6B
 1F E5 8D 67 AB 36 6F A4 B5 E5 B0 FE 45 60 29 4C
 AB 43 D6 2E E7 13 D4 77 3B 55 4B 4F 6E 1F E9 52
 22 BE 46 C7 7C 08 40 1C 0F 4D 5A F5 61 55 6C E6
 61 08 21 0E 75 B7 00 70 CE 9D 74 C3 24 5A EA F2
 1E AB 6F 8F 7A 22 5D 64 B6 33 77 8C E5 EA D2 FD
 6E A7 5E 80 C8 0D 43 7F B7 00 39 CA 02 A1 93 0E
 5C 74 AF 86 37 DD 9B 7C C0 43 D3 1D 5C F5 0F 0B
 0F 25 7E DC 1B 6F 65 40 3C A3 D3 A3 DF C5 70 8C
 69 5A 51 27 FD 50 B3 5F 05 86 D2 85 9B 61 D7 9B
 8F 66 FD D9 53 4D C9 12 E3 A0 15 DC D9 43 72 4F
 53 C5 E4 7D D8 E9 72 63 E3 B3 38 B9 8C 19 FF 19
 38 5B D5 A2 93 0A 07 ED BD 58 B0 C3 06 C6 FE D8
 F0 E6 70 33 1A 37 8B F9 DA 4B 47 C5 94 07 BF B7
 00 8E 36 F7 C2 78 71 05 2A 66 88 12 A8 C2 84 32
 B0 34 53 51 C6 E0 F7 26 B1 DA FB 5A 57 93 74 73
 94 0C 28 8D 6F A6 56 3C 7A 6B 7D F1 C2 67 12 70
 0C B4 40 EE 17 A2 5C 79 C7 E8 04 E2 3F 4C EB FC
 3A 6C 3A 94 EB AE 26 7B 3B 27 59 61 1C 90 F0 A2
 3B 57 55 83 49 FF 80 85 24 0A 1C B8 76 4F F2 EF
 AD B7 83 D1 1D EF 96 86 2A 70 51 66 CF 98 D9 E0
 54 1A 65 5E 18 53 C6 BB 82 E1 5C 7E C5 FA CF 17
 F5 D4 4C 17 2E 7B C4 2E 84 0A ED AB 02 0C 44 5D
 70 1D FE 14 EB 2D E6 E1 48 C9 01 FA BF AA 2E 6A
 A6 36 D5 E6 72 1A DA D0 6C E1 19 19 2F E5 5C 28
 78 8F F5 7C 9C 8F 75 B6 F1 62 C0 50 08 6E 57 A2
 CE 50 CF 34 FF C2 94 AC 22 85 C4 4C E7 06 B0 63
 AA E7 1B CA 16 A3 B4 8E 03 F9 23 FD AA 85 36 4C
 B1 BE 8F 2A 4C A4 E5 63 AB 22 10 FD CB 7E 7A 04
 AA A1 63 4D E5 6F 47 22 BB 07 83 FD 1F 08 47 99
 37 CD FA 96 4B 0F 39 E8 17 42 B4 58 2F B0 F0 25
 09 29 4A 7E F0 B6 FA 1E BB 94 0A 80 D0 4E 4A BD
 79 5C 8C DA D3 01 C6 BC 24 BF 7C EB 6A 74 88 A4
 AB AA E2 58 05 34 47 4C A3 7A 07 7B 56 4A 77 8C
 C0 AA 5E 18 39 24 E0 F7 4B 24 E5 B1 19 C3 3D DD
 A9 FF D9 70 30 F5 E1 64 D6 18 ED 8B A8 66 F2 8B
 AC D8 29 83 8A 7A F6 00 EB 54 6C F6 4C 8F 03 B6
 1D E2 3F 2A CD 4B 52 7D 29 10 5B B1 BA 39 84 5B
 DD 2E 5D A4 9B 60 22 CE 6F A6 F9 40 FF 3A B5 3C
 60 8C 7C 3A CE 71 99 47 08 F5 7D E0 E3 E3 C2 93
 8F 1B E2 22 C4 FD A3 D6 CC 47 34 13 10 41 2B C4
 31 B5 ED 1A F7 18 B8 0D 35 8B 5E E8 9D 54 73 BA
 21 04 66 19 B9 E5 99 3F DB AD 91 6B DC CB 07 86
 0D 26 B9 63 4F F1 4F A0 75 93 27 5E 7E 7C B0 3E
 0B 9A 54 65 D3 34 ED BC 30 78 1B 5A 83 3D 80 D5
 E4 98 B7 D1 D0 B2 EE 02 AF 10 19 76 00 14 CA 53
 92 45 F1 69 28 7F EC D7 2E 42 D9 50 ED EB A3 97
 39 E5 51 C0 EC 61 9C B4 0E 40 FC F6 75 C6 90 15
 44 36 56 F4 73 EA 55 2A 42 53 F4 E1 21 48 5C 6F
 37 27 99 3C 1D 03 7E 3B 3E E2 18 2A 97 BE E4 4E
 C8 4E F2 5B 5B 1D 0F 3A AF B3 BA FC AD 51 AE 11
 AD 15 7D 3A AE E4 5D 79 E9 26 B0 94 84 E0 9B D3
 3F 8B AF EB 82 FB F0 4F E9 1C 36 1D A3 CE D4 0A
 FD 73 68 32 26 A7 CD 6D 79 88 9D C2 C5 84 A6 B4
 FC 14 77 56 41 F0 60 2F 58 33 39 9D 45 3F 4C 4A
 78 97 AA F3 4E F7 30 6E 83 50 E7 15 D0 48 88 43
 5A 3A 5D 14 D1 44 32 79 E9 D7 DB 02 58 E1 54 23
 7C 91 55 B6 27 78 B2 B2 06 DA B8 D0 26 36 49 2F
 DE 89 A0 7A 4E 2B 38 81 E4 16 4D E4 DA 4B 36 46
 42 FC ED FC 11 6D B1 48 AF 99 C1 7E 90 26 2D 9A
 7B DB 6B 10 AB 0B E6 A2 84 5B 54 35 D4 9C 78 BD
 68 8C 9F 0E 0B BA AE 95 91 C1 BD 85 85 3B 23 6F
 D1 04 25 B6 DD C0 46 F3 6D 23 68 3B EC EC 4E 63
 F0 81 2F AF D6 7D 5D 84 95 48 05 DD 88 A8 1B 7C
 28 36 AE BB F6 9E 09 9C 32 F4 A6 74 25 52 25 CA
 36 EC E7 F2 56 1E 85 74 B6 47 BB DB EC A5 62 E9
 86 D3 1A 3C CC 7D C9 60 43 A7 E0 EA 56 62 06 3C
 DE FF 5C 5E A9 87 85 44 AA 05 6B B0 90 CA 09 DE
 DC C9 40 90 AA 0B 10 69 2F 55 7A 5D 75 8A 49 A1
 99 FC 4D 5C DC CE 3A 1C 1F 02 8A F0 72 18 EA F3
 E4 D3 9E 4D FD BA 40 B2 A9 29 63 19 0E 34 F9 89
 DD 1B 35 29 9C C4 3D 26 89 92 73 28 AE 71 FE 6C
 75 3C 34 36 95 94 BC A8 48 A7 55 A7 96 88 3F 51
 3C 32 C8 85 8E 03 43 79 90 E5 DD B0 49 73 53 CA
 49 51 F0 2C 91 18 4D AC D3 68 C2 91 D8 A4 D5 A3
 22 94 25 61 1D 35 35 67 FE 4A C0 0E 4F C3 78 1B
 E9 24 4A 0E 0B 5B A9 EE AB 2C 8D 09 CB AC E1 BE
 16 8D 60 7A 63 00 E4 AF AE 58 EF 97 21 9F FD 8E
 3B 4A CB CC 13 B4 A6 0C 43 C7 97 9A A7 A9 8D DF
 9D F5 D4 18 76 7C B0 5E 52 DF 62 B2 B4 72 E2 AE
 25 D2 9F E3 19 D3 8E 97 2F C0 C2 80 A7 ED 82 5A
 58 D0 DA E2 AD 47 DB 63 15 29 86 37 81 82 94 19
 66 E1 ED BE 24 DA CD F1 2A 78 A4 FD 98 F7 2B 64
 A6 46 5A FC BB C8 BB D1 21 C1 F6 1C 88 16 3B F1
 3C F6 D3 20 5D F0 74 3A 58 C3 2A 68 45 BB 77 D0
 CF 63 A1 61 E0 C9 2A 64 58 55 12 35 87 2C D5 EB
 55 C4 84 8C 0D 23 1A F6 D1 15 95 AE 99 73 40 32
 3E 16 D0 66 7B E6 C4 E2 57 EF BC 8D 89 99 9E A1
 95 83 CB 7B 75 71 25 5F F5 4D 70 54 4E 3E EA FA
 32 9E 82 B6 25 3E 6E 8E ED 85 65 8B E6 C7 0C 04
 34 BE 81 C3 25 A3 C0 FF C0 55 FB 41 77 F7 AA 3F
 99 23 FA FA 33 3D 4F 50 90 DE 60 FE E5 F8 C6 C5
 FD 75 D1 B8 03 46 77 87 A7 BF 4B A1 29 7D F5 A9
 12 8A 2A D5 EE 51 80 8F 2F 17 8F C7 05 74 1B F4
 8A 56 0A 4E 41 D8 DB A0 AB C7 CB A0 C7 E9 F7 83
 5D 35 14 F3 98 58 9C 5D 6D F9 70 4C 7E 73 D2 F5
 CA 95 17 88 E2 60 9E E0 84 0D 08 E6 C4 3A CA B8
 E2 C0 A6 5E 43 8C A2 BB 46 A7 C8 25 48 99 2D F4
 08 79 9C 5C 8A 11 46 6C 92 9F 08 FA 31 94 2D 41
 66 D6 69 A3 E6 49 68 65 33 2B BC 64 46 46 4A 81
 4A 11 33 90 DE 94 D7 45 C8 E4 51 D6 B6 9F 6A 47
 FC 00 AE 61 68 BF 41 C7 49 6E 02 0A FA 77 DF 12
 D8 86 9F 3F C1 7B 07 FC CC 38 9F E6 09 87 94 CB
 DF 75 3A 27 AF 32 35 19 E1 01 64 91 D7 89 D3 F0
 2E 8E C7 56 A1 FA F9 3E E9 4D 4D 55 B5 8A F3 C8
 EA 99 76 51 8B 77 98 4B AE B2 4F 89 8C 88 4E 80
 24 68 5B 84 FB F7 94 56 67 A0 DE 02 D6 E1 74 0F
 F0 B6 6C E7 90 A5 6A 01 8D 54 D6 62 8E 59 28 59
 35 DC 64 EC 98 3D A1 11 F5 F4 A3 3B 2E 3B A4 EB
 3A D5 2B 7B A0 E2 C4 7D 68 7A 63 37 6D 89 F7 5E
 C2 AD 17 10 D5 37 83 92 D1 A3 26 77 A6 F9 CD 7F
 3C 9B 02 C2 E4 F1 00 4E CC 68 85 B7 9E 2B 4E BB
 07 D3 49 02 EA 82 F0 16 A0 14 80 70 19 3B DE 4A
 DF B3 B8 AA B4 56 90 47 37 D7 26 C8 B5 14 94 9D
 E5 5C 5E 49 A4 31 9B 2B 4A B0 0E 2C 8F CD 8B 10
 6E 68 8D B6 ED BF 46 F0 A2 36 13 0D 01 F3 42 BF
 06 8B 1A A3 4D 4C 28 38 A1 0C 94 78 D5 5F 2B 43
 6F FC 23 E7 8D 33 63 BF F5 47 C1 53 6E 83 6B 70
 5D AD 15 D4 AA 50 FE 9A 4B F5 38 B1 6A 17 6D B5
 64 50 E4 13 5B 74 EC 9F 0A 89 5F 32 8E 62 B5 BA
 38 8C 37 0A 83 30 24 86 2A EF 5D 60 21 7F D1 25
 DC E5 C7 8A 9D 31 F6 94 64 F1 C9 B9 F8 5C 1B 16
 7A 0F B4 1D B3 03 CE AE 92 94 AD 76 BB A7 C2 70
 AC 1B DC A7 1F C6 47 D4 F4 80 38 86 1C 1C E3 81
 22 AC 56 21 91 75 12 1D 9A 68 33 68 12 3C D0 9C
 D3 3C 37 24 CE 68 1F 1D CF 0F EC 55 A4 02 73 5B
 A5 16 E0 4E D8 E2 C0 97 55 06 0C 83 A5 84 1E 44
 36 9C 2C 62 56 8A FF 41 8B 24 7C FC F1 F8 5E 37
 72 09 18 D2 73 69 02 47 53 82 65 8A 1D A1 80 63
 53 99 CE 63 0D 4E 14 FE 16 F7 E0 BB 09 AF 6A 17
 B6 A5 C4 34 C7 45 6C 8C 52 46 1F 8A 03 49 43 26
 AB D8 41 53 66 0F 8B 06 5F 2B 49 7C 1D FE 91 47
 A9 A9 88 3D 57 B5 8B C1 FA 39 75 AE F5 60 8E 94
 58 C3 94 94 F6 BF A4 22 AC 98 BD BF 00 43 52 D9
 67 63 3D F7 B4 E1 84 84 F3 9A 1A 59 28 86 C6 B4
 3C EE 61 A3 6D C9 B0 69 E8 57 40 3E 94 90 18 35
 A5 9B 27 2A F1 DD 3E 13 46 25 6B FE 8F 83 D8 D0
 F8 C0 79 91 F6 70 06 91 EC 6F 33 CC 21 61 52 CF
 61 4A 7D 3E 3A 1C 57 FF E4 1A 22 F3 77 5D 10 E3
 3F 24 15 CE 9E E0 15 BA 28 FD 32 A1 11 49 40 91
 34 54 47 40 66 DF FD 9A EF BA 69 A5 F9 B9 C5 31
 0C B7 56 F5 3C B2 0B 08 03 3B 5F 57 4C 7B A6 0D
 C7 F4 0F 05 6B E1 85 4C 71 52 AA 15 2B 1B 54 C0
 FB 41 8E 25 79 B0 CB 7A 9F 98 8F F9 7A 2F 54 04
 D8 6B 14 E1 36 C5 36 DE A2 E7 B7 BA EF EE 9E EE
 28 AB 0D F4 22 DD D5 A9 9C 7F 61 89 CC 8C A6 AC
 93 94 D4 C6 46 62 C8 C7 57 7F 84 D7 CC 5F CA D4
 69 CF 08 15 6C 32 12 DF CC 80 DD 48 2C 3C 57 84
 F0 AB 91 C2 4D FA 56 26 05 7C 0B 29 17 42 82 97
 58 9E 25 6E 5B 35 C2 F1 7B 18 6B 77 60 50 67 CA
 AB 99 66 44 CE C3 8E 0E A0 95 C9 E8 17 D2 39 9C
 81 10 ED 9D 43 82 8A 48 5A C7 70 36 AD 37 22 B3
 85 04 CB E8 E3 2C 6D 58 30 A7 0E 7A D6 3D 98 36
 D3 10 57 84 F3 27 6B 8E 81 0B 33 82 7D 3E BA 60
 7E EA 63 AE 5D FD 4F 05 0C C6 1D AC 52 56 E3 40
 8F 10 D8 2D 4B 00 A8 76 71 00 19 85 C2 E9 57 77
 BF DC 70 D8 C3 D0 76 BD D3 BE 5B 1A A5 DE 64 C4
 37 8A C7 D2 B2 94 48 91 DB 34 34 50 E5 E6 36 BB
 76 FA 85 4F 7F BA 76 E5 06 60 46 3F EB D4 44 B3
 C4 E7 9F 4F 62 67 C9 DE 70 68 BA 31 C0 8C F1 4E
 A3 6C 67 E3 6B D5 AD 37 0F 0B 50 05 EE 5D 98 04
 24 B7 35 35 2E 4A 8C 55 2D 1D 61 C5 FC 35 C3 0B
 C8 EB 76 D8 4A 40 F4 B1 B0 65 0F 77 2D 9B CE 38
 C7 D8 80 86 9B A5 EB D2 FC 17 3F 5C F9 9F D0 70
 07 50 C5 AE 07 D8 71 78 B7 96 E4 22 73 16 52 31
 AB 74 8B A7 38 DF BE E6 DF 28 BB EE E8 61 04 76
 B5 9B 9A 30 C7 49 5F 63 96 58 1C 75 5E 46 5F EA
 EA 65 F4 F8 10 4F 8D 1E DB 14 F5 E6 2E C8 FE 23
 40 EE 9F 4A 69 F1 1E 7D 97 22 AD E6 BB 05 FB 0A
 56 83 C1 45 55 BF D7 37 DB 14 19 40 86 92 C3 7E
 AF 3D 36 0B 8E CA 3E 6E 95 DF 81 DC 02 5F 83 07
 01 BB 58 EC 4F 4D B7 6C BE B6 07 E3 D5 5C D8 69
 5A D3 19 1E E9 56 4F 6A C5 12 B6 EC 5D 47 63 D8
 5E 1B 92 3B 57 D2 CA F5 42 A8 99 2D C6 D9 74 68
 44 6A 38 E2 FB CE 0F FF C9 18 87 3B 83 03 D0 D1
 12 BA 19 E0 39 EE D9 73 39 ED A7 56 0A F1 FC 59
 9C B2 38 B0 B4 60 32 D2 89 9A 95 A4 76 DB 10 60
 72 DC C9 4C D6 91 2D D9 7B 69 A7 4F F8 24 E9 34
 A2 A6 9C 57 28 04 98 60 79 31 3C 08 AF F6 D2 20
 45 7B 66 F6 81 39 6F 3E E2 58 A5 79 A3 16 8C 7F
 9B 4E B2 8F F3 42 45 AE B1 97 85 57 7D 11 6A BA
 12 B5 15 A7 FB BD 4F 73 C7 A9 14 60 13 AF 5A C3
 95 CB 04 11 33 90 D1 BB 2A B3 17 14 CA 8A AB 3B
 68 0E B7 C8 39 D0 6E A4 BD DC F2 C4 E6 EF 86 77
 14 0D 7A 0C 01 91 0A 04 F2 49 92 96 60 94 5E EE
 71 AF 86 33 A8 2F F1 FA D7 CA E8 E7 9E EB 65 40
 01 09 27 58 F9 67 9D B3 DC 8F 6F 84 51 2F 8D 6B
 26 6A 3F 22 45 8B 5F 42 CC 50 08 7D A9 FA 22 E9
 71 98 E9 DE C2 7A FC C1 08 D4 83 A9 89 2D 2B B8
 31 D5 FB 0C 33 0B 02 9C A5 BB 10 FC A2 1E 5A C9
 8A 0C 0A 67 E5 36 7A 50 04 09 08 2A 38 AE C5 57
 57 7C 45 DC C2 84 C3 9F C6 4C EF E1 4B 87 A6 51
 CE 8F 07 F2 C6 F9 EC D5 BA 45 8A 85 25 CD 19 8C
 A0 ED E4 9B DC 92 76 01 0D 12 69 93 F3 E5 88 54
 CE 21 70 5C CE 3F AC 62 F1 B5 20 8C 7F 37 E4 A5
 18 BC CD B5 F6 48 31 D7 96 7D 61 BF FC AD 2B C0
 8B 53 99 1C FE 15 29 E9 33 41 82 30 52 4D 57 4C
 F0 12 B9 0E B1 59 6D 09 CB C3 CB 00 5A 95 F3 F1
 59 92 D5 F2 B6 21 BF 90 F2 5D C1 6C 72 A2 E4 E2
 29 4D 62 92 6E 51 EF 3D 24 1E E3 61 5C C0 28 5C
 AD 17 40 F7 99 F8 06 92 CB 6D BA E9 EA 08 9F A3
 D3 17 8F 3D 4A 94 81 3C 3E 63 55 8B EB CD AB 1A
 39 AC 35 73 E4 D1 49 5E 05 CF DD 23 E9 40 9C E1
 C4 12 8C A2 F0 44 11 84 8F B7 6D B2 2C 4F 03 98
 ED 2B 6B 34 97 D7 C3 4B 8C 77 C7 FA 6C 68 CF A7
 23 3F 54 3D 27 B7 30 68 20 E5 3E 04 A6 B6 CE C4
 09 AA 67 AA 34 99 44 06 AF 2E 6F 6F 90 4E B4 05
 87 D7 28 2C 73 0F FB 8C 74 7C 91 D1 51 DD A1 13
 D8 44 4F A1 A7 D2 BA 13 69 00 C1 FB 4D EE EA BD
 CA 6F 50 E2 3A 4F 40 73 55 76 38 BB 71 BF 28 67
 46 0B 98 B4 AC A2 E2 37 24 3F 80 00 36 1F A3 BF
 7B 53 3D 2C 04 75 BF D1 64 95 54 B6 4B 12 DD EB
 25 A8 F8 10 8F BC 87 1A 4D 9F 69 29 86 6A CA 52
 41 84 DA 54 92 07 1F 3B EC A1 96 83 54 F5 0F 2B
 8F E1 32 92 66 1F A9 69 DD 3D E3 36 FC A4 DA 9A
 1D 10 7F D8 4F F6 5B 63 D3 D6 43 51 F8 9C 05 3D
 FE 08 6C 8A BD 6D 7D 02 17 78 6D C8 F1 56 24 C2
 A7 77 5E 20 1E F2 35 D4 A7 23 57 6B 0D C0 56 EA
 85 4D F7 10 1B A9 F8 20 7D 74 86 9A B3 68 1A 64
 EA 97 9F 16 4B DB 1C 6B 8A 50 E6 F5 DD 84 3D A6
 69 3C CC 15 8B BF 12 65 F0 7A C9 4C C4 EB FA 40
 00 13 8F 6A 5F FF F6 82 67 A6 D4 3D 15 38 01 D6
 60 79 22 8E F3 48 6C 1B 47 A2 0D C5 D2 6F 81 3E
 78 51 0A 05 71 5E D4 5D 9C F9 94 32 6B 5D 80 E1
 FA 41 EA 78 3D 48 7D 88 20 91 2C 6E C6 6C 5F E2
 FB 5E DA F1 F6 63 22 39 47 69 61 32 DA D8 2A 05
 E7 77 FF AE 5E DB B3 D6 4C FD 68 19 8A B3 48 CC
 57 1D 1C 8C 75 4A 28 56 A1 34 A9 1D 39 17 09 54
 52 9C 4B BA 60 41 90 17 22 72 B3 8C 53 81 7A AC
 D4 FE F8 38 6F 48 D8 F6 88 DF 41 93 C9 17 D4 BF
 BD 40 0E AD E2 6C 77 61 33 07 A3 56 4C 28 D7 56
 2C 59 73 EC B6 81 F1 66 E2 2C 98 C3 18 43 FA BC
 72 9C 2A 7C 7D 80 A7 EC 73 14 20 E1 14 D4 8C 6E
 8B 6B C3 EB 65 BD 06 5D 9A 40 E2 2E 25 D5 51 C4
 48 0F EA 58 D0 14 52 6B 01 73 98 48 3D 5D 00 0C
 80 AA 5F 08 9F F6 A8 AB 8B 82 9F FD A7 4C 81 CB
 8A AD A4 01 61 85 FA C2 4A EA 48 C7 A8 79 99 1C
 56 2F 34 DA 25 08 52 8C 9E 01 FA 96 74 52 F1 7F
 EE 97 61 37 5B AC 9F B1 19 C1 47 03 E4 33 84 99
 43 43 D5 64 7A F2 42 2A 0C 9F 0B 2E 13 04 C6 06
 4C B3 10 DE 06 7E 30 CE 5F 8D 6A 44 E2 30 D9 CE
 7C B8 51 0B 68 CD 16 EA 6C 38 03 DF 5C 0B 65 94
 6D F9 49 D5 7A AD 3F 00 78 BB 33 71 38 E8 BE 3F
 7A 26 C7 81 02 61 E0 28 23 73 2B D0 40 4F 4B F6
 03 75 E4 70 72 4B D7 B5 EA D1 D5 9F ED B7 9D 29
 93 90 76 43 B7 7A A3 D3 81 01 AA 86 39 E9 CE 72
 E3 68 B6 27 BF 56 7F 61 2A DA A0 C4 02 86 B7 6A
 34 6D 43 5D 77 1A 26 42 23 2E EB 7C 18 64 4E 39
 66 95 98 A8 28 EC B0 AF D8 EC 9C 37 28 C3 AA C7
 58 B4 EA E4 18 B1 51 26 3A 9D CD A0 6F 86 36 BF
 B1 A5 AB 22 05 F8 E5 2F 7F AB E4 5E D7 8A 11 AC
 CB 80 4A D1 E9 E3 4C 19 75 79 7E 19 D5 64 A3 D5
 8D 62 0E A7 93 AB C3 46 0C CA 0F 81 EB 82 B6 6F
 C1 08 86 29 B7 0C 8A 4E C8 53 E3 51 65 04 51 9D
 CA 13 C4 AC 17 07 36 FE 4C 37 67 C3 F0 7C 78 8E
 38 9B 7D 00 38 01 EA 9A 2D DB F0 77 A0 C2 25 F8
 FB 61 84 E0 A6 48 1B 27 83 4E 09 A3 55 90 2A AB
 C0 0B D6 2B F1 52 9C 6F 91 5D A0 FD 45 6C BE 0C
 6E 2B 35 45 A5 5F 3F 06 3B 3B EF E7 55 58 2B AA
 B6 0D D7 E7 E0 68 79 06 92 A4 46 0F 9F A5 49 32
 C2 2B CD 64 12 4E 84 3B 71 97 D9 28 B9 66 29 F0
 0B D8 F5 C1 9E 80 D6 83 9A CA D8 09 C2 AE E7 63
 C2 3B 1B AB 16 FC FA 8B 5D 42 50 2F 94 98 77 EE
 49 90 C8 3A 65 9F 77 3F 65 BF B1 AC C1 EA 10 25
 D9 98 74 EF D6 B7 F1 9D 76 1F B1 58 13 A1 10 80
 26 AC 87 B2 54 73 94 B9 08 FC 23 07 7F 43 E1 AF
 44 28 8D FA 60 46 CC A4 F3 F9 25 4C C3 5C A2 C9
 A0 8E C3 A0 E0 15 43 9A 09 A3 51 1C 92 BC B9 0F
 21 6C D5 CD 30 F0 88 E0 F8 8A 1B 63 B7 C9 C2 C2
 D1 2B 39 83 2A E4 E5 BE 73 A3 EB D4 9F A6 80 E2
 E1 51 4E 5C EA 28 3E 5B BD D1 EC 45 73 B6 5B B7
 E0 49 81 22 56 AA 54 00 D9 F8 D6 AD 58 9C 63 C4
 2B A2 CA AD 79 4F 12 8A B4 82 AE 73 BD F0 84 C9
 E2 D2 B5 F3 27 E3 87 C3 AC 4D 95 2E CC C2 DE 19
 76 99 83 1B 80 96 89 BE F5 2F A5 21 F4 7D 6D 20
 8E 19 AA A5 34 E3 67 40 09 90 1E 24 23 08 5C 7F
 14 83 13 1C 27 5E ED CD B6 A2 CE 10 8B 78 B8 61
 70 F4 7E 2C 46 35 1A F9 B9 44 17 E2 0C CE 4F 9D
 14 40 24 E0 89 34 CD D2 CD 87 CA 57 5D 79 2E 5E
 F2 79 3E 60 05 28 4A 56 75 F4 C5 CA 10 AB 18 45
 D7 8C 2D 27 B9 AA 81 2F 0B 87 1E FE BA C0 DE 0F
 97 8E 12 E8 52 7E 0B B0 49 BD 39 60 5A F0 14 0E
 0F F0 8F 8F 74 BB EB 3A 03 CC A2 F5 6D 0D 81 F8
 44 B7 70 F8 7C 79 0F CE 8F 76 6C E7 46 B7 A6 24
 54 2B 03 09 D1 79 3F 89 66 B2 D7 ED 4C 92 8F 87
 EF EA E4 92 2E F0 BD 28 CE 58 DC 48 BA 52 3B C5
 7F 3D F1 5C 3B DC 88 C0 6F B8 8D FA 4B A0 EA F6
 E3 73 F5 4D 97 1F 55 21 1A C7 A6 59 1B 80 BC ED
 35 E2 FE 1A 43 8A 4D F5 78 9A 1C 95 D3 93 CA BA
 5E 66 BA 25 68 65 F4 70 62 13 F3 2A 79 92 49 21
 35 62 21 F9 5C 77 9B 74 02 E5 A2 84 95 E2 DE 3A
 F4 F5 16 C1 C3 F2 77 8D 58 92 65 B5 96 7C 21 8F
 30 29 FF 88 C2 0C 8C 37 D0 0F 89 B2 08 2C 74 BB
 2C 5E 18 F9 10 E1 2F 01 4F 25 02 FE 73 50 CE 76
 51 26 36 3E CE AE FC F1 77 A0 81 08 8A C7 15 DD
 FA 17 07 66 29 77 D5 AB 55 0F A1 67 76 F7 1E 5A
 73 E9 88 F3 18 E6 FB 05 60 A2 8D 60 A3 BA A0 5A
 A5 3E AC 57 50 89 EA 70 96 B4 1F 45 3C FF 88 A3
 3F F1 F7 09 5A 97 26 64 29 34 40 CF 87 6A 59 E5
 65 29 1F E2 A6 18 A5 B5 C2 16 CC 29 CF 90 00 32
 E2 A0 7D AB 6E CD 0F 01 00 19 4F F9 F9 E2 C8 E5
 CF AA 4F E3 C3 35 3A FF 06 EF A3 4F 62 D8 52 18
 1E 43 7E 3A BE C1 A0 9D AC 78 6D 48 7A 4B 4E 8C
 69 5D F7 CF D8 80 4C 24 4A 3B 34 40 DD C1 41 F5
 4B 9C 9E 06 69 C7 F2 1C B2 19 F5 FE 3E 4F 26 9B
 11 38 C9 70 8F FD B7 31 67 23 B7 63 99 C7 CE 22
 01 D5 FA BB 26 58 3C E1 AE 26 83 A2 2C DD BC 31
 91 40 33 15 8E 89 0E 99 9C 1A A7 32 13 44 85 F4
 AA 35 C1 31 7C ED B8 D1 D5 44 66 11 5D 96 4A 68
 9D 68 F5 C9 71 4B 76 51 7D 27 0A BE 03 7C CC C0
 C0 E3 88 4D F4 86 46 98 21 75 90 62 24 87 F0 31
 00 A1 37 45 E2 C4 57 D3 41 53 4B 0F 6D C4 4A 59
 43 64 BA EB 6A F0 F4 95 92 7D 14 B4 EE C2 C0 C8
 FD D7 37 6F AB 3B BD AC BB F5 42 09 77 4C FA 5F
 73 00 5E F9 07 F2 60 3C A6 45 85 AA 07 A2 3E C7
 F4 24 3E 90 72 6F B3 A0 17 5E C0 4E 35 23 BA AE
 3F 9E 9A D7 36 F5 34 65 74 4A 90 9D 81 4A 50 36
 01 75 95 29 28 F4 63 29 52 AA 5E 80 65 FD 61 53
 77 12 C4 74 FA 7E B9 0D 6B 55 76 24 9D E6 85 81
 9F 1B 13 0C B3 EF 89 57 20 ED 57 E5 89 D4 76 68
 FE C2 2E 5A 93 CE 2C 21 B9 6B 05 7C 0E E7 77 49
 74 6C 99 E5 00 18 82 E3 B6 13 05 83 65 C4 07 4B
 C2 80 C1 65 68 A4 E2 26 98 F8 4D B3 D1 45 93 FB
 BC F2 4F 1F 12 EE 87 DE 76 AD D5 D3 63 12 0C BC
 A1 62 0F E0 F1 D0 41 25 FB 9E 9E 2B 9F 29 A3 83
 43 52 69 91 EF 1C DB 96 F4 9C EA 47 6F 76 6B 90
 19 7A 71 A3 E6 E0 4F CE 63 21 7D 7C C0 B3 BB EA
 AA F9 CD 7B 66 E2 F3 F9 C8 CA 47 65 AF D3 D9 92
 4E 94 7F CF 54 0A 6B 30 33 09 0A 0F 63 1F 99 7A
 F2 0E 29 26 D9 72 24 08 A8 B4 46 61 9F 31 96 2E
 A5 49 56 EF F3 EE 0A B2 E6 81 98 C0 54 67 B5 AE
 FD C2 B9 88 4D FC 34 04 41 4C C4 80 37 EA 17 A9
 0C 9E C3 32 9B C9 7E CF 81 DB 7B 13 BC DA EE 05
 FE E5 4C 6B 95 13 73 04 F2 C4 A5 AF EA 7F 7F DA
 E0 07 AB FC 33 8D 50 08 8D F4 8D 3B 64 83 D8 36
 1B FC D9 11 8A DD BC F6 10 8F 84 DE 74 3B ED A0
 77 88 E2 17 4B 77 C3 9A 9B 22 27 EB 2B 68 4C 08
 4F 53 F0 94 40 1A 1F 82 F8 B4 67 27 0C 0B E9 D1
 82 FF 22 BF A7 5B FA 86 CA 9D B4 3C 41 70 92 27
 6E 66 72 9B 4E C4 44 0E 95 C4 69 1D C9 CD 9C CF
 A2 B3 7A 28 58 97 3F 98 C9 93 F7 35 1D 4A 34 B7
 8F 95 AD AB 83 8F 01 B1 5F BE C6 C6 22 82 72 34
 62 C3 D8 D4 6D 11 9E 9D E9 8A 67 DF 57 6B 58 36
 29 83 FE BA 58 91 52 ED E8 A4 5C 97 6F F2 19 ED
 04 76 AA 11 C3 7C 6A 4A 48 9A 35 EF 2A 74 58 9E
 B0 3F 33 B3 91 A2 D9 57 EA CC FF 49 25 AF 3E D5
 72 79 51 EC 1A DC 6F 96 20 B8 96 B6 A8 A0 29 A3
 E4 EF A2 2B 86 D5 44 1A A6 77 1D 63 36 A4 27 1B
 30 1D E3 70 54 CD 9C 07 C2 3A 35 3F FE 16 1B A6
 EF 90 21 17 8B 0A CC 8F 67 4F 78 CA E6 CC 2E E5
 1F 39 2E 4D FC E1 40 79 49 7F B1 97 28 25 69 2C
 A5 EE 03 D4 53 0D 0E 94 55 94 2B 26 32 4C 34 A8
 B1 81 29 20 E9 AA 83 F8 38 58 AC 2F 16 65 6D 79
 A4 32 AD C4 C1 24 A3 5B 88 D8 FD 2D FC 9B 85 F8
 D9 41 88 E6 6E 31 02 45 7F 5E B7 A7 BF 59 59 3F
 58 DC F3 08 45 6B F7 E7 9D 11 89 24 14 BD B0 50
 9B A1 5D 42 25 E9 42 85 8F 2B A3 F1 2B 2A D8 13
 CD 57 DB 40 78 30 83 6B EF 41 5A E8 3D 3C 0C E0
 69 93 18 65 99 F6 0F 0A E6 99 23 32 3E 5A 99 3B
 D9 71 2A 51 B4 09 EB EA 85 C6 86 CA 62 DF 08 D4
 B7 2C 76 ED A9 F9 65 6D 07 4D 29 3B C2 1A AA 3E
 E1 ED 77 60 5D 98 38 F6 4C BA 1C 06 1A 9B 70 2F
 0D 16 92 DD CD AD 00 AC 61 CA DF 57 8B 9E A1 46
 07 68 6E E1 F0 B4 87 74 61 F8 B1 8E 60 D5 98 CE
 64 59 CE 47 F2 4F 8F E7 82 BE 29 E5 B1 8C CD A0
 FF F1 FE 1D 8D 6B B5 D4 75 87 66 60 62 62 4C ED
 22 E7 C9 81 73 CE 88 95 35 E8 67 B1 B6 D7 86 45
 21 65 9B EA 03 34 C9 76 35 C7 D1 19 6B A2 CE 6A
 88 66 46 EF D3 2D 14 29 9F 5D 78 D5 FD FB 9D C7
 2D BD 5B E3 F5 58 14 14 25 20 46 C7 0F 28 41 09
 64 F6 23 B1 A5 3E E9 52 4D E7 5C 80 93 28 E5 E2
 E4 96 05 33 4A 40 E0 16 3B 16 54 7C 30 6E 15 D3
 61 FD DE B4 A8 B5 E8 A1 2D 9F 25 1A 96 51 96 A6
 11 59 08 C0 59 4A 2C 48 A7 7C 2C 6B 0E 3D 17 A4
 EE DA 83 E8 79 9D 9D 8F 76 A1 AC 68 FE 3C 85 CC
 92 F4 D2 57 5A 0E 2B 2C A0 FA A4 14 79 22 36 F8
 71 BE 3D BB F8 19 EE 7B 7B 1A 88 9F 7D 54 0D 21
 92 71 D1 86 2F C4 16 C2 60 99 43 04 95 18 5C 65
 59 43 A9 D3 93 0C 34 BC 0B 2E 5C A8 F0 15 F9 33
 48 3D FE 48 35 AE 84 77 CE 0F 91 B5 70 3F 60 B8
 D2 20 14 5A E7 3D 08 A2 97 0C C8 2C B1 F4 D7 FB
 AE 39 73 98 70 E0 71 A1 6B DD 74 F2 99 5E FB BC
 D2 61 72 69 3B 9A E6 4B 7C 53 E9 28 29 7F 96 06
 98 16 E4 8B 14 63 D8 5C FE D6 9D 20 7D EB CD 04
 2B 23 7D 61 62 7D 54 3E 76 86 50 AC AA BB CB A9
 C5 41 90 4E 6B 84 6D A8 73 FC C3 3B 31 2B D3 BB
 87 AE 8A B8 E0 9B 01 8E 3A 6D 08 A0 EE 52 BB 87
 80 9B C7 0C EA A8 27 7A CB A8 A2 27 E2 D4 E4 00
 30 FE 56 6F 5C 0F F8 41 BF 16 D3 E0 BC FF 8E 36
 31 C8 25 88 93 C1 1F 7E 90 31 B8 C3 65 62 43 B5
 B5 1D 8D E3 E0 AE 47 7A 0C 4F 5C DA 91 42 76 CB
 58 0D 95 F5 97 0E 60 09 AF D6 07 13 95 2E 5D 87
 FC 07 64 AB 9E 4A AC 16 BE CB 52 E4 53 B1 DE AB
 09 97 C5 83 CB B9 9D 2B 66 31 8C 10 EC 81 A7 0D
 E7 96 0C 5A E2 A6 F0 54 3E A2 8D E2 7B EB C7 B8
 DE B1 6E C3 CA DF A0 B0 E1 74 18 0A 1A 9A AB 8B
 3D 2B B0 37 40 77 3E 32 49 82 E3 57 BE 19 64 DD
 5A 19 17 09 DF D3 93 03 8E 6E 16 E7 64 00 26 7D
 78 80 A5 07 C2 87 76 15 A4 97 F2 3B 61 38 8E 70
 D7 DD 31 28 CC 73 5B 8A F5 D8 0B CE A3 6A 73 79
 31 52 58 1E 71 55 44 39 9A E6 E2 CF 08 56 A1 68
 40 78 CE E9 05 A7 A7 1C 40 0A 58 78 88 62 35 EF
 C4 33 12 AD 3E DD AD 68 E0 15 9D 7B 95 03 5F 34
 7C 1A 48 28 31 B3 86 EF AD 98 C7 CB 37 D4 6E 59
 60 ED 5B B0 51 73 C9 E9 19 73 F1 21 FC 1A 93 8E
 DF C8 60 DF 36 F1 D2 6E 1C 59 A9 A2 90 CC 09 42
 6D 63 6F 42 2C 06 42 9D 2F 0E 2A 5B F9 BD 78 96
 12 54 48 79 B9 D4 C4 5A 55 6D 94 A3 7C 3B 56 EA
 4A 78 86 F8 7D 55 32 ED AA 12 7E 39 35 46 53 18
 30 B1 28 FD 7E 00 51 9A D7 2B 3B EA 52 59 FD C7
 AF B9 EA B4 99 50 C0 C0 6D 69 04 73 3F 89 00 77
 57 A2 8A 28 95 D9 56 40 51 36 E2 B0 0C 55 32 97
 5C 49 EB AA F6 FC 80 1F DA 2C B7 3F 7C 5E 5B F8
 53 45 03 1A 06 6C 44 61 8C A0 8E 19 36 C4 55 DC
 D5 DD C7 D7 8B 2F 4C 90 EB D1 A3 AB 3C 73 42 FA
 61 B7 E1 4E 66 EB 60 E7 63 E4 EB DC 66 11 E4 23
 B7 62 BC 53 46 7A F2 AC 5A 05 D1 76 E1 C0 A4 E7
 70 9B 68 8E F6 3D 3D C0 6F 5C 98 91 DF 36 0B 19
 F3 36 8F 39 11 5A 94 C0 04 C7 2E 16 59 0F 69 E9
 80 CF 08 56 42 27 F5 22 3F 69 0C 91 D7 8B 66 59
 51 A2 15 5E 14 A3 1D 64 01 D2 D9 92 FC FE 69 37
 F1 DC C0 9A 84 77 84 F4 55 4C 09 D1 D8 D7 52 07
 24 7E AA 7F 13 4D 61 72 93 65 61 72 D6 C7 65 74
 0B A9 1A 46 F7 54 63 CA 63 A1 15 22 BD 93 64 1C
 6F 3C 3E 78 71 11 41 74 AD 73 BD 89 36 A2 50 B4
 77 D2 65 9F F6 72 BE 94 21 86 51 BB 12 0F 0B 0B
 DD 2F 72 9E 50 C8 64 72 44 4A 5D 18 2B F7 F7 6B
 DC 94 AA 8D F1 6A 36 6B BA F9 BD C2 94 16 BF FB
 B7 4D 12 95 EB 47 96 73 D2 6A A0 08 EF 96 1A 39
 21 02 05 50 59 5D 04 CA 5A 75 B0 34 6B B6 C8 C4
 82 1C 79 F0 94 4E B0 62 F6 96 6A 06 DD 91 EB 49
 17 47 94 61 49 7D 52 15 4B 09 64 BE 37 1C E6 08
 C2 66 F8 24 F6 A8 A3 C2 6A 6E 77 6E 6D 70 C9 1C
 8B 00 49 6B 68 99 A4 4C B1 9F A7 C5 43 E9 2C 5F
 0D 16 B4 1A BC 84 4B 17 21 09 D6 BA D4 4A 8D CF
 E0 4F 9E F8 D9 D2 30 C2 48 04 74 99 68 16 BD C7
 CE CA A4 64 D7 2A B7 D1 6A F6 D5 15 1B 5C 91 0E
 05 D4 68 53 CF 70 92 23 CE D7 34 4B 93 14 62 10
 85 B0 87 CE BD 48 93 E6 14 C2 48 04 5B 55 7F 34
 2C BF 4D 1E B3 EF 3B 1D 55 E9 A8 FF 39 B6 D2 4A
 B2 FD 3D 88 70 DB C8 2A FE CB B2 76 6F 18 2B E9
 C9 AB A0 4F 53 DC 2F 35 C7 11 14 69 D6 C7 D5 06
 BF 0B 58 CA 32 A6 23 D6 1D AA CC 3D B4 D2 38 5C
 FA 7F D0 5B E7 91 80 A9 09 57 BE C6 EF F2 F6 F6
 17 E3 84 50 43 19 1A 16 98 26 31 89 60 6E C6 85
 B7 77 17 30 57 E9 DD 98 B8 49 AE AC E2 0E 48 B5
 D4 CB 57 54 EE 77 0E 19 34 12 26 C3 B3 64 62 62
 11 EF C0 EB 55 0E 0A B3 31 6B 74 3C 6E 86 F0 7C
 A5 77 D7 16 13 B8 05 41 4F 76 44 21 42 18 69 8B
 6A A1 AC A1 86 DC CA 21 E8 22 B5 A0 AD 7E 1A 70
 93 5F 4C 26 8B 0B ED A4 AF 7C 33 07 1A D8 CA A1
 24 81 42 4B 16 46 EF F4 EA DA 20 92 CB A7 60 D4
 89 76 B8 F1 A0 23 FC 0B EB EA 82 D0 9C 1F FB 4F
 00 42 7A 75 31 96 50 B1 20 F5 B5 95 38 4A BA A7
 99 8C B5 3F 27 12 90 92 93 B0 7D C2 10 04 87 99
 7A B5 D6 94 DA 3B 2B 12 64 0A FA 08 DC E8 32 37
 F7 69 17 F9 E7 76 82 CD A4 DE CD 81 BE 9A C9 17
 D2 7F 6D D6 29 A6 8D 01 2C 2E 83 BF 05 86 1A F7
 3D 05 16 33 CE 05 3B 23 71 70 FC CF 17 4C 02 D9
 ED EF 81 FF F1 99 82 44 84 3B 0A 85 31 7A 52 2B
 D6 84 E6 DD 23 E0 0D 50 E9 7F 7E BA 6B E5 DB 00
 F0 50 67 79 A2 2E E0 DF D3 D1 22 B8 42 F1 BF EB
 44 9A 43 70 02 D7 51 44 77 B7 C8 9A 00 17 59 BF
 44 BF 56 F0 7F A1 1C 57 2B 10 36 A7 73 F9 49 9A
 FA CC 19 99 5B A6 93 39 C8 CD CB 49 7D 70 E6 C8
 2F CF BD 90 7F 2F B7 35 58 F5 18 6F D9 ED 01 2A
 C6 EA C4 9F 0D 64 02 C8 3A 30 5D FB 68 F3 D2 69
 A9 C2 67 92 49 27 EE 11 52 0A B0 68 9E 1D FE CB
 65 C0 A7 C0 61 82 B8 43 BA 81 34 C3 B6 10 42 00
 8C D7 D5 AF 51 BD 37 AF 0D 30 51 01 C5 9C 0D EC
 3B 98 57 B5 1C 54 C7 B8 ED D3 4B 44 13 51 D6 69
 C2 C0 76 A2 CF 13 67 3F 71 13 BD 12 0E 40 65 C2
 97 3D 09 23 90 1F EE 69 80 B7 3A CB 2F 82 F7 27
 3D 83 86 10 B9 F1 33 C4 43 15 29 39 58 C3 57 84
 0C 43 97 4A 81 B8 1D 1F A3 9B ED 57 3D AD DA FC
 F7 20 02 55 B7 48 B5 FC 6C 55 FF 82 15 44 96 6A
 D5 B1 FE 6E 1A 7C 8F A3 34 50 51 AC B6 6B 5E 0C
 36 DA CB 94 1E E3 98 07 75 49 A0 3F B3 34 C2 71
 D3 3A D7 4A 8A DB 01 82 17 FF B7 A5 3F 08 B6 21
 6E 0D F1 FB 21 0D 7B DC 4D AB 07 C6 0E CC 27 28
 E9 33 50 5D 4D EF 30 93 E7 56 39 12 5E DC 07 7F
 90 B0 5F 85 7C C2 24 7D A6 B2 FA 68 46 00 85 D9
 39 7F 05 F4 9B D7 E3 25 73 89 72 EE 06 13 D3 F6
 B5 34 89 AC E5 30 7C 95 32 51 C0 D1 2F 42 3F 5A
 4E 15 69 D9 29 03 48 C0 1B AA B2 9F E7 25 D1 3B
 35 E5 BA AE 92 C8 45 B7 81 C0 ED 2C 5D 4D 34 37
 5A F6 B2 51 D8 15 26 9E 2A C1 E9 0B AD B9 EF 0F
 2F 83 7B B1 20 11 5A 8D 95 E4 C9 5D 50 F9 B0 E2
 A5 42 23 D6 79 DE 76 9F 9D 0F 6B B0 43 AB A5 13
 FB 0B 49 55 83 76 8E 39 12 96 7C 4E EF 89 3A 2B
 FF 6A 43 5A 22 7A 67 B7 3C CF 23 3C 17 8D 62 1D
 34 73 4E 4F F4 CD B1 02 48 94 5C 84 FC 46 79 B7
 9D C5 8F 03 AD 81 25 D4 7C 9A 7B EA EE 76 EE 6B
 F0 4D 51 DD 42 81 11 7D 12 FA 4F 1C 9D 5D 8C 7D
 B8 E5 C1 DE 16 59 9D AF E6 4C 4F 3A 49 02 B3 31
 05 6F 7F 0E 75 6D 03 98 51 90 FF B7 08 12 8C FD
 78 45 28 5B 49 B1 68 C8 63 17 D4 22 55 F9 82 EB
 80 47 AA 6D C1 39 38 85 0F 38 C1 8E BA F9 BC B6
 F6 61 E8 46 84 97 DF 5B 39 0B F1 6E 6D 37 DD 61
 CD 1F 97 B9 7C 86 4F A3 47 17 36 FF 83 88 E5 81
 43 0E 21 9D 63 E3 3B 1B D2 72 07 FD F6 34 F0 69
 90 EE 3D E1 62 E0 AC AC 6A 72 5B 3B 66 78 9B A9
 3F 87 73 DA 29 CC 5B 0C 09 1A 93 32 1D A9 DA A9
 F7 63 E1 E1 E3 F9 E3 08 E3 26 D7 DB 22 50 4C B5
 89 EC 7B 24 A3 2B 48 CA C5 E5 77 99 93 EE B3 F2
 85 4D 4F FA F6 B7 0B 40 EE 9B 9A 4E 98 32 6E 52
 AD 95 41 A1 30 4E F3 1B BC 12 5A 04 06 04 43 E1
 CC 91 D4 C1 BB 47 0F AE DB AA 11 95 78 D0 E4 35
 A5 D9 3C A0 8E 14 B2 41 B4 49 E5 07 95 99 58 02
 A4 F5 64 6F 47 2B 06 92 3C E0 64 2D F8 48 6C B8
 0C 56 F0 DE 78 A5 96 9E F5 59 B9 26 BB 65 16 75
 0F 26 DC 51 91 47 AB 3D 03 CA 6A 1E 9E 56 DD A7
 7E 9C 22 B7 60 60 81 3A 3E E6 47 D3 E9 C1 95 F5
 EA FE F8 51 A5 51 B1 8C 2E 39 74 A9 50 A3 EA 3C
 68 4B EE E7 79 B5 41 1E 94 11 68 BA 38 6D C9 EC
 A5 4A F0 50 4D FE 14 FF 5C C1 4F B8 CC A4 E5 6F
 E6 8C C0 A2 1C 97 E3 02 C3 9C 83 27 54 5E 3C 84
 FF 24 C2 13 E0 2A AE 19 39 9A 3B C1 AD 50 91 DE
 AA D7 E3 21 F4 F3 B8 2A FB 7F D5 C2 1D 37 61 42
 09 2C 4A 4E CB FB 58 69 BA E8 71 BC F7 B2 79 1B
 B4 88 B2 C2 7A 7C 5A 87 84 36 F4 18 20 D8 30 C2
 CF 29 D3 4A D1 58 39 28 E6 0A 3F 89 CC 87 97 47
 B8 CA D1 43 33 C6 E1 DF 10 D6 B1 27 6A 43 D8 73
 27 E9 99 D0 AC F2 7F 3C 2F C8 69 44 F4 C5 74 C7
 8B 7E D5 48 BD 98 83 5A C3 F4 00 27 F3 9C DE 06
 FF 5B E0 01 8B 76 F5 5E B0 BD 55 DB 3E 60 AA E3
 BE 7B 61 C6 B7 E9 88 DF 96 57 83 58 5E 17 1D 01
 81 EC D1 80 95 25 3E 63 B2 1B 86 79 7B DF B3 4B
 A0 D1 4A 31 85 E2 C5 84 C3 AD EA 81 81 E4 60 FB
 3B F3 77 7E 30 DF E8 78 BB 53 40 70 46 E9 87 D9
 F9 0B FD 85 E8 0E C2 06 F4 18 1C EF 22 79 ED 90
 09 F8 24 24 BF 46 07 F3 3D 8A C5 AB 23 A9 17 F7
 EB 59 D3 EE FB 2C 42 1B D9 86 06 3F 48 D5 6F C5
 D6 23 87 59 8B 6E 87 6E AC BE D2 E6 03 82 E2 66
 24 F0 C7 A7 3F 06 13 7A 01 3C F3 E6 2C 3B 63 0B
 D6 D3 15 81 71 89 42 F1 6D A6 5F 08 88 7B 7C F7
 E5 45 22 B7 70 21 86 0A F0 D2 BA 64 F6 C7 BD A1
 96 B5 D4 5A 36 2B 28 63 A3 91 E0 1B 89 DE 8D CC
 B1 04 B5 4B 12 6E 49 8A B7 C0 2C 48 28 6C 89 AE
 0F 16 5E 06 A8 3C 9F 7F C2 80 0E 9E 63 1D E1 DC
 24 7E C4 D9 44 BF BB 61 47 DA AB A0 BF 12 E2 DF
 52 3B 2A E2 E2 14 A2 4C 04 00 F2 AA 82 7D 78 30
 BB 66 29 D1 5F B4 FE 0C 70 D2 BF C2 88 0C 34 07
 DD A2 6A A1 18 8E 22 A7 B1 0A A3 B3 35 39 B2 4E
 F4 75 E0 10 C5 CA F1 D6 98 AC D8 C8 74 70 8B 53
 B7 7E 27 E5 6C 3D F5 90 CA 76 2F 1B 63 0D C2 3B
 BD F2 66 99 DC 61 01 A2 D1 08 D7 77 FB 34 3E DA
 1A 5F F4 62 7A 93 2F 52 D4 02 10 EF 8B 1F 5F 59
 97 1A CD 58 EF 2D D9 78 D1 70 B7 40 E5 8A 97 7D
 F0 02 BA 14 74 98 94 4A D1 20 D2 90 34 A4 AF 56
 A1 A6 FA AF 8F 58 30 5B AF 1A 12 37 62 D3 CF 1C
 D3 6C 0A AB A0 9D 42 5F 6E 72 1E CF 2A E7 BD 6A
 22 9F 8C EA 66 94 43 2F 5A 0B 77 A0 A0 DD 96 72
 E4 9E 55 36 06 3F 25 7B 55 94 07 AF BC 1A E7 57
 8E C4 F9 EA 5F DB A2 83 AB 80 FC D1 E9 A4 A7 1F
 9E 15 24 BB 0B 67 65 A3 F5 4E 73 CC DC C5 0F 6F
 81 6B A9 10 DF 13 C5 DB F0 CF 16 8F 09 ED D9 E9
 04 61 47 38 43 57 FA FB A7 D3 76 10 21 76 2C BF
 36 71 2D 0F 09 A6 00 06 D9 63 AE BF 29 5D 44 3D
 D1 F8 56 FB 04 E3 1D 27 9E 88 65 AD 2F 6B 6D 2F
 FA 59 08 70 4D D7 56 93 F5 D2 FC E3 A1 0C B7 6D
 D7 39 1F B7 7D 51 30 0D 94 C5 E2 ED 46 E7 7B 3F
 05 6F 94 0C AA 6E 54 08 E2 EE 1C D5 EC ED EE C3
 9F FB 05 F1 93 5B 5B 0F A4 A0 8C 7D DE 3C 4F FF
 78 32 96 EE 33 BC 42 CA F1 8D A7 04 61 18 44 92
 F8 7C 56 19 BE 05 B7 96 DE 4A 34 B1 B8 53 F6 33
 78 6C 49 DA BB A7 90 10 46 A6 D1 E5 3E B8 7F 7B
 9C 99 82 16 F6 3F 44 A6 81 29 FC 03 A1 09 65 05
 24 8C B1 C0 55 BB CE 26 72 0C 9B F4 60 39 E5 71
 22 C3 99 F4 A2 EF BD 85 BF B9 C7 F9 59 79 E7 25
 5E 25 F7 BB 9D E1 4C F7 0C 14 67 C0 E5 61 AC 75
 6A FC CD A1 74 83 BB C7 09 FA FB 4F F4 73 2D 40
 4B 1C 51 A5 71 FF E4 94 0C 28 43 94 35 D2 35 D6
 DF A7 A6 63 2D 10 F8 FC B4 AC AF D7 28 E5 EE E0
 48 D6 B9 42 91 7B 3B 57 43 4C 1F 2C 45 E1 D2 48
 51 81 AE 91 EB 60 25 63 4E F6 33 65 9E C3 C1 9E
 32 05 C6 4C EF 3E 90 C1 4D B2 CD C9 A3 5B FD CE
 A3 D3 74 8D 85 A3 BC F3 E9 AC 6B E0 F5 9A 84 B4
 3B 20 2C 24 7F 04 4F 62 19 F1 DA F1 2E ED 99 FF
 0F FB 2B C9 16 21 DD 87 2C 7E A9 2F E7 06 CF 2E
 10 70 70 06 18 26 A2 73 09 87 D9 99 18 71 30 30
 4B 83 9D 4C B5 B0 91 77 26 42 FD 33 4F EC AD DC
 0B FA 3A 07 82 7D 4E 69 84 15 AF E2 22 93 8B 3A
 A9 5C 40 D9 29 F3 7D 9B 70 23 0D C8 8A C7 F3 32
 54 C5 BE 33 E7 AF 46 86 13 3C 68 96 FF 6E 95 72
 1B CB 4A B3 21 22 A7 DE E3 C1 6A 7A B2 AF B8 C5
 D5 1A 65 C1 3E 70 E6 F2 A7 D9 F3 B0 20 7D 02 09
 12 81 50 3D 5A 51 B0 7E 84 50 64 99 4C 90 0A EC
 F3 8E 2F 4E AC FB 68 DE 34 31 14 E4 1A 6C 1E 22
 66 1E 51 73 CC E2 B5 C8 90 80 80 D7 A5 FE 50 8D
 DA 3E DB 54 9C C7 D1 AD E9 0F 31 42 DA 51 43 EF
 95 C6 BD AD DA 09 AE 2E BC 4C 22 AD F0 9C 9A AB
 E1 B4 32 45 E9 61 F9 23 08 B8 B7 64 8F 8B 38 16
 70 90 C2 20 AB 56 DC CA 47 B2 37 A6 6B 30 16 37
 3F 1C BE 4E FB 29 2B B3 C3 C7 1E 37 06 A6 07 F1
 57 88 E7 EC 09 0C 51 67 F6 59 D1 64 BD 19 45 10
 2F 27 57 37 E9 A5 58 1B D6 47 E4 BD D6 14 23 13
 BA A7 A7 83 E1 F7 94 49 3A B1 A3 40 37 FD 2D 9E
 32 65 45 6D 22 0C FB 5B E2 E6 52 9A 04 2B FF C9
 64 0C D1 8B 58 53 AF 7E DF C6 92 6D 54 41 EC 9D
 32 C6 91 F7 0C 51 C2 F6 D7 22 91 C6 2B FF AD 05
 43 D0 C0 1E 39 66 06 31 EA AF F1 0D 21 1D 93 4E
 99 03 31 03 E1 01 D0 29 28 E6 35 3A 6B 0E 6A 0B
 D8 5D C5 FF 9D 8A 1A 3C 64 80 0B F3 A5 16 79 9A
 56 75 E5 44 43 AA 15 D3 65 39 30 94 BD 45 E0 7F
 5E AC B9 CF 7F 57 B3 17 67 BA AE 0D CE 3F 0D 80
 EC 95 8F 28 D8 84 84 FC ED E1 97 E8 37 8F 7F 16
 48 85 51 AD 84 FB 1C E7 73 23 6D 61 87 EF 79 E5
 4D FA 9F 25 96 AC 42 5F 33 71 E9 D5 8B 34 F1 FA
 CD DE AE 98 52 AD 1C 4D 22 29 E3 4F 29 DB 93 BC
 6A CD 4D 40 AA 1F 9D 4D A2 AA F6 FD ED E6 12 89
 10 CD CE DB C7 7E 2B A7 94 B2 78 20 E0 9F F1 6F
 6E 7F 4B 36 FC 5A 16 AD 9C 37 78 70 2F 13 E2 BE
 7D 45 BA E1 EE 60 E3 BF C6 D2 A6 A0 71 00 EF 44
 00 7D 4E 70 27 8F 36 3A F3 93 E4 73 A7 CA C7 DB
 53 F5 11 58 D2 76 A4 08 02 21 92 50 1D E7 BE AC
 4F E5 1D EC 7B DE 84 D2 F9 A0 FF 35 CD 5E 87 29
 FF DA 4D 9B 21 48 0E CA 6F D1 12 FB C4 37 C0 11
 E6 5C 03 33 EE 46 AF 77 4C B9 1B B6 F5 66 C1 2C
 5C 43 ED 7A 09 8E FD 8F ED 95 99 A0 33 6E 2D 22
 4C F7 8B 9E 57 3D 39 02 87 ED 39 0D 10 D4 E9 C7
 64 AF 65 D7 04 2C A9 85 EB CC BE 59 36 2A 2A F6
 40 CB 89 36 CB E5 AF 80 B4 B7 EB 31 57 EC 7E CD
 60 7D 5B 6B 50 04 00 91 7D E4 C3 75 01 92 05 C4
 C2 DF 0E 67 49 61 4D 54 4C A7 F3 81 2B 9F D1 EF
 8F E5 CC 5C F7 5C 3A 10 73 21 7A 7E AF 1B 1D A9
 AE 3E 6B B5 50 49 BD 23 0E E1 19 51 8B 92 57 BA
 E0 76 F9 BB EE 61 D3 EF 39 49 1B 4E 8E AE FE 75
 1A 25 83 04 99 BE 29 D1 A3 F6 05 73 2F B6 3D 32
 26 14 CC D4 3A 23 6E CB 6E BB B2 76 4E C4 F6 E6
 A5 E8 41 42 B5 67 08 F1 56 9D 56 37 CF 09 9D E6
 33 11 AE 2E 4A 52 D4 AB 47 E8 45 D9 77 D5 49 21
 BF 53 3A C8 16 CB 81 74 74 58 EB 7D 13 35 79 17
 EE E7 77 9E CF D6 AA AD 80 A4 04 1B 1E E9 7D 46
 ED B7 46 FD 48 03 EA B2 91 80 49 6B C7 F8 C8 0B
 2F 8A 90 FD 93 DF 4A C7 4D 19 B8 0B C9 C8 0B 37
 1F 5E 1F 89 A2 5F F6 CB 37 2C A7 7A 5E AD E3 51
 F1 3C 21 6D 30 3C F9 8B 12 45 FA C1 17 7C 7E F0
 B9 58 0A 6F DE 3E AF 8A 0C F7 66 D5 F3 5B 0F BA
 B5 79 77 2C 41 67 D0 2F 01 D5 53 AE 26 40 73 E9
 9F D0 FC 7A 51 3D 95 09 48 62 3E 94 51 63 AC 06
 DB 99 72 F3 DF 28 45 2B 05 71 71 D3 BA CC FA A2
 69 7D 07 56 B9 9C 3C F4 73 A4 80 A0 1B 46 2A 25
 F1 0A 1A D4 CB 2F D2 0A DC C7 90 0E 59 00 B6 79
 5F A5 A3 39 12 EC 0F D6 F7 4E 7E 56 DE 9F 9A 5C
 E0 38 9C 01 99 71 DA 52 F1 4C 74 A1 D9 63 5B E6
 EA 86 E2 4B F3 51 88 F0 39 67 4B 37 B3 36 98 4E
 FC F5 D5 13 06 E9 0E 41 46 D2 7B 88 62 9C 54 30
 76 14 CD BA C3 94 F3 D6 26 B7 90 00 61 76 EA C9
 18 65 17 A8 A2 4D A3 8A 0C 0A 34 29 48 58 31 42
 BA 5A 30 75 8E 7C F2 6F 68 8A 6F 20 2E 8B 39 F7
 9F CB C0 E0 35 FD 64 FF A6 30 B8 36 45 3E 37 07
 43 F3 9E 53 2D 32 61 E0 1F C9 FC 6C 9C D3 21 02
 45 57 8F 7B 9C 4A 75 43 26 D3 4B 51 AA C6 8A 55
 9B B1 EB 10 76 2A ED 0A 3E EF 82 21 C1 E7 82 B7
 6E E3 CF FA 4E 1D CC C0 68 2C 8F B0 1E B8 28 B8
 1F 13 C5 8E FE 3F EB 2B 8B 61 CA 2D C2 D9 A3 FC
 2B A7 9A 26 03 52 5A 9C 02 BC C3 42 C8 B5 A8 33
 C0 BE 53 59 97 B8 A6 FE 1E 15 15 9E 01 32 A7 2F
 6A 91 8B 26 FF 11 31 47 70 3E 72 46 60 D0 C1 43
 01 5B 26 69 DE 4C 4E 8C 16 55 4B 6E 65 0D 0D C1
 75 34 F0 86 F4 DC B2 04 EF 64 15 3E FE 61 D2 CD
 E2 14 5A 8C 5D 43 3A 91 1D 0B E4 42 48 76 30 CB
 A5 A9 0F DB 2A CB BC 1F 67 3A EF 12 CA C4 77 40
 67 B8 63 F8 80 55 4D CF 95 69 EA D0 55 1B 52 8E
 C3 C3 FD 30 17 43 8D E9 AA E7 DC DB B2 3F E7 7D
 72 2E 76 BD DA FD 07 14 03 B6 D7 3E 19 B7 16 61
 35 45 2E 83 C8 C2 16 BE 2C 9D ED 62 77 D4 E0 4D
 B6 98 F5 C0 9F E2 23 A2 8E D9 0E B2 9C 6A 90 D8
 EC 3D E3 5E 12 7F 36 F1 1A 5C BE 74 D5 43 C9 CD
 04 C8 77 3B D7 1F D7 73 18 EC 6A 8F FE 41 39 21
 B2 5A D9 16 67 15 A1 75 D3 53 A5 85 C6 B1 1D 80
 C7 B9 F1 68 7C BB 71 F7 1C 26 64 1D 13 CC 41 BF
 CF 9F 0B A5 65 85 1A 44 3F 2E C7 00 36 93 B2 EA
 27 52 67 A1 FB 7F 24 29 5C 2D 81 87 87 9B D0 B3
 5C 30 CE A8 84 98 A8 D3 AE CB 06 AD EC 90 03 22
 C9 B0 6A EC FF 76 78 49 63 26 FF 34 3B 49 7C D7
 85 38 E4 CE AA ED C0 78 27 7D 14 1B A0 AC BB 10
 0C 36 1D DB 96 69 C1 11 D8 B2 B2 95 73 34 F5 C3
 E8 3F CE 9F 51 62 84 76 A3 50 49 16 F3 F1 36 B6
 1D 38 BA 5D 20 B9 96 CA C2 B8 C3 E1 9E 0C 0E 4C
 E3 DD 25 06 95 E3 7E 46 D6 E3 19 D6 B9 7A CF F8
 8A 39 7E 10 A1 72 50 4E B5 5A 9D 54 45 CE 22 C6
 E4 AF 09 C7 E7 D5 DA 3B 85 F6 CD A0 DD 7E 35 C0
 94 6D 9A 89 9D AF 9F B4 EC 07 58 28 CA 2D CF 1F
 EE 43 A4 68 A5 ED 19 F3 0B FD 56 36 62 24 DD 99
 CB 41 84 CA 85 A9 53 D3 48 EF E3 66 59 71 35 FF
 48 92 B3 82 0D 16 55 40 55 DB 09 2F FD 5E 00 8C
 90 97 C5 F5 BA 6C 45 06 89 15 75 DC 2D 88 2E 77
 5C 1A 02 4D 44 F7 8E 02 2F F4 08 B9 0C 27 0F A6
 86 01 FF 90 60 09 BA B6 82 5B 56 81 0C 48 FC 6F
 D1 0A 07 46 5C 45 04 35 3C DF E4 4C EE 03 76 23
 A6 77 18 FA FA FA 16 7E D6 9B F5 3E BD 33 6E 49
 42 4A 48 6E A7 55 44 82 20 0B F8 6D 47 90 40 3D
 B0 45 45 6D 05 70 89 07 42 CB 04 13 36 C4 47 B3
 2C 3B 62 90 7B 61 DA F7 DE BA 7C C4 70 42 C2 EB
 A1 D8 9C A8 0C 41 26 25 69 72 01 4B D9 8B 21 C6
 94 66 66 6C 52 0F 51 DF A2 DF 10 93 A0 5E 54 BF
 7D 17 B5 DB 98 C4 FA 7B 46 EE 7C 05 CF BD E4 BE
 B2 AA 04 6E A1 35 7F 70 88 65 CD B7 86 1B 61 03
 92 FD AD 45 BE D4 4C 5B 3D 80 CB 10 A6 B5 AF 86
 6E B0 17 AC 7D 2B 77 51 B1 E7 54 61 CF 93 15 D6
 F9 60 29 5C 59 97 8B DB 6F 5E 87 72 47 82 63 BC
 63 93 D1 E3 10 46 78 FE 95 04 8F CE CF BD 48 A2
 33 FE BA ED 56 75 47 A7 DF 13 91 8C F4 40 B1 8F
 A0 49 A3 F5 3A EB CB AD 12 77 3F 19 C1 13 DA CE
 F3 BC 72 45 0E 86 5D 31 29 09 00 D4 D7 EB F9 2B
 A5 6D D1 C2 01 3F 89 1E 54 58 F8 7D 48 87 8A D4
 42 D8 DD C0 8E 5B 11 4B 48 15 AB FB D1 59 98 DD
 60 6E 49 45 96 EA F1 15 E0 8C 5C C8 BF 0A 27 E1
 BD 23 94 1E 1F 0A 2B C2 29 29 2D 1C B9 57 0C 09
 21 4A FC 01 05 DB 30 78 A0 94 2C 63 4F 6F 4A F0
 91 B5 F8 EA 93 49 ED D2 ED 2D DB C7 8A 30 98 0A
 A0 5B F5 CD 35 54 E4 62 7F 8E BE BC 45 33 F4 23
 ED 49 98 AC 88 CC BA 0C F6 60 2D 18 46 65 7C BF
 E2 84 C4 20 FA C8 D3 F2 71 65 04 60 C6 1D 78 09
 9F 40 F2 47 84 2F 11 A4 09 9E BC ED E7 17 E6 42
 95 83 D2 69 00 C0 A5 F1 08 E5 2E 7D A5 7C F2 51
 FF EB 13 83 ED 70 1A 97 8A 79 D5 2B 9B 6C A3 EE
 28 80 6E B1 88 EF 31 EA 51 48 AE 8E DB BE DD 1F
 51 C9 13 45 85 3B F1 7B 36 37 FC 64 90 50 A8 C9
 A8 76 39 84 63 AA 48 95 00 20 A5 F9 9A DB 2D 7F
 F0 06 18 FA 47 DE 5A 02 0B CA 49 BD 0E 7F 07 0B
 D6 E3 F0 A2 34 EC 80 1E 8D 30 1A 63 D1 34 73 94
 36 A4 B4 16 04 1F 1F EE A9 73 03 12 0F E1 21 F4
 5C 97 1F 24 A9 8E 25 8C 18 A5 90 58 B8 70 59 58
 5A C2 A1 C4 98 43 8A D8 B8 7B 1A B7 DF FE 48 0D
 6A 83 05 E5 88 F3 90 C4 22 CF E7 C8 B7 6F E9 AD
 DA 7E 31 08 48 58 99 55 E6 FD 6C A6 8E FB B0 DC
 68 D3 5D C0 55 18 72 FE D0 8E 21 A9 26 4A 12 AE
 F5 3B 18 16 C3 68 AC C8 BC 7A 2B 25 72 3B A6 27
 12 07 04 23 29 F0 22 1C C7 BC 30 CD 09 79 34 8E
 A0 CC A6 73 03 0F 01 96 3B 3D 81 B6 21 DF 06 0E
 6C 99 34 28 10 4E 3F BC C4 31 81 08 92 59 DD 4E
 88 28 C3 D4 AB 13 D7 42 03 50 BD 70 01 AC DB 20
 6D 70 DD F4 AD 97 3A D5 11 56 11 F6 77 C5 0B D9
 84 AC 96 B2 23 1F 96 0A 6F A1 70 F8 1C D3 59 8E
 C0 B8 4F C0 BB 8D FA B5 CF 95 DC E7 41 CB 21 28
 AE 2E 64 90 D4 9F C4 FE D2 88 04 5D 20 43 DD E3
 EC 40 CC EE 92 4B E2 F2 03 74 AB 29 0D DC 1F 45
 74 EF 90 EC 45 E7 90 0A F5 58 D1 F6 7B 74 1F F5
 69 73 AB AB 40 90 C5 BE 0F 97 58 83 C3 3A C9 FB
 04 CA 71 F1 C0 A5 6F 8C 5F 2A A0 84 ED 47 8D 2B
 A9 E0 AF AC 4C DF 77 26 B5 30 2C 00 BC 6E 7A 94
 22 DE 40 AD E0 60 32 E8 42 4C EB 1D FB C0 3F 96
 A7 50 41 57 9E 83 88 D1 A8 F1 24 FC 24 7C D7 5A
 FF 7F 0D 1D 1F 15 F2 23 35 58 2F AC 50 0C C2 3F
 FA 92 F7 EF 35 AB 25 18 35 0E 49 81 4E 00 2A 1F
 3E 6C A5 18 DC 9D C5 1F 77 DA 6B D4 4B 03 C1 AB
 24 BA 8C E3 2C 6E 58 6E 23 C7 FB 93 2C 67 F9 3B
 A7 8C 5E 74 CC D6 A3 1A 76 75 D7 F6 06 5A 25 83
 88 4D 6C 36 A1 FD 20 78 9A E8 3B AE A3 D3 71 1B
 6D 4F EE 28 BF 88 9B A3 F0 3C 19 83 27 A5 71 CB
 26 04 C4 F6 A3 C1 CC 6D 6B 54 3D D6 2C E4 FB A6
 BC A3 30 60 41 E8 54 BC 43 78 42 AB 18 BD 10 49
 3B AA D8 49 9D ED B8 27 4A 02 CA B1 5D 32 B9 CD
 D5 9D F0 D1 51 BB F7 8E FC 1A 5A C0 97 96 B9 CA
 E9 EA 4F 2E AE FF 51 AE 98 DC 00 C2 9E A5 7D 8E
 B7 78 8E 09 E8 66 C2 E6 61 81 6D 9A 53 AF 25 E2
 29 F5 83 B8 7B 35 1D 35 F7 B1 B7 36 75 8C 6B 4B
 66 33 89 AF 56 3A 39 D2 D3 00 2C 8E BE C7 1F A4
 A4 D5 92 AE 10 52 CE 6F F0 A6 C0 E9 75 D6 AB 66
 ED 58 6A 0B D3 A9 B0 9B 60 2C 09 B4 89 D0 6E 4E
 CC 0C 8B 2E 3A 47 91 DB 08 69 08 4A 87 CB 8A 70
 DC A2 12 DA CE 39 92 7F B5 F5 5D 52 29 83 62 E9
 6D D4 98 C1 B6 62 7D B0 DB 48 20 5C 98 2C 0A 99
 E3 F2 48 FE 66 F8 29 13 49 90 A4 AE 7A 1C FE 57
 28 32 13 89 1B B5 45 08 A6 35 CC 4B 60 83 A5 9C
 9C 16 E7 1E 8E AB 23 73 2E B7 84 0A D9 FF 76 94
 A8 68 DB C6 4C C9 9F B6 55 76 0E 3D BF 29 43 E1
 EF F2 75 81 42 13 61 01 35 8C F6 C7 2F 2F BA 6A
 9B 9E D0 0D 53 28 FD 99 62 8F 7C 13 24 DB 4A 74
 55 EE 19 FB 10 81 C6 E7 64 53 9A CD FA 6D 9B ED
 43 B5 A0 5B A9 EF F2 BF 7B 53 C0 FB 2A 27 4C 4C
 CC DF CF 8B 1E 51 B3 E2 66 22 EB 59 D6 B8 6D 20
 A7 67 C8 05 8F 4A 2D 25 79 92 FF 07 BB 00 02 EB
 4B 84 4F 11 2E A4 36 74 21 11 31 58 0C 93 2F 98
 BD 6A A4 A8 F7 8C F0 23 EA 15 33 5A 7D F3 67 BF
 93 96 45 A6 49 69 5B 76 5A 1F A9 53 A9 1B F5 70
 85 17 0C F1 AC E9 55 04 E2 70 FD DD 15 32 96 9C
 84 7D EF A3 FB EF 6C 7B A0 C1 18 9D 85 68 87 60
 00 FA 63 34 F4 D6 04 37 1A 22 00 DE CF F4 A3 FF
 CC EC 08 97 0E 08 5A 2C 7F A6 57 B8 D2 73 F2 F0
 52 FD 09 8F DD F0 D3 DE 12 3F 85 71 02 E2 1E 3F
 1B 20 2D 76 6B D8 F1 5C F9 2B 90 D1 23 6A 18 9F
 97 A6 23 B7 9E B9 04 C3 96 32 05 5D 44 7E B0 89
 E6 69 F5 A6 99 0B 58 54 4F FA 6B 07 C0 F1 FB CB
 D0 A3 DC 1E 3A 3A 28 C8 72 8B 2B 7E FC 50 19 2A
 7A D3 C5 91 03 65 83 24 7D 85 27 BE B1 2E 6A C0
 0B E7 A3 32 8F E1 2A 49 06 CF 14 53 F4 45 98 9A
 5C A5 34 4B 11 99 EC E6 0C D0 3C 5F A0 6F B8 79
 0F 28 81 63 38 82 FB 6D 9C 22 C6 3A 67 65 9D 17
 90 42 B0 98 D8 66 70 EB BE EC 52 D4 B3 D8 8A E3
 92 2D A4 25 3D C3 EB C8 5A 71 97 41 69 F6 37 5B
 78 75 C1 0D D9 A9 F9 1F C2 BE 3A 39 1B E1 D2 3F
 43 DA 42 55 EE CA 9C 1F BF E8 38 03 AF AB 4C 53
 63 4C 02 89 36 18 31 C9 C4 6A E7 F2 CD 65 9C 1F
 5A 2B 6F 84 71 EF 22 2F F6 04 19 B8 F7 C0 D1 7F
 51 CA CD 0B C7 F2 1B 74 7A CE 3F E0 A2 69 59 92
 60 A7 D4 6D 08 75 46 E7 9E 47 77 5D 60 A3 0A 97
 F0 E6 FF 12 AC 47 2A 68 05 2E 81 F4 46 73 0B D8
 4D 7C ED D1 38 CA 25 FC 22 B9 E2 FD 48 F6 21 B5
 7F F1 D3 76 B9 29 C9 24 86 D8 5B 76 DC 2A 16 69
 45 B6 41 1B 54 09 DB CD DA 5D C2 CD B3 8F 26 06
 39 5A C0 1C E1 80 35 22 91 FD AE 1F 8B 2A B6 7D
 76 DF C9 8C F3 C8 F2 DE BE A8 4B 3C DC 22 A2 61
 55 44 05 DA B2 CE AE 49 35 E3 FF E5 9D F4 E9 3C
 FF 9D D7 0B 8A B6 91 76 C0 35 3F D9 18 F8 8C 8E
 7A 0F 4B A3 A3 EC C8 37 C8 4E 95 A8 37 EA DC 45
 DA AC 46 98 F3 33 84 F6 4F 03 21 9C F4 54 E5 67
 46 B7 3E 3E 42 22 91 16 B3 2D A9 B2 AC 1D F4 0B
 C1 8D 34 66 56 AE 46 74 91 47 8F 90 1F 59 39 DB
 A6 00 53 2D 91 9D 30 16 A0 54 30 A3 6F 68 7A B1
 C0 6A F4 95 DA EC BB 17 5D 8E 03 2C 6A 11 99 C2
 68 CE C0 46 91 7D 59 64 7F 17 74 FC B3 3C E9 83
 EE 79 EB E6 55 22 87 C1 A0 40 27 CA F5 EA C5 42
 DF 04 24 7A 14 2A A9 27 64 68 96 A5 9A 5E 1A BD
 FF 5E 56 FC CF 18 01 45 71 0B A5 AD 81 85 5A 1D
 AD 0E 56 D0 8C 90 3B C9 84 1E 04 B5 9A E5 0C 6E
 99 E3 F7 47 D0 04 2D 36 DD B1 F6 A6 80 04 75 33
 E6 DC D8 7A D8 B1 49 41 8A 46 D4 57 9F 1D AC 52
 F2 B7 7D 73 FF 1B C8 37 08 DC 65 D3 2D 75 4C 47
 3B FD 56 A9 D3 CC 89 72 09 50 06 F0 11 BD 31 A8
 4C 17 93 17 F5 54 1B 76 60 DE 94 D4 16 54 EC BC
 D4 0D 18 51 5F 5E A4 8A 09 6F 90 8C CC AD 1D 19
 64 8B 7C 90 5C 10 14 37 BA 7C 67 13 C1 81 74 FC
 CE 7C 4D B6 86 63 FC 2A 88 B5 04 DA AE AF 74 0D
 14 77 A2 76 D6 50 AF 81 52 65 C4 79 49 AE 82 A1
 92 1F 3F 43 EE F0 42 25 B6 A4 A2 A6 ED DA BD F0
 E0 27 BA BF 92 53 CC 9D D9 B7 0A E6 7A 8F 65 D1
 BD 19 4B 47 67 88 F0 D9 A3 58 D5 92 6D A1 1A C2
 75 22 3C 9F 96 BC 92 ED F7 A9 BB C6 D0 1E D2 27
 41 28 4C 9A 02 BD C5 1D 4A 08 22 BB 6C 4C 8D 32
 03 3B 84 C5 47 73 4F 15 E2 49 E1 A7 7F 0D FF 02
 D7 04 41 D9 1E 0C BA 03 AB 91 B4 7D DC 41 4C EE
 59 C7 A9 3E 5D CA 8A 10 13 74 82 EA AF 5D 15 0B
 6C 66 95 48 73 CE D1 82 0D 12 D3 89 72 01 80 2E
 4F 12 96 D7 D9 6F 31 C0 54 BD 37 AB 78 4D 2A 53
 13 01 8C B5 0D AF 6F 80 AF BA AA 6C E2 11 AA 39
 C5 9F 30 C7 61 BC 9D E6 91 22 EF BE B0 C1 30 2B
 0C F0 37 61 3B 79 33 F0 05 7F 38 9B CE 3F 32 63
 3B F1 2D 0A 62 A2 57 66 90 4C CF 39 46 AE 6F 65
 2B 45 A3 B1 FD 82 33 D4 43 C3 2C DC B2 56 98 1F
 1A 73 E4 24 23 74 AE 42 6D B2 A6 D7 9C A8 F2 99
 EC DD AF EF 60 55 E1 0B C3 63 04 4C ED 0E 66 0D
 A2 9F 17 C8 26 0F 70 83 E3 FD D8 95 86 44 3E 3D
 39 23 9D F2 61 2E AF 8C A7 14 B4 83 2C B5 9C A6
 39 15 54 30 18 94 16 86 A6 39 89 5B 16 6F 5D A1
 EF 86 FD 4C 0C 54 C9 FC 59 30 5C 06 BB 94 C0 6E
 13 A3 56 A7 E0 1C 91 AB 48 8E BF FA 7D 44 6B 91
 23 D0 E2 42 F9 ED B5 A0 37 C9 B0 7E A3 88 F7 65
 A2 72 3A B4 80 01 1A 23 53 54 B5 DB CF F1 33 8F
 D4 15 FA 44 52 13 C5 85 C6 50 3B DD 7C 34 A8 68
 7B F0 BF 83 58 F7 1F 40 EC 2A 74 75 A2 1F FE A7
 2A 61 2F 18 5D 9A 89 6C 88 09 D0 8C 15 F1 17 62
 17 79 0F B1 DC 17 89 29 83 95 0B ED AA 59 F6 DF
 6E 58 68 4C 19 70 03 F2 0B BE D7 AC 2F 7A 63 60
 A0 9F 0B 11 09 30 CB 2B C5 8D 2B 07 DC 92 9A F2
 49 CF 40 6C B3 B2 5D FD C3 51 45 82 73 96 F1 6E
 AE 34 7E 6F 9E AB 13 93 62 13 AD 39 E2 80 5A 9F
 AD 1E B8 85 E6 34 38 4F 60 B7 A8 9A E0 B5 00 A1
 A1 82 FF A8 72 DE CF 19 23 C7 D0 68 ED 75 1A 13
 29 C9 9A F4 5F F8 E2 69 28 CC A7 5D 7E 38 C1 81
 27 43 1E DE 5E 2A 28 4C 35 81 AD F0 D2 E8 CD F6
 62 48 72 62 51 19 40 AC A4 F7 A2 CC B9 05 91 C8
 23 E9 3F DC D6 85 A6 F1 CF DA 6C 86 89 9B E1 68
 1E EE 92 0E D0 90 65 61 47 58 8D 92 07 89 CC 4A
 03 84 AD BA CE BC FD A1 5C CE 90 DF B1 CF 11 25
 81 02 2E 5C CE 32 B6 72 27 60 47 64 5E 99 A7 72
 41 6E 7B 64 56 04 D1 98 93 27 D4 C2 E7 55 54 BD
 5E 84 EE CA 4B 8E 65 F4 70 98 92 73 1F 74 BF 8A
 1B 76 19 42 C7 A2 8F 42 A2 4F F0 6D 94 AB D0 C1
 3A FE 50 8C C2 71 B7 C2 F2 8B 72 22 03 D7 A9 B0
 82 D3 08 60 5C 0F A9 C2 DA 61 C5 4A 79 51 71 C4
 F1 DC 5B B7 78 F0 FA 3C 51 E9 27 CD EA D2 CC DA
 DD 52 0A 2D 56 65 1E 7C EC 1F B8 DA AE DB 15 3D
 B8 19 50 DF 0E 21 99 95 FC 29 AD 5A 37 07 F4 D1
 5F 79 35 53 FC 61 0E 26 9D 23 44 07 ED 47 75 E8
 37 7D 26 A5 2E F1 A6 01 DB D4 DA 60 73 86 4C 7E
 32 0A 52 7A DE 70 BC 97 12 17 05 B7 DB C8 E5 A0
 16 8C FA 73 FB C7 24 91 17 CC 8A C8 3D 36 8D 67
 B1 83 EA BE 76 D5 2F A2 1C 13 9F F4 2A CB 54 11
 EB D8 67 08 36 5D 4F EF 83 DD EF 70 29 D2 95 78
 C6 5B E5 C6 38 43 F3 AD A2 B7 EC 24 83 A4 01 13
 30 74 06 8A 78 A3 EA 21 62 2F 30 DD 4C 25 CF B9
 E4 9E 29 25 C3 70 CF 38 3A C5 BD 59 B8 98 15 02
 F7 64 E0 8E 32 BF BA B3 5F 19 D4 D8 DE D9 C6 52
 96 60 BB 0A 1F 8D 01 F3 5C 81 14 CA 1B 20 43 C1
 1D BC 66 8C 5F 7D 7C 5D D0 65 A0 DD EB 0D 35 09
 CB 17 49 44 E7 A2 B8 34 E7 1F 17 DC C2 6A 2C E0
 A5 6B 28 D0 E1 4D 39 DD 98 CB F8 5F B1 6A EA A2
 45 B6 FF 93 64 7A 71 EE 23 EE BD C4 CD C1 61 F2
 82 50 7D B0 7B FD 8D 41 D0 DB CC 71 8C 67 67 7A
 7F F6 EF 02 A5 DC DF 4F DD A4 C2 DB AA 15 25 7E
 F3 5F 41 8B 01 9E 1E DA DD 72 83 AD A1 72 25 00
 BF 25 F6 0A F9 C3 5A D7 EF 40 5B 66 A5 67 FA 1C
 DF A2 52 3F E5 D6 3E CA 4D 29 66 07 D4 D5 D6 4E
 61 2A A2 CB A6 97 84 35 A1 12 BD 1F 4B 71 9C 9B
 2A 44 07 3E 45 26 DC AC ED 43 02 02 0C 0D 64 D1
 DB CD 9D AB 11 17 56 48 FF 56 D9 AD FA 38 12 3A
 57 EA 05 B5 6F A0 73 E1 AD D6 D4 56 36 A1 20 08
 21 D6 53 F5 EF 0F 29 E1 18 EA 87 BB F3 FA DE E8
 33 7A 45 2B 2A C0 1B 66 EF 31 F4 0F C7 62 C0 87
 EF D6 FD D9 8D 43 3D 2A F3 74 39 94 AE 52 94 1F
 58 28 01 CD D1 B8 D8 D3 D5 CC 7A 09 40 CA 74 35
 50 C7 C3 AA 08 33 06 69 4E 52 8B E6 81 09 65 EF
 DC 1E F0 7A 83 EB 9D B9 4D C8 0E 79 63 4F 1E 96
 15 88 CE AF BD AB 27 5B 9A BE 41 8D 02 93 F1 1A
 9B 1E A2 84 03 D6 05 AC 0B 62 F1 BA B1 E0 78 6F
 EA 63 2C 29 89 4A 4C 8B 56 2B 29 29 86 54 B7 61
 B1 BA 8E EE 6D E5 F3 32 6A C4 9D BE AE C2 E9 9F
 CC 5E 25 D5 B2 10 D2 F7 0E 2D 13 FA 6A BA B7 A4
 6C 3D BA 0C C9 24 73 D1 25 50 DE C7 82 C9 7D 1E
 D1 80 9D EB 1C D3 CC 5D 09 56 76 97 D5 38 F6 7F
 A4 16 3E 38 CE C1 16 38 17 90 1E 97 DB 67 92 9E
 E6 60 A1 60 99 ED 52 59 39 16 4B D7 41 18 11 20
 F2 31 FF D0 DD EF FF 15 21 C5 EB 7D 76 D2 70 C3
 B4 B5 36 CD 2F F4 9F F8 AD D8 AB D9 BD 1A 39 B9
 2B F3 A7 2E 07 6C EF 01 B7 8F 6E 2A D7 FD 88 3A
 55 5E 99 ED 2D 3B E3 CB DF EA FD 46 69 01 D0 C6
 3D 5A 8C B2 C9 C5 8F 1F B9 0B 99 5B 45 63 A3 DA
 E0 FF DB 93 EF CD 0C E9 55 C8 C9 51 1D F8 2D 6A
 F7 75 51 D9 5C 32 53 B8 27 D1 96 83 0B 3A 20 DD
 DE CD 3C DF 6D 77 06 75 0A 70 D6 46 77 D7 C7 5B
 18 B6 34 BE ED 7B 40 98 67 F9 04 E1 89 61 BD CD
 F9 2F 9F 5E BD E8 EB C8 0B DD 00 FD 97 63 A8 FE
 C8 D3 51 08 2D 95 63 85 F2 E2 16 01 35 80 D8 31
 02 76 C8 62 A2 2B 5D 3A 13 D9 4C E7 58 93 16 80
 05 32 43 FF F1 1B B5 5B E2 47 83 5D DE E6 FE 87
 1C 6F BD 56 89 ED 48 F0 44 9F 6D 0F EE CE BD CF
 D8 CC 55 18 8C 18 87 F3 C5 45 9B A9 62 64 21 51
 74 BA 7D 67 00 06 3B 2B 9B 92 DC A2 B3 B7 D1 15
 DB BC 8A 17 25 89 75 B1 88 C4 B0 42 CD AE B8 01
 47 4B E4 DD 18 DE 6B A1 5B 1C D2 10 E3 81 B5 89
 D1 33 95 38 69 23 DD D5 6C 6A 2C 8E 95 43 A3 41
 E0 DC 73 88 CB C9 D1 94 87 CD 3D 0B B3 8D 5F EE
 C3 73 05 BC A8 3E EE 74 D6 0B C6 C0 90 93 C8 A4
 55 53 33 16 73 38 53 9E B0 E4 EE 88 96 76 94 4F
 4B DC 5C 60 E3 A0 43 8C E2 92 E1 1B B4 76 84 18
 06 E0 38 B2 C1 6B 43 DC CD 04 59 FD 5B 38 6D 91
 00 76 43 FD 38 B3 00 6F 62 69 DF 5B 54 32 93 7D
 F0 DC 9B 94 5F 02 9A A7 2E 7A 39 B0 CD 80 BD 6D
 79 06 AE E9 7F 37 E3 C8 02 35 07 04 29 22 8A 58
 0A DF 6E 72 31 5E FE 82 36 81 7E F1 69 47 A5 00
 F5 D5 79 A6 89 FD 34 76 02 97 0A 9B F3 E9 D7 2E
 4C 1A CC 44 9C 57 A9 87 66 E2 59 7C E0 36 DE 0E
 4B CD C3 09 63 D7 26 D5 51 DA 0A 06 EF 14 04 56
 7E 41 19 08 7D 34 D5 17 BC 2A 6C D9 C5 0C B2 CE
 D9 AC C8 1B 3F 43 CB 10 AB 2D BF 20 7E 0B 09 21
 84 9A FC 18 1D F8 95 67 C5 97 52 32 FD 5F E6 5D
 94 01 1E 36 BC CC 75 8B 0B CE E9 00 CD 60 18 63
 DF A6 2B 14 EB 14 99 C0 19 66 93 D5 4E 12 0E D1
 EC D2 15 C3 ED 66 4F D1 D0 F5 B7 C5 ED A7 B8 5A
 79 33 ED EF 81 31 97 FB AC 66 CA 01 F4 7F 01 5B
 70 12 BD 0F 10 E8 77 A3 91 13 A9 58 0C 8A 7B 0C
 1F E9 FF 70 DD 8B FE 9F 32 98 69 8A 03 89 13 96
 6F 1A 4C 1D 45 76 97 EF 50 C0 1B 4B 8F D6 B9 BE
 1D 02 BC 7D 03 C0 18 E7 58 33 EE 03 DD AB 1B D3
 4B DA 45 CE BC 18 B6 12 9C CC DC 7D 7B 58 44 46
 2C 27 00 E8 68 71 25 B1 53 6E B5 75 97 FD 43 29
 33 04 CC 54 66 D5 76 28 54 4E 55 82 69 82 2D EA
 5D 28 BB 4A 9D 2F C0 99 FF 89 D8 F4 B1 7C 00 6E
 E2 46 19 F6 48 0E 31 A0 25 6D F0 D7 0F 24 85 49
 92 A7 65 60 FA 37 59 DA 36 57 CB 2E 14 66 E7 0F
 81 D3 F9 86 4B D4 E6 C6 27 06 2D DC B6 86 D3 2E
 A3 3D 1C BC 89 16 C8 BA 85 52 B4 C7 EF 2D B0 54
 59 51 99 B7 7A 2C 1A 48 CF 9A A3 DF DB 03 7A 10
 ED EC 70 C8 0B EE B9 7F 35 8D 4A E3 04 49 BD 71
 D6 90 3D C9 64 EE 6C 67 03 8C 31 D8 22 30 B6 54
 B4 38 E2 C7 88 63 04 CC 90 96 1C BF 30 A7 12 89
 F9 65 2E 72 17 D3 8B DD 28 40 DA 15 C0 AE B9 68
 49 35 56 D6 C3 B6 DB 7F 1B 81 89 0F 4D 80 CE D8
 11 FC 99 2B EA C6 8C 7D AA 05 4F 1C 2A A8 13 7A
 09 DF CD 13 8D 57 E3 34 7E 8E 4F 59 DD A9 2E E5
 F6 4D 4C A5 41 3E 1C B9 44 28 8E 38 C4 4F 47 97
 93 1F 90 93 30 46 E7 FB BB 3F C3 F7 51 50 68 17
 8F 58 34 75 3E 21 61 3F 60 4E E4 24 96 13 84 34
 4C A6 29 58 CE 15 8A B4 0C E5 A7 C3 1E 45 F5 60
 F4 C0 88 03 13 DD 57 0D F9 E6 D6 4B 0E D5 F3 2D
 41 5B 05 F1 78 A9 56 74 40 23 52 2A B1 46 EA 98
 09 F1 6B 1B 58 8C D5 15 09 AA 50 AD 51 EE 2D 84
 CA 18 20 9D 3F 01 04 AC BA F4 B3 C8 8B FA A2 77
 ED 41 4D B3 9C 89 70 AF 2C E8 CB A2 F1 87 E2 A2
 D9 09 D0 B5 5A 3C 75 57 07 A2 66 B7 3F 48 45 56
 59 12 C7 76 23 27 41 48 DB A9 5C 5C D1 A6 54 F9
 6E 53 3A E7 03 69 88 38 A4 7A D0 01 64 0E 6C 3F
 65 FF B1 06 24 B4 37 98 30 AA 6A 58 7F F6 B3 E2
 99 A0 ED A1 C7 84 4A 37 1F 9F 9A FC 28 F7 7F 77
 EE 14 D0 F7 4A A4 56 FF 0F D8 25 17 01 D9 02 38
 B5 78 99 7B 48 99 34 AA A7 1A 72 02 51 FC CC AB
 61 EC 3D 37 F8 5D 70 96 E7 60 3B BB A6 2C 07 56
 CC 65 3E 3A 8F 78 A5 90 FE EF 20 6D 60 37 7D 77
 42 17 BF 66 E2 36 D6 C0 F3 55 E3 FC 41 47 52 A6
 7C BD 45 7D 16 1D BB F1 79 58 28 45 B0 EA AB 77
 A9 9E 6E 23 A9 0D 3B 30 F9 FB 51 15 10 0C 29 A2
 FB 92 08 3F 6C 04 B3 3D 0C 19 5B 84 49 70 A3 27
 E4 E3 CD B9 C9 3F 1A 70 72 B6 A6 69 EB CE 3C 27
 A8 BF 34 AD 05 43 5B FD 8A 25 E8 54 27 48 73 FF
 24 90 35 2E DB 15 F3 A7 0B 06 6F C0 B7 D9 94 75
 F8 3D 45 53 3F B9 37 F9 15 9D ED 79 7A FA 84 6F
 B7 1B AA D6 15 F8 50 6A 9F 7C 11 FA C6 ED 81 8E
 FC DE 19 2A EA F1 49 AE 4B A6 2D 45 47 30 28 F4
 FD E2 2A 33 E5 E5 D0 2F 96 BF 33 27 04 E9 8F EB
 39 8B BB C2 83 C7 2A 4D E2 02 07 8D CB 13 DC 9E
 9D 8E 4E 1F 94 DC 1A F6 FC 91 90 58 D4 9C FE 76
 9C 84 E4 EA D9 9D AE BA D9 13 8D 54 E1 D7 D4 E3
 E8 E6 E0 B6 C4 27 E8 E5 9C 9B F0 99 63 4F 9D C8
 97 F6 AE 2C 0D 4C 29 EB 96 16 CD E1 E0 D8 CD 94
 19 FE 92 94 43 5A C5 ED F6 61 1C F4 A3 40 05 E8
 E3 D4 B1 4A E1 AF 21 2A 97 6A 99 FE 3B 91 5F 5C
 A4 AA 1F D9 58 26 7E 30 32 3C 3E 51 85 62 47 00
 A8 0F 5A DA 63 8D B4 6E C9 D3 1A 14 F7 86 B0 09
 96 97 B7 82 EF D5 D5 E1 68 92 59 AB A3 F7 1B 92
 79 61 65 FB 15 5D B3 7A 75 69 1D F8 B6 B6 86 86
 89 97 F6 8E D5 92 F7 F0 9D 31 0C F8 AA F5 15 F7
 DA B8 FD CE 7D 6D 63 07 60 F4 E8 8E AD 43 BE 67
 72 CA E1 83 B6 82 8A FA ED BC 92 D2 30 83 0E EA
 DA 09 A3 0A 4D 3A 88 95 DB EA 7A C1 97 0A BE A6
 41 5F 2A 75 1A 6F 10 6E 7D D3 E2 0F E2 68 43 DD
 7C E4 3B 36 F7 03 E3 A8 80 01 50 B2 DC 2B A4 71
 FA 96 A6 B0 8A 9A 90 04 0A 65 C5 A1 D6 73 4A 6D
 EA 67 07 0C 0F 04 AB 25 9E C5 04 71 F3 B6 6C 0F
 22 42 C8 59 8B 82 CA 58 B0 5C F2 0D 61 EF 19 D9
 88 4E 6C 3E 63 47 F0 F3 2E 29 9B 56 11 C7 42 4F
 F6 38 8B 51 DB BD C6 8E 65 1C 9B B0 05 B0 E5 34
 F0 C6 3E 07 4C 05 FF C8 94 12 22 E6 C0 F3 64 08
 1D DC 32 79 F9 19 61 87 EC 41 E5 AA 4B 9B 20 F4
 26 A3 30 02 07 0D DC 8C A0 B0 6B 47 5A 5E B6 C7
 8A 1D 41 BF 43 57 61 B1 A6 2B 38 FD 24 E6 AB BE
 29 C3 50 68 79 9A 6C 21 17 C9 48 5A C5 30 FD 9E
 11 79 9E 24 07 32 F2 F0 B6 16 17 37 00 21 D0 12
 61 22 E2 A3 45 5B F5 AA 3C 3F DA 8C F4 AE C2 D9
 AA 99 46 87 A1 96 EC E7 59 86 52 60 2F 2F E8 77
 F2 E6 98 41 6E C1 08 16 DE 78 23 FA B3 84 13 2B
 C4 21 1B 56 E9 FB D1 B9 3C D1 89 7A 09 C9 7B D4
 08 EF 7C 5A AD CE E8 05 71 84 EB 26 77 4C 39 CB
 5F 0E BF CD C7 A8 AB 94 D9 13 3F 6B 25 80 1A CF
 61 D9 8B C5 0E 4D F5 E6 B3 F5 4D 82 15 9E 29 10
 81 17 1B 38 A1 C0 3C 5E 65 CE 03 29 97 CF DB F1
 FE B4 0F 20 E4 3C 7F AD 10 81 B5 F8 59 1B 04 64
 34 C5 65 43 66 BA D3 59 62 AA 2C D1 5C 30 BF B2
 2E 37 01 E1 1E 23 C1 01 87 5A 4B 71 E9 8A 99 AB
 AA A6 65 81 E9 F4 6B 83 4A E3 83 C3 E6 8D FD 9D
 67 88 EC 68 83 AB 9B 83 22 F2 FB FC 8D B0 13 0D
 05 91 91 12 98 E2 AF BD 68 9F 9F CA 67 C0 3D 9F
 68 75 61 1D 0C 4E AA 2E 10 DB 57 58 86 7E 90 9A
 8C 26 AC 7D 8A A3 73 B6 35 21 1E 46 06 A5 93 C4
 AC ED 27 E5 E2 F7 79 42 DD 05 6D 4C D9 44 F7 14
 BD D5 C6 8A 3F 23 F6 CC FF 79 96 D4 17 3A 2E 8D
 EF DB F0 ED 13 56 C8 FC D9 17 CD 99 72 B1 CC 1D
 39 A0 55 EA 84 DF 77 36 3E 90 8E 90 65 20 A0 07
 B6 96 74 CC 6F 72 56 64 4C 0E 95 41 61 D0 D9 38
 06 0D A3 53 C3 96 C1 3E 33 A2 5E 54 EA 83 F5 12
 A5 5A 8C 56 BD 1D 5A EF B8 59 E4 3F 0C DE A2 53
 BA 7C D2 4A 59 BA 71 45 3B 4F 17 1F 35 E5 D5 B1
 DF F8 95 44 9A A1 F2 99 B9 68 AE B6 90 E0 AA F0
 39 A2 E6 C3 BB 85 6A DD 86 6B 81 EC D9 35 15 98
 B0 51 AC 08 11 B9 25 0A DB 49 C4 FC 4B B4 D7 97
 2D DE 54 2B 43 AF 3C 35 65 89 B2 76 42 90 C8 48
 C6 BB F6 4C D0 23 55 79 1E 38 07 81 95 3F 3E 15
 91 D5 A7 DE 86 49 4A 93 9C 94 A0 02 7A 7C DF 13
 20 9E 9D B3 5F C3 F0 86 5F DA 27 CA 5A F2 62 C3
 DE 15 CB 52 A6 76 8C B6 B9 1E DC D7 8C 78 02 6C
 E0 5A 33 BD F6 7C 88 D1 F1 92 FF 5C CE 80 B7 FB
 86 3D 7D A4 49 05 84 FC CC 09 4B 36 5D 31 CB 6E
 BA 4A 99 F1 43 D1 DA 18 20 D0 D1 FC D6 8B EE 1C
 1A 23 A3 2F 68 17 29 ED 37 C0 BF E4 45 5E D2 2C
 69 47 36 D2 84 56 C8 7B 4B 7F FA 93 80 26 BE 6C
 95 A5 27 76 0A 70 AB D6 FD F5 36 5C EE 8F 80 D7
 1A 9D 4A F4 51 DF A5 DE 78 3F 0C 55 6A FF ED C5
 E5 90 90 D9 A7 14 9A 66 1C 58 95 F7 A3 B9 57 23
 D8 8F 5E 73 27 E2 4E 70 4F C5 0B 8D C6 76 C5 1C
 0E 05 40 4D C7 17 1B 82 D5 F1 0D F2 D2 D5 9B EF
 76 68 29 ED 16 2D 12 F4 EA 00 5E 7F E4 D5 6E 0E
 02 75 E5 1F BB 1D 89 2F 04 41 49 27 94 85 1A 18
 52 7B 90 D5 E7 6F 80 BF 4A 0E E9 43 52 6F 63 57
 29 08 69 90 B5 8A B4 B0 C6 2F 44 BA 4A 7A 13 9D
 51 6B 4F 7C 40 AB D1 73 4E 92 AE A9 F0 E9 DF 1D
 7B E6 BC EB 31 25 E0 9B AC E0 2F 6A E6 37 7C 3E
 60 44 28 F3 E5 97 D3 D8 00 DC 86 8E 04 D2 7C C1
 7D C2 9E 52 6C 94 A2 7E F5 B5 1F 6B 92 D3 FA 21
 78 84 F4 C4 0A 5F 8C 12 96 FF B6 CD 36 1C 96 A1
 CD 79 45 D6 53 9C 1E 2E C4 8A 6E 08 CA 1C B9 8F
 D3 35 06 7A 95 55 CF E5 6B 32 1B BB E2 94 00 9F
 2D 2F 5E AB 7F BE 89 FC 87 EE AE 3A 38 26 13 37
 C2 E2 3A 14 B7 53 8A 8C C6 AF 48 94 6A 62 F4 77
 D1 C3 0D E6 05 69 A7 03 19 91 8C 6B 98 77 07 4F
 C8 4C 16 FA 48 70 3B 84 6E 96 6D 43 1C B3 2F 7D
 69 98 E5 A4 C9 A2 11 E6 A1 F5 45 CB C3 F5 D0 26
 6F C9 5A 19 C8 F8 42 00 DD 44 9C 61 BA 51 01 1B
 62 42 33 69 30 98 6D F6 0F 46 05 15 BE 78 D0 C9
 D1 D2 79 BF 96 A4 0E 6A CB 41 AA 51 26 73 BA 10
 6C 94 0A BD FE C8 10 46 86 0D 3C 24 F7 92 47 FF
 87 8C 13 D3 7E 97 85 9C 0D 9A E8 E0 7C A1 45 AD
 5A 0E 50 34 7C 97 20 90 C6 EE 1B B8 6D EC 4A D2
 5B 02 77 DE B9 DB 63 9B 93 CC 33 71 D4 FC CC 2B
 0D 6B C1 EA 6D C0 CD E6 D4 4E A5 4A 1B E8 4B E9
 DC A7 2C 39 FC A8 D1 79 F8 3D 02 BD 0F EB 04 BA
 7A 8F 96 B8 A2 BF 74 A6 33 4C 4B 5C 04 8D 09 77
 06 AD 1E 81 1A D2 BA 75 3E B7 D0 FA 59 91 4F BA
 D9 F6 9E 1E 49 6F 54 DA CC 93 B1 1B 79 BD 8F 5C
 FE EB 5A AA E7 1E 9A CD DE EB 7A 5D 83 97 99 3B
 95 45 17 2E 0A 7F 24 6C 24 F6 79 46 16 38 CF 09
 C3 CE 16 A4 3D AE 5C 8D 52 58 3C 8F 1B 01 36 72
 60 E0 4E DD D8 46 E5 7A 22 9A 9D 62 BF 6C 96 AE
 CB 32 ED FA A7 58 85 24 A0 9D DD 62 95 41 EC 76
 CE D6 A5 90 B6 BE C9 87 88 C1 9B 55 FB 54 38 27
 5A E0 27 50 CA A5 25 3C EA 12 81 99 4D 8C 76 35
 69 1F 2E BB C7 64 B5 AC 03 30 4D C6 96 D9 6E BC
 76 BC 6F 95 78 71 4D 0F E1 23 DB 22 ED E2 AE 39
 2F 63 83 7F DE 91 A6 A0 BC E6 97 93 9C 13 4C 9B
 57 9A 68 BB 1C 8A 12 D5 08 E1 68 46 37 44 D3 12
 C4 F5 86 83 BC 2E 45 1A BC 69 A3 7A AA 15 D3 23
 DB 1C 9C AE 6C 1F C9 38 AC 28 52 F8 93 3C 45 2F
 B5 B3 15 22 11 80 19 F3 96 38 86 97 82 20 B2 06
 BA 6B A1 F4 8E 8C 34 97 8F 90 1C 31 2F E4 94 35
 C1 F7 97 E7 05 3F 34 EF E8 E6 D0 99 B1 CE A6 47
 F7 D3 8F 86 84 30 64 58 A4 DD 99 BF 93 6B 1F 75
 B0 E4 15 20 04 C5 DE D2 52 E3 A2 23 A3 61 C5 ED
 C7 3B 13 24 8D 6C 80 6D 6E 31 D1 85 BB A4 BB CD
 34 BB B5 3A F2 95 3C 9F C3 1F 8F 2C A1 2E 75 9C
 87 E1 DE 3A FB 2E D4 BC DC F5 3F D3 F3 42 27 2D
 03 00 A1 78 E1 71 F5 2B 5D B4 74 25 EE 38 A9 A3
 4F 4A 0A 82 F4 A6 F4 7C 77 38 71 76 37 61 2A 12
 53 99 B6 54 28 E4 41 11 73 1B 69 38 22 D5 AF C0
 76 33 93 CD 03 0F 71 25 3E ED D6 BB A7 A9 08 4F
 FB B2 5D 3F 63 1C 74 82 F8 B7 E6 8D EB 2B 95 94
 F5 D4 9A 68 33 E6 4D 39 85 1B AA 21 4E C1 54 5E
 84 81 0A 19 4E BE 32 A6 A0 DC 46 10 68 6A 56 52
 3F 8F 02 90 0B 52 0E 72 B1 F9 94 9A 55 5F 56 EA
 A0 B9 E9 7A 2B D2 FB F2 DB A1 F5 2B 5D E6 B0 14
 65 08 43 9E 4B 75 BE 8E 5F 2C 82 73 76 F0 90 DD
 B9 57 96 51 2C DB E3 4B CF 6E FD F3 69 BC 02 8B
 20 05 0D 31 A2 5B B2 AB B9 D5 62 C1 3C F0 1B AA
 E0 EA 43 C3 D1 8C EB 00 85 D3 CB 4B C3 EF EE 12
 6E 84 CD A2 50 64 5A 6F A0 20 6E 4B 19 DB 10 07
 32 10 6A C6 86 98 8E 6B C7 4E AE 0B 2E C2 D5 BF
 EE 88 BB E4 55 E3 96 6C 5C 2B 00 11 4F 21 6E 3B
 E0 04 6B DB B5 DF E0 A4 2C 36 44 82 46 71 CE 82
 46 91 75 45 D7 78 FA 4E C0 D3 2B 03 C1 6E AF 3D
 1F 3D 0B 88 F7 EA 9D C9 A2 F9 60 F1 EF 28 E7 32
 9B E1 A2 B8 FF 15 62 E1 71 FE FF 72 AF 2B CF D1
 A7 25 91 DD 3E AF FD 7B F7 1F 4F 4A E7 59 0D 2C
 F5 77 C6 A5 29 E5 84 E0 1A EE 9D 90 F0 C2 ED 56
 67 F7 87 03 25 43 A2 8C 4F A0 F4 69 CC 18 33 2A
 FF 6F 9B E7 D8 3E 64 AE 94 54 A8 33 38 4E DD 52
 A0 DA 6D 94 E1 87 58 0A F6 6C 4B 49 8A E6 23 EC
 88 F2 33 D5 DE 34 A0 51 D4 A0 52 E6 EE 3C 06 59
 6F CF 88 3A 8B 14 C5 6C 2C 04 8B 78 DB AA D7 85
 EC E8 AF 0C 09 D9 2A 55 9A 1C EE 87 AF F8 6B 1C
 9E CF ED A0 BF B4 4B 43 EA 30 EC 3A AD EC 77 4A
 ED 8F 94 19 4D 7B F1 0F 47 94 4E 36 39 12 27 8C
 30 F0 4E 7B D9 09 F9 2B 7F A2 44 77 91 D7 1D 11
 56 A9 C2 A2 30 7B 0C B3 CD EA 2A 66 6F 39 41 BD
 7E 14 B5 3F CE 7D B2 F5 32 92 C2 C8 EB 64 D5 34
 EE 74 7E 6F C9 70 4F 4C DA D7 64 AB 1E D5 FF CE
 8F 9A 67 13 67 82 6B 14 26 AE 19 1F 0F 16 C7 68
 77 8E 6A B0 DE C4 6B 3B CF 97 B1 34 2B 2F 76 23
 A8 4C 19 63 39 36 DD 60 D9 69 EE 31 EE DD 52 62
 5E 12 DE 0B 97 31 38 2A 42 60 9C 26 88 04 32 DF
 37 7A B5 1A BD 66 B8 20 33 FB BC 1E 6D 0D 5B 79
 D3 BC 1B D0 63 A4 36 E2 AE 85 B9 1B A0 8C 88 37
 3B 92 E1 B6 63 A3 C2 63 17 03 68 D9 A4 11 CB C4
 16 47 BA C9 1F 00 4F 7E 9D 7F D0 B8 97 11 7B 52
 30 EC 70 78 FD 04 25 06 F8 08 12 66 3E EA A9 94
 6A 65 6F DC 51 38 F4 D1 94 4B 0A D8 A6 04 70 23
 86 CF 82 27 FB EF 12 98 F9 E4 01 77 25 CC 75 B3
 5A 1B 2C A2 9F 90 A9 85 62 00 F7 14 33 09 C2 65
 2B 09 2A A0 AA E4 C6 32 E1 63 FE 9D B2 87 AA E0
 AB B8 28 47 9B 5E 0A CF 5B FB 81 52 23 08 7E 39
 24 CE BA 96 D0 BA 85 16 A4 DC 3A 0E 20 1E E0 ED
 83 8F E5 9A FC BB 04 00 CC 63 73 34 9E E0 CA 9F
 37 50 C2 2A 59 CA CE 3F EB A1 81 0B 3C B6 21 5B
 4F 1E 1E 24 E8 70 8E A4 3A 74 8A BF 8F 33 54 75
 15 AA 51 80 CB 0B B4 F1 6D 6C B3 15 A7 2A F9 08
 76 4B C2 23 3A B6 88 25 0E D5 BE A5 32 7F 08 70
 EB 58 74 DB 07 FB DE F7 F9 21 9C 22 48 5C 8E 5D
 6E AF B4 D8 99 85 63 D0 09 01 3E 6A 93 9C E6 C8
 A3 86 02 56 F6 8A 02 F2 9F 6A AD CC 2D CA 7F 6B
 D3 FD 74 63 8F 27 7A 5F 9B 0A AC 2D 15 38 61 77
 55 88 63 EE C2 5C D8 EB AC A5 3F E4 AC D9 F7 74
 DB 01 D1 E4 C8 6C 31 4D 4B 33 52 00 32 93 BB FC
 13 EB 66 D1 83 E2 B8 FA 86 3D A7 9E 8D EC BB 41
 24 F0 D3 BF 8D F7 0A 45 5C 86 F6 80 95 7A 10 A0
 23 29 0C FE 68 28 1E 9B B0 3F C7 78 FA A5 7A B0
 B2 A0 5F 50 63 3A CB 8F 69 8B 92 FE D2 8C 9B 75
 47 0B D4 FC 66 50 2B C2 1A 37 29 C4 23 1E 6E 9D
 9A 7A 97 D4 BD A4 C4 7F B8 12 FE 50 CE B7 03 1A
 59 DE 02 FD 2E 65 15 00 9B 46 1C D3 F6 F5 EC 7F
 6C FC 71 FD B1 31 59 AB E0 7C 78 2C CC 30 57 8C
 19 9F AC 43 49 3B 9C E5 1D D3 ED 81 13 67 FB C3
 F1 C9 18 4A 32 15 3F E7 05 40 D9 E2 61 17 A8 BD
 7C 4C 0A 52 3B 02 EC A9 22 78 2D D7 F6 34 2F 10
 52 00 53 B4 92 3C C4 E1 7B AC 47 DD D0 08 65 7D
 22 7D 62 AE D7 B0 68 F1 7A 1E 29 F4 6D 8E C8 F3
 E2 48 1C CA 23 F0 0F 44 01 7B 07 31 1D DE E7 87
 4C E3 2F D5 2B 94 3C D8 5F 0C 87 E3 DA 11 9D 5F
 09 8D 43 DB 3C 26 CC 6B EF 59 BB 99 DE A9 4B 2B
 64 08 3B 3E 4A 33 18 01 B7 72 F1 7C 38 0C DA 50
 68 C1 F4 F9 9A D2 9A 1D 10 F2 17 C3 DE 00 37 4E
 07 7E 1A 11 FC CB 65 3A 59 F8 8D 4E D8 BF 32 FC
 55 DA 52 5E EC 74 E6 14 B0 44 A8 D2 45 93 4F DC
 88 64 A5 14 0D E7 57 E9 37 E7 19 89 DD 14 7B 83
 5E 4C 73 2B 90 73 39 43 B6 BF 04 87 7E F7 74 B9
 16 2D B7 F9 8F 45 09 7B B9 7C BF BD 79 41 6A 1D
 17 BD 64 A8 2C F0 DF AD F7 37 7A B4 C5 3C BD AC
 D4 AC 67 D8 24 8A 46 06 E5 DE A0 E0 99 F2 49 F2
 DE 8B 97 5F 55 FC 7F EE 1E 0B 22 C5 61 C7 AE D5
 BB F0 DA 29 AE D6 DC DC B5 0B 3E 2B 57 99 A0 F8
 3D 05 71 68 F5 2B B8 F1 22 FA C2 CF FE E7 DB 4D
 29 65 12 51 EF 32 8B 36 34 4A 04 49 97 0D 0F 5D
 A9 BF 71 3B 7D 78 68 90 D8 36 2A E9 37 74 6D 2F
 86 BD DF 62 22 2F 00 F1 C5 72 4B 94 86 3E 1E 28
 6B 1B 7E 28 C6 10 0E EF 72 96 40 B0 4C 84 D2 F5
 53 71 AC D8 F5 25 DE 5D CA B2 BE 0B E0 2E 0D 79
 8B 02 0E 3B FE CC 9C 48 F1 5B E4 B4 DE 92 BB A9
 63 59 1F 53 12 5B 7E F4 E3 FF 0F BF 1F B3 7B 81
 CB 9B 20 35 60 5A 62 C8 F8 BD 1C D8 4A 85 80 9D
 3D C1 85 B7 2E 00 E2 61 D1 61 54 27 61 5D C2 D7
 83 3C D5 B7 A0 A3 78 35 58 8D 57 86 7F 0B 68 3F
 01 EC 5E 01 FA E5 FC F5 3F EA 01 39 B6 EF 3A 9F
 2C 27 75 EE 3F 36 3E E8 69 9E 3F 6C 25 F1 5C 5D
 F0 5A CC A1 51 C4 70 DB 17 39 72 CB 43 28 40 9C
 3B A4 54 D7 35 34 DF 3B 57 0B 06 6C 20 2A 66 8D
 83 73 0A 89 96 A8 15 A6 F3 7F 76 FC 97 B6 36 F4
 C3 5B 5A 94 43 14 DE C5 2F 96 5A 96 57 44 6D E2
 47 32 E7 19 38 0C F7 80 71 79 25 1D A1 05 1E 05
 70 FE 21 E5 D0 E8 C5 3E 27 46 71 5A 56 52 90 4F
 86 06 F2 3B 9A D4 73 AD 7B 50 4D 2F D4 E0 3F 11
 7E 77 52 92 A1 14 FD 67 7F 07 5E F8 86 E6 D1 C6
 80 92 8A 93 79 5F 64 83 C6 19 5E 19 FF 73 C9 68
 67 DC C3 F1 12 69 7F 0E C8 DC 29 94 6B 74 95 59
 1F 20 50 8E E5 35 8C 02 31 75 E2 D5 67 97 73 05
 3D 42 AA 68 FB F8 08 A9 96 DC 3F 1B 5F C9 4B C1
 F8 1D 1E 9C 76 33 53 14 B0 8D 60 91 64 02 54 66
 6E 45 21 DE 55 65 42 C3 2C 82 25 2A 47 62 0C 55
 23 EC 4B FA 52 15 9C 86 01 28 01 6C 2A AD F2 72
 11 80 01 5C 6A 45 1D 30 33 1B 87 DE 82 62 08 29
 B0 AB C5 3F FD C3 51 44 D3 6F 4D 11 8F C0 23 F6
 C5 C4 91 96 BF 66 B3 5B 91 C2 91 AA 3E D1 E7 D3
 5C 73 58 20 0D 1F 1F E0 90 AA C7 7F DB 68 C4 1C
 36 3C C3 ED 12 2F 71 2A 91 2E AA 52 A9 4D 70 B0
 AB 6A 9C 19 37 1C 12 58 0A 35 F3 A2 BF 0D 4C B2
 68 E7 14 4B BE 3B CA F1 6F 4B F4 26 70 11 FA 2B
 1B 39 95 FF 3E 5F 64 7F C6 DF BD F9 08 3A 0A 03
 E2 EE 3C DC FA 7D F5 99 E9 B9 F7 93 49 4B 2C 22
 C6 E4 62 76 CF ED E5 78 03 AD F0 7E 05 B8 A5 67
 42 DB FD BF B9 5C B4 06 FD 49 92 AA E3 A5 95 1F
 F6 88 BE 71 6A 6A C7 28 90 6B D7 B6 AE E6 5F 67
 FC 3A 3E 02 0A 2C 69 98 89 2C EB 6E 98 89 03 09
 1C 11 EB 1F 4B B6 D9 E3 0B CB 67 A2 83 40 26 A2
 5F 3B A9 11 BF 32 E0 6F 59 14 04 F7 1A D5 CD 37
 29 70 CB 00 63 64 C1 CE DE BE 4D 5C 9D 9C FF E5
 D3 00 A1 F1 09 BE 22 21 EB 62 CE CD 1B 48 60 7C
 D9 A0 F2 6B BA B3 D2 8E 61 4F A9 C9 1F B7 E4 8C
 1D 56 B6 56 05 10 C0 6F 4D 38 50 49 3C 06 A7 A9
 B6 C3 DF 59 53 F5 F4 5F 02 66 78 01 02 6B 8B 48
 41 23 13 BB A1 66 35 33 A1 F8 D9 B3 7C 4A DD 87
 20 B4 E2 EE 00 24 58 C1 4A 07 67 C1 A4 71 54 5B
 B1 04 78 3B 60 1D DB 1E D3 EE 1A 0A 4D D7 F5 FB
 9B 65 FC AC EB 5D 21 5D 98 FC C4 D7 CC 05 82 DF
 C0 E8 96 C4 64 AA 86 52 6F 4D CC F6 30 ED 97 15
 4C E2 E9 01 70 25 F7 D0 6F 71 EE 34 BD ED 18 A9
 93 9F 79 D7 8F 3B 63 50 EF 1F 47 A4 9F 1B 08 70
 42 94 95 DB 40 3F 8B 4F 21 F9 5C C4 10 95 15 63
 15 E0 AD EC D2 B9 D5 42 6B 1B FC 2F 1C EF 46 B2
 45 F9 70 36 20 AF 53 02 6B FE 39 71 A1 40 FF 28
 E1 6D 6E 85 35 B7 8C CE 93 FF 3E 11 EB 72 A5 E7
 87 C6 28 80 B9 8A 4E 5C EB 0F DA E6 1B 4D 42 EF
 48 86 CB 04 7C 4C 8C 26 10 99 D2 27 26 02 E4 32
 B3 BF 35 DF 85 6B B0 E7 95 0E DC 52 BF 35 F1 83
 ED 45 B9 5E 2A F3 26 1C 0F 59 45 82 59 D4 A0 D2
 2C AA F2 E7 74 F5 4D 72 AF 9B 06 E6 C5 BA 4E 16
 6B 8B 3A 26 B4 E0 9E 73 AF 16 A4 4E 82 D9 44 14
 C8 51 0B 6E 6E 36 FF 3C 68 BA 34 10 18 AD A6 97
 DF EE EB 60 CC 46 E3 C9 32 67 22 AC AF 8B A1 7D
 4F 43 C1 B6 F4 11 F1 E1 E3 4D DB E7 41 B6 B0 DF
 C7 2C 1B 1A A4 28 F5 5E 29 35 74 7F 8E 2C C4 EA
 16 12 7E 26 26 CB DC F1 B7 6D 03 9B 2B 47 52 4B
 52 15 2A 6C 31 4A 80 FD E2 A8 1B A1 99 16 72 F2
 95 3A C8 C0 EE F7 3D AC 39 4F 98 61 4D 55 95 31
 36 27 35 19 F3 DE 5B DB D9 8A 5E 2F C0 42 DC 70
 07 E1 BA 94 19 6E A7 E9 C4 AA 42 96 EB 0A FB 74
 30 E0 0E B2 CD DC 86 AD 92 27 71 4B 69 63 8D 79
 CC 19 46 A9 B1 1F 68 08 DA 46 DA 3C 8C 15 BB 1A
 FE CE 6A 07 F1 B0 A5 F0 FD C4 DF 7D 1A F4 4C ED
 4D 85 6C A1 29 4C DD 2D D4 4E 9A 95 D8 69 46 E8
 82 4F 09 9F 03 4D A5 91 3B 96 05 E8 DA 2E 32 C0
 9D F1 46 DD 8E E6 2E C2 3B 63 BB 9F AF C5 D3 8E
 F7 97 C3 C0 94 B0 BC 4D 29 37 92 7B 52 D4 CC 6D
 82 DA 03 63 F1 3B 49 4E 7D B2 78 04 A3 AE EA 56
 46 05 F8 63 B7 BB 32 44 2C A4 02 F1 6C B6 99 BB
 CC 4E DC 64 FC D9 5B DB EA 4C 5E 5C 78 72 45 D5
 5F 0A 90 8B F9 B2 F0 96 F9 02 BA 89 B7 0B 9B E7
 3E B4 DA 4D 04 B9 08 BF DE 76 85 AD ED 81 5E 32
 28 45 36 03 37 D6 FE 33 FC 98 FB 92 88 C8 86 90
 DC 5B D7 E6 FF 02 0E 7C B7 1C 71 D9 DA B5 C5 B3
 8B 26 84 A5 F1 3B A9 BC 16 92 8B 21 D3 CC 9F 83
 EB 3E 9A 0B 67 4F 01 EF 0C 87 73 D6 C0 EC B1 BD
 92 BD 90 A8 8E 09 7D F1 8B BC AC 1A EF 8C 63 B4
 94 24 58 2E 2E BB 67 94 8D C3 E2 1D D2 27 B9 64
 0B 72 B4 92 D0 C9 F8 78 5A 2F D8 8E C4 93 5B B8
 B1 BC 00 37 F7 7F 12 2E D3 51 91 6F 88 43 9C 72
 19 98 1B DC C8 81 9F 1F D4 8C A4 95 1D 1C 31 23
 4B 73 2B 7D 6A 05 0B 4C 33 F7 DA 91 EE 0E F0 F7
 69 79 25 AE B4 B6 75 20 4B 9E A7 7B 6F 25 71 7F
 8B A3 AA 92 CA 8C EB 47 F8 B6 DF B0 8C 26 B8 8A
 71 6D 6F 3C E4 C1 3D 7D 15 E0 02 D5 73 64 A6 64
 9E 27 9F A1 7F DF 5D ED 69 FF 21 99 D8 52 85 9B
 9B 55 6C 98 D2 71 A8 F1 3A 74 C5 0B 74 80 2F AD
 A5 83 D3 D3 27 67 EB A7 32 91 50 1A 09 76 36 0F
 6A 29 BA 3A 16 5C 35 3A 72 BF 56 FC 1E 18 8A 5A
 6A D6 89 B9 64 CF 60 3D 53 4B 88 A1 B9 12 B6 07
 F3 BE 5B D1 CF F0 BB D0 D5 6B 34 37 0C 48 B6 28
 69 6B 48 E7 4B 50 93 02 FE AF 37 68 44 90 85 28
 40 ED 4A D5 67 92 56 B7 0C CD 63 84 23 4E 9A ED
 6A A3 9E 18 47 2B 54 BB BD C9 8F E5 80 B5 0C 7C
 44 53 2A 4D 00 EC 54 94 6E A7 DA C1 17 09 3B 62
 86 02 E8 8A 29 47 11 36 88 4E 87 1C AA A3 71 10
 EE C9 6C 81 50 78 EA 8E 91 E0 37 03 CB 0D 39 B4
 5E F6 FB 2A C5 0A 57 B3 21 53 F4 02 9B 97 81 85
 4F 3A B5 29 69 59 D9 84 D2 01 F3 62 C3 5D 53 A6
 BB 61 4F 45 0A 5A C0 E0 CA 12 FE 97 24 C9 83 FF
 D4 92 D8 85 E7 37 76 9A 8F 3C 0A 72 3A 91 04 12
 DB C2 41 81 B1 4D 1B 07 2D D0 52 CC A4 AF E4 CC
 E3 8E 4B 38 D5 39 A2 CA F0 AE A6 67 A5 4B D9 3F
 45 14 FE FB 49 55 37 A4 D9 7C 43 9C 56 9D 35 77
 10 CC 80 FE A5 62 B1 32 BA 2B 46 B9 C6 65 92 E7
 7C 0A E8 3B 20 12 EA C2 42 BD 68 66 24 F9 DC 2E
 49 C7 5A 6F 00 F8 F4 4B 37 A7 9A A4 AD 0C 74 99
 26 87 47 C5 7A 89 BB 86 AA 25 44 08 4C F8 D8 A0
 DE AD 9D C8 14 30 4D 67 7E C4 16 B1 1B EC 5A 51
 39 33 39 88 A7 4B CA EF 6D 16 2C CB 1E B6 C8 7C
 CB 5E A1 F0 72 13 65 80 69 51 67 72 96 B9 A7 B7
 D2 56 B4 01 65 92 95 FF 21 66 08 7B 1D BD B7 01
 84 66 75 3A B8 E4 7A 34 DD C7 5E FB 25 FB 71 EC
 77 F7 1E CE 5B 44 96 95 91 D3 07 46 AF DD EA A3
 AB E7 C4 DD E5 53 BD 9C D8 2A C6 CB A0 0E 4F 85
 01 61 00 57 5B D8 12 E6 8A C0 D4 85 43 44 F3 BB
 59 EB 0A 21 B1 21 26 4A 11 C8 E9 A0 83 D1 54 34
 48 B6 52 4A A9 89 FF 4F 27 AF FE 98 31 53 BA 4A
 68 5D 6D 53 1A 7A E2 9F B3 47 CD 34 88 D2 0C AE
 D3 D9 68 BC E6 28 B9 1F 9C DC 7A 56 5E BA 29 70
 D3 BC A7 04 46 27 81 9F A2 5A 35 B3 47 5B 44 15
 F6 27 3F 1C 0B B9 F2 0D C6 25 C4 29 40 DF E0 B3
 0A 82 EC 5D 83 B2 8E 5B 52 6B 53 C9 6F DB 7E 48
 29 06 64 8C B3 62 C7 9D 6E BA 7A D2 44 0B D5 7C
 62 63 91 39 AA 69 54 C6 24 7F D1 E2 D0 A3 DA 3F
 9E 83 26 3C 19 A2 07 E6 EB 46 41 04 31 4E EB 10
 5E CE F2 9D D0 0C 79 35 77 4F A5 8C 73 DB F5 81
 3A 87 A8 53 FC 80 D4 8A 0A 26 37 70 B4 0B 01 04
 18 C3 97 91 FE 2E C9 19 9E 84 5E 3D DE 55 27 8F
 CC A7 9F 02 E7 44 4B 52 F9 8D 7C E9 7F 6D 50 48
 47 07 FC 0B 6E 31 6F CA 83 9B 85 41 DB AE A4 74
 F2 6C 1B 61 37 8C A1 67 D5 E3 CE 3B 9F 3C B2 26
 8B E0 34 A0 BB 85 60 ED A8 5A 1B ED A0 2B B1 48
 27 44 74 9B 9C 3E 5E AD 50 E4 B3 91 A8 72 8F 64
 3E A2 EB BB 01 77 D4 D5 1C F2 42 63 55 01 DF 0F
 EC 4F 8E 7F DB 68 7B 79 9D 8B 04 A8 4C AE 1C F7
 3E 60 36 25 3B 1B D4 17 FD 0B 44 B8 E1 79 AC 6F
 3F D6 7B 24 39 6D E6 C1 8A 00 68 F9 EE 1A 59 3E
 0B CD 54 85 BB E8 C4 04 39 E9 13 73 C8 94 D5 DE
 5B 80 25 34 F2 6D 8D 52 7E 7F 1F 69 FC 3F E5 B3
 07 77 7F 81 0A C0 DA 99 03 C1 1E 6F 07 F6 0C 0F
 EE 9A 2C 5C C9 D1 4F D0 C4 C0 AE 1C 9A 1C 8E FC
 DB F9 31 30 67 C6 DB 19 05 66 4B DB F7 BE 10 7B
 18 31 CD 26 27 3A BA FF 0C 68 D2 AB 3C BB 78 13
 9B 3A 03 12 04 CD 93 27 F2 39 00 7A 26 AA 99 ED
 79 F3 B0 17 E6 67 EA 8B F1 8F FB 48 31 0D 30 E7
 D5 F8 11 74 DE 76 FC 89 9C 0B CA 64 7D 44 30 DC
 E4 04 EB 35 EB 11 1C 30 4C E5 BD BE 37 2C D7 9F
 F6 2F 77 77 54 C0 18 10 FD FF F6 07 B9 95 EB 03
 9C 30 D2 32 BB 4D E6 90 B7 E1 65 37 5D 2D FD AD
 FB E9 61 80 76 6A 16 C7 72 BA 1E B2 48 CF 76 9D
 3B 5B 08 AE CF CB CD 23 BF 33 CE DD 76 3C C2 94
 63 2F 15 2A 06 BB C6 76 F2 F7 80 71 DA 2B 5F E4
 D6 AB DD 06 FF 36 93 AB 1A 47 C0 7C 4B 0C 17 50
 8B 25 FF FC 95 09 49 BD 42 3F F5 D7 CE 84 7A BD
 34 69 93 C6 FB 30 10 E5 D2 0F 3E 66 A9 D7 07 B5
 73 A9 FF 32 DF A0 90 60 2F AB F9 FE 8D 37 49 D1
 B0 F9 4D 6A 45 8F 09 A2 86 5B 7A E1 45 02 82 03
 0C 0B 7D D1 77 48 31 EA 68 75 92 6E 27 6B 89 65
 B9 5D 3C D0 94 48 31 14 D6 5C DC 52 D9 1E AC FB
 92 7C 77 DC 4B 68 26 55 96 D8 FC CA BD A2 B5 97
 FB E5 BB 10 0D 40 96 DA 66 40 78 C9 67 30 95 12
 DA 37 45 DC 6B FA EE 2B 2D F5 4A 1E 6A F9 87 23
 3F 27 22 9F 8F 64 51 F4 EB 39 A9 38 1F AA 6A 84
 86 4E A6 BD EE A4 7B B9 77 D7 4E 70 79 4E 6A F2
 69 78 65 8F CF FE 93 91 5B CC BB 02 FA E9 62 00
 69 64 F0 89 E7 6E 8E 8B AD FB 18 7C 75 C4 4F 9E
 6F B7 22 A1 D7 D9 DC 49 0C 2B DA DD A8 73 D4 28
 DB 9A 6C AC 05 30 34 CC 5D D2 56 4C 9A 7F C4 56
 6D 58 F9 6E EA 60 8C EC 30 A4 CF B2 AE 23 20 0D
 BB 3C 99 AA 08 FD A8 ED 56 56 5F 8B AB 2F 5F D9
 7F 95 BD 6B EC E2 1E 25 3B D5 CC 4D 7C 24 7F ED
 EC 70 57 AB 87 CA 89 DB 50 A2 EC 15 7C 7F EB B3
 5D A6 E8 3E A7 48 D0 EE E4 EC 81 6B 25 2E 9C 60
 7F 20 F6 7C 2F 5A 16 FC 10 CD AD A2 D5 9A 3B D0
 8F 32 13 FB AE 55 66 E3 C7 7C D2 0E 43 9D F9 97
 2B C6 D1 88 AB 09 99 01 F4 69 92 99 AE 0A 4A 6B
 89 B0 D5 2E B3 B0 93 1E D1 8B E6 85 31 CD 1C 1C
 3D 45 4E A9 3B F4 2B 0A 0A 27 E4 46 14 74 F2 58
 68 4F C8 22 88 F0 C6 1D DE 8C 06 D1 A6 46 E4 13
 CB EB C3 13 4D 4C 7E 7A 52 FC EF 72 BD 2E BB 1C
 D6 AF 6A EF 81 F4 82 D3 0A C9 17 8B BB F4 B2 3F
 DF 4B F7 57 1A D6 17 02 D1 F5 F1 01 1B 6F 1A 22
 F8 EF 78 ED A2 96 DE 0C F9 76 02 65 6D 7A EE 8F
 34 CF 68 9A 2B F2 FE CE 26 B3 89 99 FA 1E 48 D1
 64 8A FB 0C 99 6A D7 71 69 0E 95 67 20 A0 AE C6
 5F 94 15 9A 05 9B 43 B5 66 9D D5 C3 CA 24 C6 4B
 28 62 66 D1 77 B3 FB E4 E4 47 0C EF C9 93 9D 52
 E3 D8 5D C4 EA D2 5F 01 42 B8 73 54 56 14 A4 C5
 30 A9 AE 73 EB 9B 2E 2F 25 48 9F 0B AD 9E FE 83
 31 B0 CE 5E 29 0C 24 45 61 16 C3 AA E7 52 B2 F0
 5D 69 02 85 02 BE 3E EF EA BB E8 9E A8 D2 75 45
 9A 52 A4 35 3B 39 57 3F 42 4D 75 1A 5D 89 81 C8
 E3 E9 07 CE 5B 01 64 8E 55 07 47 E2 71 5C 8F A9
 10 DF 64 72 22 03 38 C7 C4 FF 45 49 DA 0A A6 2F
 FD 2C 1E 2F 2A FD 86 8D D2 F8 BF 98 F0 84 76 3E
 01 46 02 3B 34 0A C4 41 49 3F 1F EC 0B 7F F7 1B
 E1 A7 A9 3E 4A 48 8F 6A 2C 35 7B 53 DF 35 ED 3D
 DF 29 F3 8A D4 EF E5 D8 58 8A 61 F8 0E 09 75 D2
 5A 3E BC DB 53 21 E4 BF 3A C4 D9 3E 1B 13 7B F3
 DB A8 82 E4 E6 21 FC 65 45 2B F9 8D E2 B2 8F 0B
 E1 BF 04 24 B0 35 AA 91 2B AE 5C B3 2E A5 EE 21
 BA 1F 72 B7 CA EE 2C 75 81 0E 65 65 39 2B A1 17
 C5 EE C1 4B D8 19 BD 0E A7 91 BA 60 66 D6 F8 FA
 01 25 0F F0 96 39 21 66 0E 79 61 1E 61 E3 0F 10
 C4 B1 CA 3C C5 0A 0B B8 35 81 83 CC 91 F2 3A 40
 A7 AB DA CC CB 5F 88 45 D3 40 63 D8 87 2B 19 EB
 5B 61 8A 25 DE DC FD C7 E3 2C 5F 89 19 8E 92 9C
 1B C6 A1 23 B9 7E B3 80 BA 8E 45 3B 2F 0A 3D C1
 DE F8 9A D7 7C 56 84 6E 76 07 D0 EF A8 C9 92 A4
 5C 65 6C 9A 53 5E 2A 94 6A 1F 6F BB 19 95 29 02
 52 E3 7C 57 63 BE 48 C7 93 9C A5 3D E1 2F 67 C2
 73 31 B7 54 29 D3 6F BA 36 40 29 61 44 41 E8 BF
 1E 5F E5 1A EA 3B 86 47 86 BF 0E B0 23 F8 81 45
 D0 CB 63 06 A0 4A 44 4F 98 5E A7 75 F6 95 2C E0
 BF BE 7D A1 07 B5 D6 8F D8 72 41 8B C6 65 62 D2
 56 51 FB 38 89 96 A8 4D D5 F5 18 58 56 7B FC 3C
 B2 85 6B 6C DD 40 3F 67 A3 B6 38 FE A7 DD 68 AA
 A0 69 6E B3 B5 4E AF A5 6C F3 86 E5 8C BF 95 BD
 CE E9 40 48 7D 47 9D DC B3 74 A3 78 BD 69 1A E1
 42 DA 61 5F 62 83 F7 A7 AE A6 23 93 B1 D4 54 77
 DA F4 13 48 5E FD 2D 56 AE F3 C7 64 A1 D2 1E 0A
 08 20 E3 9B 33 36 57 C4 21 CC 88 87 6D 00 ED 0A
 94 93 76 D4 40 6C DE D7 01 4E 61 80 4F 16 61 A6
 EC F1 44 61 E5 CE B4 95 28 46 38 52 BB 10 BA DE
 62 AA 83 F9 B8 B7 C4 DA BC B2 B2 B0 7B 8F F9 16
 DF AE 45 97 67 58 8F AF AC 98 98 28 93 B6 A7 F8
 0D 39 D7 AD A2 8B 54 CC A0 E4 BD CB 87 5C B2 F8
 B2 7C 7C D5 55 D4 3D B3 4C 5D FD 66 A9 D2 49 3E
 CA B7 52 B0 C8 A4 58 2E 0C 47 DB CC AE D0 44 52
 08 CA 85 F2 26 89 AD 26 36 72 72 96 89 9A 9D CF
 03 93 2D 80 FD 36 1E 49 03 F8 62 4C 1A 85 93 3E
 FE D6 73 07 FA 70 DD 33 49 D8 CF 42 8D 03 F3 5C
 13 BA 70 BA 11 20 72 46 15 1D 86 A4 95 EF 12 1F
 07 7C 77 81 44 62 03 DA 35 D5 4A A4 EB 1A 31 87
 18 51 4D 53 B5 4D AD 5C 43 79 EB CA 4A 15 A5 8A
 AC 9B 58 EA 71 1B DF 13 F9 5A 95 C8 E6 2C 79 BB
 2F 47 F4 8B 7C FE 40 D8 D5 B5 63 9A 54 DF AC 7E
 99 8B 3D C4 FA 8A 49 FF 29 29 A2 D4 5B C0 9F 67
 43 A3 BB 3A C3 F4 DD 60 BE 94 58 16 07 2F CE F8
 61 33 1B E8 16 BB A5 AE FB 61 01 08 6B A6 0E 1D
 45 91 C1 EB C9 F7 83 E4 4F 6A 0B 78 D8 5D 07 4E
 F6 BF 22 A8 8D B5 28 13 D4 84 48 67 58 CD 93 61
 0A 2A AE 6C D9 B3 C0 3F 0A EF 14 55 A2 66 F9 60
 9C 8F B8 8B E1 29 41 CB B4 5B CE FE 8A B3 DB DC
 7B C3 37 27 A6 F1 64 ED 30 78 06 5C 9A FC B5 06
 91 7A F0 83 0D 69 26 69 9F E0 AD F0 45 DA ED DB
 DA DE 2E E9 CF 5D FD CA 3E 37 2F AF 59 AF FE 66
 2D 98 0C EA 0F 4E 97 19 56 9D FF 9F BE D7 68 F0
 BA FB F1 6D D6 3A 5B 83 65 94 F8 82 95 04 53 01
 CF 3F D6 3C 14 D1 C5 DB 62 2B F7 2A A8 D3 19 8A
 13 93 75 85 E5 A8 B5 DA 02 D3 53 7E 92 9B EC D1
 25 47 B1 F4 F0 4D D4 E3 A8 BF 1C D6 EA 4C 07 77
 97 74 15 16 2F 87 01 1D D3 F3 91 71 E2 49 29 2D
 9A 6E 8B FB 56 DE 5B 44 4D 1B 0B F4 2A C0 C9 E6
 C1 B3 B2 10 DE C3 40 B6 DF F4 34 07 27 13 19 49
 8A 20 EA 48 CF 7A C7 61 63 E0 28 1F 5E F5 6C BC
 CA E7 66 0E 7B 26 29 28 1C 38 26 E3 82 A6 82 F7
 82 35 43 90 17 2E 8F 9E 94 F4 C7 23 30 A6 C2 9A
 6F A3 54 DF D3 26 2C BD A5 16 11 F9 82 18 B4 0D
 EC 17 29 BC 0C 83 C8 F9 96 8A B2 86 A2 4B 04 05
 E4 91 61 36 4F 3C 35 59 03 54 61 DB 21 6E 76 52
 CB 69 73 DA C4 34 1E AF E6 65 01 2E 49 51 BC E5
 EC 2D FD F0 83 4A D5 D3 6A B7 B9 68 37 94 A5 0A
 D2 B5 55 41 D8 A1 3B D4 6C 4A E3 28 6F CC C6 CD
 9E C6 F6 CA 2C A8 01 DC 1B A0 EC EF FF 87 FE 22
 38 2A 91 B1 00 5F 98 68 00 7D E4 0D E9 D5 54 B6
 FB 82 82 15 27 29 F9 89 3C 91 43 0D A8 EC FE 24
 3F F5 6A F4 38 CA AB 31 59 FE 54 B8 B3 3A 3C 3A
 42 CA AB CC 50 6A 2E F1 91 EB E7 AE 46 7C 8D 6F
 F4 C8 E1 02 05 51 01 23 24 D3 4B B9 C9 8E 67 E9
 29 1E 67 A4 67 E2 34 46 7B CC 39 DA 2C AC DE 5F
 1C 7E 1E CA 54 42 C5 33 B9 D5 F7 D2 C9 0D 1E 13
 0D 68 BA 09 94 FE E9 CD EA FE 3F 43 37 4C EF D1
 C1 74 82 F9 42 ED 4A DF 0D 91 9B 1A A8 14 1A F4
 C6 F9 3E 02 C6 53 B9 CC 22 9A 1C F8 D7 22 FC 57
 8A 2E 24 DF B0 87 51 87 1E 40 03 C3 34 97 ED 8C
 E3 54 A0 5F 2B 4C 58 B8 88 30 35 02 83 68 9C F8
 9C 2E E2 6A AC 8A EE 51 EC F4 F6 FE C6 9C F7 A8
 EE 5C B7 22 B9 C3 E7 B0 AA 2C 9A 73 49 94 C9 87
 E5 41 2E 72 18 32 2E B5 AA 54 51 B2 08 68 47 CB
 7B 67 56 3F 92 7F 53 D6 6B 71 DB 3E 04 7C F0 53
 C7 22 80 A4 99 61 A2 D4 37 05 5D 3A 80 5D B4 03
 B0 15 D4 AC 02 33 45 05 63 4C 4E 0A 34 FE 96 01
 85 41 DB 55 59 D6 65 BF 74 9C 2F B1 EF 5F 1D 56
 15 58 43 7F 22 C9 49 43 CD 91 41 BE 14 57 E4 72
 8D 43 FC 43 D9 62 83 E0 93 0F 80 AE 90 A3 D3 1F
 A2 2E AD 17 AC D4 6C 59 3A 91 E0 EE 6E 32 6E E8
 3B C1 B7 F6 74 52 68 F0 B6 E3 5E CD 8C 6A E7 DB
 3C 6B 31 90 95 C4 5A 5B 58 EA EF C9 F1 41 FA 13
 5C 7C 59 F0 78 F4 19 07 14 4D 1E 82 12 00 A3 95
 F8 34 06 08 B5 25 EB B2 65 4A E0 50 0E B8 8E 30
 B7 7C C8 A7 7C 33 B5 49 27 9D A5 98 D2 39 51 B0
 06 80 D8 D6 FD 7C 97 B4 09 47 07 6C BB F3 00 37
 45 61 89 3B 6C BF 71 46 A3 80 DA 4A 5B 4C 03 BC
 4B B8 B7 06 5C 3F 97 59 CE F2 08 F3 B9 21 50 08
 69 4C E2 D6 CC 76 E8 8E AF 18 9E 2D 9C ED 28 88
 B3 AE 93 20 4F C0 8D 90 CE 0A 44 98 C4 15 38 15
 0F 3E 4D 44 19 5F 77 3A 5A EA FC A7 20 A2 E2 0F
 1B CC BC E4 CB 89 F8 07 6D 56 FD C3 0C E1 7D 7A
 BB 4C 6A E1 33 25 ED E6 E5 2E D2 68 49 C5 21 EF
 97 EF 6F F3 48 E8 F0 50 B9 34 E5 9C 2F 66 1F 85
 DC 87 F6 57 25 44 4C 6C 07 6F D6 68 B6 EE 12 1D
 21 23 1A 21 0D 84 FD 20 7D 1B 24 32 4E B7 21 5F
 10 A6 C5 35 72 F8 E2 CC 2F 6C D9 A2 B6 D3 61 94
 B8 E6 37 B1 E5 28 D9 8A 35 C4 DD 48 07 6A BE 59
 FF A3 B8 D9 5F B4 54 48 FD CE 0A C4 A9 DB 5C 5D
 B2 D9 2C FA 4A FF B1 E3 9A 98 27 6C 2F F0 AC FE
 21 4A AC CC 04 04 02 66 99 81 9C 18 E9 3B 94 1F
 D2 4E 49 41 8D 73 38 C1 A7 8E 9D 70 A5 ED 3D 12
 8D 56 CB 73 4A 65 23 3B EF 32 DD AD 34 A6 E6 AE
 F2 13 3F FB 44 F0 64 6D BD 0C CC D3 67 B4 C8 93
 DA 2E 39 14 53 14 D4 A5 B4 C5 62 8E 78 96 DD 66
 4E F8 B3 AF 06 CB 3A CE F0 04 24 CA 92 E6 97 7F
 F5 15 5D CD CE CB B8 E8 79 82 EA F8 AD 62 06 9E
 7B 08 10 66 1A 7E 23 F5 19 8C 4E 38 ED BC D4 A6
 BB 23 02 7A 71 61 71 7A CE DC C7 A7 F4 A0 F9 17
 32 F2 68 C3 76 51 42 69 C3 97 24 F8 AB 99 3B 98
 17 8B 3F 6F 0D 4E 8E 01 A9 2F E3 83 79 58 CF BE
 2A 4D EE 8C 4D E8 D7 B5 8B 88 E8 7C D4 BA 01 67
 2C 6F 2D 97 C5 62 03 84 C5 B7 89 30 B3 8E CA 6B
 BE FE C9 64 BD D1 AD 86 46 B7 D3 DE 95 D6 29 2C
 CC 58 03 90 06 23 EC 67 6D 51 A6 3A 48 B0 95 4B
 93 01 09 42 4C CB 78 13 F7 C0 2F 2E 57 27 6E DA
 5E E8 43 FC 26 32 10 B6 45 00 A4 27 3A E1 21 89
 30 CA A4 22 BD 56 F4 D0 53 CB D1 97 1A 43 65 7A
 8A 0E 4D 6E EC 92 C6 24 7D B8 91 64 95 CE 78 9F
 70 42 FE 69 D5 7C 89 A7 A7 BB 4E 96 1F 30 55 B8
 4C 12 A3 5C 38 6A 83 E4 A9 2D 06 10 4B 40 A7 4E
 7D 6A A2 A3 F3 8A F9 51 1C 62 F5 C9 A9 B2 3F FC
 52 22 93 A6 64 61 82 2F 24 F1 61 EB 52 4E F2 E2
 EF 2C E2 F5 95 4C A5 5D 7B 3C B1 5A 48 CF BA EA
 B0 6C 2E 8C 9E B9 25 85 5E FA 2F 6B 12 6B 48 D4
 29 B7 D9 36 F0 D6 D7 D1 F9 2D 7B 77 20 BC 2A 08
 F6 D2 FE 4E B7 FF 66 AC 5A C9 1B 1D C2 AA AE 2E
 1E 5B DE 76 98 22 4E 33 4D 0F 3B 08 FB 7F F6 76
 DA 7C 07 85 0D DD A5 47 F1 48 7E FA 82 BD 8D BF
 00 18 A3 8D D8 20 4B E3 15 0F A4 18 36 21 7B EC
 6F 0B 93 BC 02 B4 E0 7D C0 0A C8 26 BF DF 1A 29
 1E 1B B2 89 9E B1 C8 25 6A B6 7E 7F 07 CF 4E DC
 D0 AC 78 69 D3 AF B0 B0 F9 84 90 69 CB 1E 1D 74
 CB 78 D2 75 5E 39 DC 04 2E EB 04 23 B9 5E 32 F6
 76 DB 6D 47 C3 82 96 9F 46 D2 8A 50 17 F4 18 47
 34 B9 C2 1A 83 F5 BE A5 72 07 F3 C3 14 6E 05 52
 64 21 E7 69 7E 95 5E B7 0F 77 08 4B 14 02 AD E4
 03 22 D9 0A E7 FD 36 AF 1D 66 AC 39 FC AE 80 2D
 4F FC 95 52 6F A7 E1 73 94 83 A6 45 75 1C 38 C2
 2B 2B 85 FF 13 7E BE 6B BA DA 63 8E 6D E0 91 F3
 ED 9C 19 96 CB 14 61 FF 4D B9 91 50 AA A0 E1 01
 79 CD D2 E4 DB 3D 8F DF B3 BA 3B 35 6B 94 1F 67
 9E BB 22 F8 F9 67 3D DC C3 45 40 67 D8 87 7F 45
 02 D8 A7 14 44 AB BD D9 23 34 4F 78 88 94 6C 12
 CE AE 7B 4D EE F1 2A CE 2B B1 3E 74 F2 FF 1B 2B
 22 0D FF 1E DB CA 41 B8 46 6B B5 88 5A A0 1E DD
 6B 23 1A 21 AB 91 2C F3 22 BF 60 B9 D7 4B 65 9C
 32 21 02 32 70 59 38 42 1D 50 67 E8 11 7D AB B9
 2D EA 57 D8 A3 12 9E A4 D0 7C C3 A4 E4 7F FD 70
 EF 13 A8 E4 11 BC A9 03 78 63 B0 C8 3B 0C 98 AF
 C1 B3 F6 37 B4 8E 57 EB F7 36 24 35 F5 1E 6D DD
 09 B1 DD AE 0C 7C DF 2C 06 11 B4 8B FF 97 D3 5F
 75 F3 36 81 0B 2C DB F6 1D F3 A9 C2 8A 90 1E 91
 C1 68 DC 9B 62 5C 90 89 66 70 A2 1D 1A B9 90 48
 F4 44 54 B4 E9 8B 2B 66 2E 36 2F 8D 49 F9 F5 CD
 22 20 4F 8C CB 4F 0B B8 9F 47 8C B7 7D 3C 45 E0
 D7 5C B5 07 AE 56 4B 5C AE 0A EF EF 32 DD FE 9D
 C1 87 8D AA 2D DD E1 02 4B CB 0E FB C7 86 38 07
 43 B4 CB 28 15 34 12 9A CC 5F 80 74 FA 74 71 F2
 5B 50 36 35 A7 D0 26 F5 12 9B 38 B1 27 D0 A0 28
 DB CC 8D A2 5F 8D 96 F5 A2 06 68 00 82 1D 9C 2B
 00 B1 2A 86 58 A8 BA 0E 7B F1 3A 72 EB 8A 9A 6D
 2F 45 CA E6 33 AA 5E A7 93 E3 76 C3 40 8E E4 42
 2A 19 B2 B5 02 8F ED 25 FD 3B 10 36 C1 CC 37 17
 13 05 42 EB 80 CF 15 85 24 26 A4 0D C4 9A DD 0A
 B5 5D 97 64 92 C3 98 FD 00 00 CD BC 17 5A 81 32
 A0 DF 1B 9F 86 6C FD B8 97 F3 7C 75 72 14 2D 3B
 7C 2B 13 CC 4A 0A 46 89 8D 7A 8C 74 E1 A4 13 40
 38 25 CB AE BE 29 1E 0F 38 4A 41 3E C4 F2 A5 56
 46 FB ED 21 85 89 A3 5B 45 AD 9F D9 33 F9 35 33
 4F A1 8D 0F 8E C5 75 25 FB 89 F8 05 23 A2 0A 60
 C9 0E 90 63 8C 6A 01 2A DF 54 6A 4F B6 2F C0 BC
 F0 EF 9B CC 2F 6D 98 CC 40 9E 39 EB 30 F1 41 56
 2F D8 A3 68 EF 96 26 25 43 34 74 04 6D A1 93 EE
 80 0C FB 4C EB 85 65 32 E7 6D E5 7D 86 F9 A9 BA
 25 CD F1 E2 74 F1 AD 03 9D E1 AD 2B 49 22 51 C0
 6E 57 2A A3 EC B7 F7 4C 48 6E 3B A1 E7 C9 C9 14
 BE 3E 85 B2 31 4F 83 E8 50 DF 55 9A 50 7D 57 3E
 E0 BC 20 E8 FB 39 AA E0 CF 1E DD 3B 8A 2D D4 54
 D4 E3 EC D7 F7 2A 79 39 C4 54 66 96 3A D1 4D 63
 B5 A8 38 15 7E 27 80 C5 F9 85 54 24 50 64 37 38
 98 C0 4D 03 0B E5 97 B0 F6 5F 42 6B FA 47 2E 26
 7A B0 77 AF 4A D3 4E C2 33 7C 26 BD CD C9 25 D2
 23 42 F6 A2 15 E6 BD 44 6A 95 62 E5 B1 85 82 D3
 42 2E 45 CB 62 3D FC 35 23 25 C5 35 72 5F E1 D4
 16 A7 A1 36 5F 7F C9 50 D7 8D A5 00 B1 D8 5E A7
 32 39 A0 A2 EA 37 F1 6C 96 EE D5 4B F0 9C 46 A6
 CD 5B AB 55 8E 55 FD B0 7B 3F B4 7D 7F 3A 27 FF
 2E A7 2A 73 A4 DC 96 A8 07 3D 3A E2 5B ED D9 35
 F2 3D 86 BF 1F D4 EB 04 07 C5 E0 41 8A 37 32 B3
 C8 2C AB 79 E1 1C 4B 12 6D 78 1B 84 63 10 0C 4D
 F4 5A 4C B9 70 BD AF 44 E7 11 74 03 69 D6 EB 8D
 FE 6A 8D 57 90 5C 29 15 4F 51 BA 4C 19 10 FD CA
 FE 05 82 82 BC D9 1D AA 8A 1E 9B 6E F7 81 15 CD
 CF 99 91 16 50 E5 F0 A3 DC 2F D5 6F 40 FA 29 C3
 5E 63 A4 2A 00 29 9F FB DD 37 59 15 30 F0 5E 82
 BE E9 49 23 07 82 FB F0 5F 73 FA 3D 40 51 4C 82
 96 60 53 D0 DD 95 E2 71 15 6B F9 91 1E 70 D1 D2
 0D 62 62 58 2F D1 8B 0E 08 46 FB 41 C5 2D DA BD
 49 AD AB 54 5C 19 40 37 C7 0A FF E1 2C 2D 61 AF
 7A F9 DE 34 B8 CC B4 65 70 7F E6 69 CD 39 F2 20
 53 55 B5 CF 2E C8 05 91 DF A1 F0 5D BE 5B A4 63
 52 FA 16 2D B6 EC 5A 4D 87 17 02 80 4A B5 99 FF
 36 74 8F 23 5F 92 18 13 57 57 F1 FD D8 8C 77 DB
 4A DB 6E 3B 87 AC 2F 01 E9 69 C0 2C 2D 16 6F 16
 A4 03 A0 98 E1 D3 B0 25 3A 91 EB 9F 73 3E 50 7D
 5C EC 0E 3C BF EB 13 0E 46 46 A3 7B 39 E2 92 4F
 1C D2 73 B7 99 20 EB 1C BB AD 52 62 E5 1C 98 16
 66 CB D9 3F 0A 46 23 3B 4C 78 B0 17 02 0A 7A E0
 EC B5 40 E2 61 D9 D9 A5 71 9B D6 E1 6E 2B F2 B1
 4E C3 DC 49 3E B5 3F 84 0B A0 FB E5 40 95 83 18
 D3 5A FD EB 6A C3 74 78 A1 BB 1C 82 FC 1D 56 A2
 6C D1 E4 94 9D 6E 51 CA 1C 82 3A D2 92 4A 28 C5
 B2 A9 3D 8C F3 F4 D8 C1 EA 5B 33 04 86 A3 D7 FD
 2D D6 36 8B 28 DB D3 FA 3C 74 90 95 FD DC A0 E5
 71 FC 9C A3 FD 12 E7 9B 87 B7 EF 03 81 B1 DA FA
 88 41 EF 3E 38 C2 28 92 6B 72 84 27 E5 26 20 F5
 C4 55 95 96 B6 07 59 BC 4F F9 FB BD 89 35 9A 53
 4D F3 48 F1 D7 86 39 10 FE F0 F7 0C A7 6F F8 F6
 DF BA D6 D1 C0 A2 23 EC 5C 85 DE 3B 9A B3 AE 8E
 4C 42 E4 BB FB B8 F0 7C 43 20 D5 29 F0 46 D5 D0
 CF CA 05 29 65 49 E4 86 6B C9 EA 02 97 6D D9 7F
 40 18 80 D4 88 D7 26 00 7B DE 4A 96 C3 59 AD 66
 12 0F 09 31 9F 0D 5E 6D 08 53 65 CD C6 65 97 AF
 85 72 66 80 62 36 17 11 E2 8B 04 FF 70 79 2E 92
 02 E6 3D 82 FD FD 94 C6 88 A5 D7 C4 FC B7 B6 D6
 59 14 2C 9A 62 09 64 45 00 91 AB 00 B4 2E 29 DC
 76 9E D0 05 EB 62 D2 47 51 DB EB B0 FD 4C 59 CB
 40 26 1C AA 94 51 61 DD B9 8F 1B FC ED 69 29 8C
 FC 42 95 EF 05 84 D1 63 F4 4D D5 4E B0 DA 2D C6
 9C BC D4 61 08 A5 A5 72 73 57 77 8C 7A 57 AB 98
 1C 9D 0B AC 56 92 BC 75 78 DA C4 5E 8A 95 48 FE
 BC 57 6E 50 CD 7F 2E B2 A4 0E 64 68 B8 34 56 33
 62 DF 71 81 D7 10 BA 4E E3 C2 7F 5D A3 AE 85 94
 96 8E 9A 79 12 F5 8B A6 D1 22 81 B1 24 CA AB 1A
 43 8A C4 7B A4 EB C6 AB 1A 05 A9 05 8F B0 45 09
 DB 1B 11 CF 44 B0 AF E3 7A B0 71 6C D9 DC 09 1C
 87 8D 38 F1 2C D7 1E 7F 00 A8 1F 85 E2 5E 55 88
 39 C8 0D 3D D1 57 C0 ED CD 7F 4B DA ED 73 B2 48
 4A 81 1A E5 7A 6E F6 40 64 66 B1 25 3B FB 62 C8
 0A 54 F8 4B 92 16 E7 FB 8D CF 3F D5 6C 12 7B C4
 88 F9 39 E9 BA F2 1B E4 F9 E7 E9 17 17 B4 ED AD
 A4 A6 76 16 01 BA 14 F0 FE 63 20 12 4F 1A 3A 04
 B1 FB 40 75 4E 44 32 B2 A2 96 96 11 6C AF B0 45
 BC 09 D7 97 DA 56 38 ED 0B E2 4D 37 39 F4 FD 41
 FA 91 C8 B1 B6 48 4D AB 01 FA 36 F1 7A A0 16 F1
 6F A6 AB 25 39 41 1D F6 AF 6E DE E5 8A 73 41 80
 33 73 00 95 1F D6 93 E7 E9 5F C4 62 EE AC 8D C1
 9B 79 C7 CD 32 9D 58 D4 5D 25 C8 30 96 88 CF 3F
 1C E2 96 D0 A7 03 3E 3A 85 C6 93 31 F1 D7 0D 36
 B3 D3 55 B4 AA 7B F9 8A E9 B9 92 C6 1F 53 19 A5
 7C 00 D0 5E 0C 28 9A BB E8 E1 D2 42 02 9B 48 87
 EE 83 48 4B BC 31 90 8E 41 4E 7D 5D 47 B4 7C D3
 60 52 71 84 F7 B3 44 A4 24 B0 6A 2A 94 1A 30 04
 4A 00 B1 5A 80 4B 07 34 FA D6 DF DD AA 96 87 30
 CC C6 70 46 04 4C EB 94 57 C7 7E 8E E4 E5 FC 88
 C0 66 4C AE E6 D0 E4 63 46 18 05 29 80 24 FD FA
 BB 07 05 D5 4C FB B3 60 7E E3 D5 48 F4 2D EE 77
 96 2B 2A 57 72 A7 F2 A8 90 96 92 65 F6 00 5C 98
 ED CA 24 E3 A0 85 2C A5 9B F0 59 F5 A6 3D 7E 41
 53 28 B6 BF 95 7F 70 9F 51 51 D4 42 66 B9 CB 8E
 61 F2 03 33 19 82 B1 92 51 D3 20 23 B0 F0 4C 50
 88 B8 8E B1 5A 11 5D 33 07 CF B8 B1 34 50 B1 02
 28 81 8B 36 F9 7F 82 D2 8A 44 F0 BF F6 93 B0 D1
 B0 53 94 C6 C1 83 2C 23 40 9F 72 19 6D 27 67 C7
 7C 44 9C 98 AA E6 10 FC D8 58 3F 61 B5 88 58 E4
 89 6B 09 7D 3B 71 F3 71 B7 0A C8 92 2F 9D C5 4A
 E0 74 81 10 6D 7B 44 71 13 C5 06 F9 DB 87 10 3D
 18 A0 D8 EF 49 0F 84 F3 94 A2 1A 6D 34 CC 66 59
 6B C6 46 78 28 CC 7C 62 BD EB 17 34 05 5B C1 83
 C2 F7 C7 E1 5A 64 CA EE 14 3E C4 F4 E0 53 7A 84
 23 10 3F 59 04 41 CA E5 42 3A 56 91 07 18 E6 1D
 4B 6A 1D AD 6C 5C E4 46 95 0E C6 BC 0C 0B 1C 8C
 9F 3A B7 BA 2B A3 1E 1D 1A 07 DB 64 A9 54 41 20
 23 E0 7A 57 9C DF B0 DA 79 D0 E6 56 9F 0B 21 3A
 E9 A7 90 BC 3E E8 59 36 F6 43 89 7E 2A BF 5B 7A
 DC FB 4B 61 D9 F4 6A BB 5A 1D E7 C9 84 A9 98 1A
 2E 49 FB 78 0C 16 92 1E 6E 51 09 63 30 D3 E6 5C
 FD BE A8 B4 A9 48 19 89 CD BF 4C A1 F0 3B B8 FC
 D1 1D 0E A7 11 DC 3E 8F 0C 18 F3 2A 68 5E 90 D9
 03 E8 EE FB 2B B9 46 A5 C0 92 5D 7F 1B 3D 01 9A
 BB 45 41 7F EA E6 B2 1F E0 AB AD 24 93 63 2B BB
 C4 AA 21 E5 89 80 0D B4 89 25 EE F4 9E FF 5F FC
 60 29 84 03 20 D9 60 B4 17 79 A6 55 0C 5B 67 F2
 4E A4 6E 4F 96 F5 5F 19 1F 26 B5 59 D5 79 30 F9
 9C 51 67 9C AE DD F9 EF 1B 88 F1 FA 83 13 BA 0B
 A4 F4 22 65 2F 03 56 62 D4 A5 CF 11 A6 38 D7 4C
 5D 5A CC 60 41 46 F8 5F 70 C7 AE 09 3C F3 0D FA
 33 8F 31 6C 12 CF F9 EE E6 6F 86 9D FF DD 2E 78
 CD C4 F2 AB F3 87 DB D8 20 77 37 93 8E BA F8 FF
 F2 6B 5C 37 31 D4 D9 81 64 5A BC 7B 68 C8 2E 16
 CA 7E 76 B2 81 B2 AD C1 4F DF 8F E2 70 83 93 11
 D8 3C D5 C2 3D C9 CC DD 11 B1 21 87 51 0E AD 2B
 05 45 D2 3B 82 EC 53 6A 6B EA 68 91 7D 7B 22 21
 CD 63 14 5F A7 FD 9A F6 41 F9 93 C1 15 C2 20 B3
 B4 4F 75 BE D6 45 C4 A9 40 7B 05 A5 47 29 16 96
 F7 96 0D BE 33 B1 D8 B2 84 9A 95 0C 78 4F 16 27
 86 BC 47 A2 BA 33 9F D4 56 7D 66 0B 49 FC EF D1
 E3 49 90 90 36 30 B4 E7 11 49 9C 0A EE CF D3 C9
 ED 63 57 90 BE 1A 9B CF F8 F9 79 30 07 3F 80 B2
 92 10 CB 91 96 30 55 5F EE 48 F4 C5 87 04 8B 45
 65 BE 3E AF 6A BC AE BA 8D 66 90 96 31 F9 D4 BE
 8B C7 2B 55 0C 89 E5 32 B3 A5 69 89 33 34 66 46
 5D 82 37 42 E0 92 43 D3 ED 33 82 14 23 27 51 9A
 0E ED 89 10 EB 4F 18 6E 66 EB 9A 88 FC BE DE B7
 57 9F FF 62 37 0F F2 0A 9B EC B3 97 C6 99 43 6A
 BE C2 43 E3 55 B4 5B E8 AE F9 FD 07 ED 7C 48 D0
 EB DA D0 FE F7 C7 0E 4E CF A6 A3 02 E2 B6 0C CA
 08 89 05 9C F7 A8 C6 75 82 FC 1D 5F 23 52 EA A9
 F3 F5 DA 39 60 91 5F 92 85 44 8F B9 ED 1E 0D 6C
 A7 26 11 AD C6 8D 71 D6 24 FC 3D E6 37 D3 7A 01
 F5 D9 C9 B4 60 6B 5D D4 52 FD 64 76 70 38 DE F0
 E7 CF 9E EE B6 3A 83 35 AC 05 BE E4 E9 23 28 EE
 7B 6B 88 E9 66 5B 6B 81 8A 23 40 10 94 77 6E FB
 E7 E5 A4 CF E1 F0 A2 A5 F5 2D 0E 3C 00 3C 9C D0
 14 47 72 E2 6B EB 11 D6 A2 99 C7 BD 33 70 B3 00
 31 AC 56 BF 51 7B 73 37 92 0A FA E1 36 A2 77 42
 0F 18 28 75 A9 49 DA 42 94 5C BE 73 BB 0B 71 3F
 65 69 F1 B3 75 C7 52 C3 72 47 5F 36 27 A8 DC 97
 B7 C8 5D DD 9F 56 FF 72 C2 08 E7 8B 13 E0 38 EF
 6E FF 45 BC EE 6A 47 FB 67 C6 9B A3 DB 7C 8A CD
 9A D2 9E 42 D2 70 E0 53 3D 5E C2 1C C8 E1 F3 4C
 30 28 FD 99 42 F4 64 A1 E4 4B 63 B6 20 EB 3B 19
 25 15 DC F3 A0 3B 72 D5 75 0E 29 57 35 89 19 7C
 C0 CF 2D F7 44 97 1D 1B D1 85 67 6B B0 7A E7 02
 F5 FD 75 01 24 AA 45 9E 8D 79 62 7B 25 6A 93 E9
 EB 30 8D 3C E8 6F 6A 76 C3 2A 42 72 73 30 D3 E8
 51 08 C8 2A DF F0 1D E9 4F 0D 7C BB C0 1E 37 61
 B7 53 8D E8 5B 36 DB 8D FC 3E 1E 48 7C 45 0E BF
 1D 83 EA BD 68 B7 61 D8 17 58 4E F8 26 9F F1 66
 76 A2 ED 27 5A 1A 45 DE 18 78 FB AF 85 5E 6A 88
 55 AE DB 10 E1 BA 15 52 12 D0 5B AF 0D 31 9E E5
 02 C5 94 3E F2 59 4D 48 1B 77 48 35 87 19 86 AC
 38 51 2D 34 FC 2F 51 F6 68 25 7F DE 5C F1 45 53
 27 7B 93 DE 23 9C 4C E5 11 9C F5 B2 F4 FC F4 B4
 6E 41 B3 A3 F8 78 8C F1 5A 70 6D E7 32 22 92 60
 4D 19 40 48 6F A2 09 5E 4A F5 6F 76 82 BC 9B 8C
 A2 8D D9 5E B5 BB 10 B8 E2 FD BD C6 63 02 4A BE
 31 39 1A 73 2B 54 33 0E 23 D8 1B D5 79 41 29 AC
 2F 56 4F 91 69 1C 1A 16 3D 98 92 66 74 E6 C5 C6
 8D 2A 87 D8 F6 CD 41 7F C8 EC F6 31 07 81 D3 68
 D9 2C 64 5C 99 34 59 F9 E6 E0 E3 95 6C 46 E3 E5
 8C 09 77 85 2D 65 DE 31 6D D6 EC 65 9C A4 3F 48
 54 EE 9B 3A D0 FD CC 47 F9 F5 F0 31 68 E7 E4 C6
 8E 0D BC 23 4B DB 8E 6F 6A 71 A4 D0 E3 BB 7D 53
 92 81 D1 5B 02 9B 48 21 09 97 4A 90 40 DC BA D9
 55 62 52 21 6C 9C E2 FE 91 1C 3C 16 43 20 B7 D4
 23 64 6E BD 49 32 4C FF A9 3F BA 40 6B 12 7A C3
 21 6D 28 2D E2 39 0D 23 9D 96 FA A2 0A 11 CC A5
 D3 4A 2D 80 8A AA 97 48 93 D5 BF 54 97 C0 95 53
 D8 DB BD B3 F3 1D 79 61 22 CE 71 AA 92 D0 43 51
 D5 2D B8 5B 89 B0 22 47 D5 FF E9 A1 12 0D 40 D0
 8F C9 E5 4C 41 67 F5 48 5E 53 65 71 82 C5 4C 13
 62 2D 35 2D D1 73 72 88 54 BB 64 9D 3B DB CC C3
 62 84 F9 F5 39 6B 7A 3E 71 6C 76 6D EF 24 3B AF
 5C 14 51 86 3B D6 1F CE 65 35 D8 F2 3A 06 CB B3
 76 65 EA 28 5C F5 8C 71 72 DD 6C D0 A0 19 29 3B
 09 C5 D5 D1 5F 4A 5D A2 57 82 90 61 BB FA F1 5C
 C1 D1 3E 80 27 FF 1A F2 EC 43 C1 4B D7 DB 48 5D
 D6 E0 97 14 6C 38 CD 83 37 D9 CD 87 BD FA 16 C9
 62 9E E6 7F 7A CA 12 1D 5A 29 30 92 84 47 9C 5B
 13 56 E5 0C 5F BE AE CB 73 4E D9 3D 97 4E 28 12
 C1 60 A5 45 37 22 C1 01 0E 1A 6C 91 2C A1 37 F0
 17 96 66 90 12 27 30 BF A1 18 0E BD 7C 86 3C 50
 B4 B3 3C 2B C8 8C 10 E1 64 32 97 10 6B 8F 98 43
 5E E9 45 D2 2A 01 09 C4 B7 51 83 15 8B F7 C7 8A
 37 B1 E4 E6 96 23 95 45 76 9C B7 2C 03 B0 C7 F5
 13 C4 65 10 8A B9 AF 0E CA 28 9C 87 8F 5C 9D B8
 1F C9 7E 2E 19 5E 1E DD 7C 36 64 10 10 DA 5D 7D
 9C C2 EB BD ED C5 DC 49 49 33 2C ED 04 92 0C C0
 01 62 73 A0 E3 79 6B 21 5C 2B 8E C1 AF AF D1 11
 13 CF 74 C9 6A 42 DC 7A A5 0B 8D 2E 67 52 76 79
 05 69 AF 26 44 22 A3 9A 44 8C 40 9E 4D E2 41 2D
 64 A4 5D 67 9B E5 84 01 97 DA D3 F7 12 56 8A 15
 F1 83 55 D4 BF 32 76 C3 DA 08 DA A8 37 B4 8A 9C
 03 0D 5C 62 FE 2F C9 16 9C C2 86 19 AE 0F 0F F2
 DB 1D F8 F6 A8 5D 89 3A 2A CE CF 9E 92 F5 A7 83
 6D 8C 82 01 A8 5B 5F F4 58 8C A8 8D 4E 80 96 67
 98 D4 F3 A8 88 5E 7A 82 F6 DF 2E B9 13 C5 E2 C9
 2F 41 0F C6 20 A0 3A 76 D8 95 DE 43 8D C8 7B 90
 6B 45 6F E9 D9 58 4B 20 09 4E AA C0 9C 91 36 8A
 B2 CB 8E FD C3 28 8B FD 18 67 AB 06 80 EF B1 C9
 49 E7 93 35 84 8C 71 B5 49 D2 FD 04 A7 A3 D6 22
 73 09 9A 88 7F 90 E5 C7 FB 9F 18 64 38 30 2D 76
 65 E4 C8 A8 D3 CF E4 B4 F1 FD C6 08 68 F1 A6 1B
 A4 E7 A2 36 BF 77 46 DC 52 9A 1C C4 B3 F4 1C 52
 58 8A 7B 85 34 E4 FB BD BF BE 45 FD DB 06 CA C5
 12 1D E7 0E 42 6E 23 96 50 75 DB E7 BA 70 2E 42
 A2 11 E9 22 F8 88 8B 02 2A E7 C6 7A E8 75 02 50
 B8 78 8E D7 A9 A2 C7 51 6C C4 90 7F 4B 03 88 36
 61 26 C0 50 3B 5D 17 05 C6 1A FF 3C 47 C1 F9 50
 3E F9 B5 79 60 D9 86 D5 3B 21 3B 9B 0D B9 FF C2
 25 B0 39 83 C5 75 E1 A8 38 ED 83 C3 D9 01 25 6B
 DC 01 0F 5C B3 21 B5 3E 83 D5 A0 C7 BB E1 3C 8A
 6F AC 8D 69 8B DD E2 15 80 A4 67 15 6C 95 A2 97
 72 39 40 9D D4 4C 81 CB 9C B9 D4 8D 13 60 BD C8
 BD F2 22 DE EE 13 5C FF 3B 0C F0 4A FA C8 1F B9
 F2 D8 F6 D2 E1 46 A0 2E A2 55 02 46 E3 08 8E 3E
 C3 15 10 64 50 26 E5 B1 DD F8 24 93 E2 AE 80 66
 5E 8A 26 F2 52 DC BD F7 B1 AC 44 D4 16 D6 7C 51
 4D 8E E5 E3 C0 38 32 F0 F1 74 DE 91 A0 3A 20 36
 D4 5D D2 EB 18 FC 07 3D 06 CA C1 34 B1 D5 08 1E
 B9 91 68 AA 04 15 66 AB F5 8E 22 91 21 C0 57 81
 34 B8 50 2D 27 F4 64 10 B2 F4 45 2E E2 49 B7 67
 2C D1 B1 D0 6B B4 1D 81 FC 03 92 BE 71 E8 20 24
 42 F8 0C C4 F1 42 AF 49 D8 63 64 10 60 36 C1 22
 16 54 3A D7 CE B3 A6 77 20 A3 BF 73 AF 02 0B 7E
 9F 84 49 E1 B7 D0 82 E5 0A A1 38 9F 7F E9 01 04
 C4 EE 63 C7 46 07 AE 20 C8 CC 97 0A 9E 94 8C D8
 C4 EA 46 F0 37 0C 76 7A 00 81 46 36 0F 4C E4 C9
 9E 0C D7 BD DF 69 18 DB 34 D8 84 1E 01 86 19 CB
 52 BF E0 D7 93 0D 43 59 CD 19 0D AB E3 76 06 93
 62 6F 50 76 D3 78 2D D3 C5 C0 50 D4 D4 13 51 F0
 51 11 F3 A5 4C 78 D7 18 B8 91 AD 7B 53 B6 7A CE
 71 97 92 05 49 FA F6 CA 0D 3E F2 E2 1F A6 48 6A
 77 D2 A6 AA CD F7 18 A2 9C C7 57 AD EB 4B B8 D4
 38 16 40 C6 6C E6 3A E3 FB 93 7C D1 DE 7B 16 89
 16 E4 58 55 2E 27 43 7A 99 88 81 82 2F D2 3A F4
 FA 6D 75 6F D0 CD 8F C4 B1 5B A7 60 49 51 C9 4F
 E2 FC 55 BD 2E A1 46 EC CC 68 35 01 72 48 90 3A
 1D 83 BF 61 93 1D FA 18 AA D2 61 54 EC 17 81 8F
 76 8A CF 5A 2A 17 ED C8 18 55 0D 92 C9 73 E8 70
 38 B8 04 01 42 48 39 FC B6 17 33 39 F7 62 58 CC
 5F 27 F1 D0 EE 09 9A DE 81 11 E2 27 38 5F 7D A2
 1D 1C E1 53 FA 40 ED 27 B2 6C 66 51 17 C5 B6 48
 02 D0 0E 2D C3 DD 06 A7 B8 7D A9 09 FB 99 F2 A0
 51 90 8C 42 BF 99 8F B2 A1 CE 19 27 5D D4 00 40
 13 CE 01 CC 36 46 5D 13 67 5C 65 BB FA 6F 4F 9B
 88 60 39 9D BD C5 0B C9 9D 55 FA B3 76 49 FC E2
 72 6D 95 11 68 B8 43 75 0C 60 C1 5C 45 3A 4C 43
 54 B5 82 88 67 B1 21 7D 30 5F 4E 49 3A 98 B1 E4
 F5 52 DD 1F 9F 53 11 1D CA 75 0C 6A A7 0A 08 AD
 FA 98 47 FA EB D8 E0 92 98 60 2E 46 48 5C C3 D8
 2A 34 3C F5 30 07 62 D7 8D FF 93 0A B9 E9 BB 00
 6B A5 54 34 32 35 97 43 6D 46 50 D2 AD 3B 2F A0
 5E E0 5A 5C 4B 78 68 B3 71 A7 7A B3 1A B2 F9 23
 0A 27 FA 77 DE 05 67 1F 5A C8 B5 68 57 54 DB 7A
 8F 6D 8E 44 49 A7 82 34 CC D0 40 9A 84 62 E7 5E
 2C 06 11 93 0B 4A F9 46 03 13 40 2A D8 BC 2C E1
 60 F1 91 16 D3 5D 8D 8E B6 CB 39 C5 99 DA AA 79
 45 D0 29 02 4A DB 0B 8F 72 6E 69 92 72 52 65 4B
 4B CF 02 E2 96 10 84 A6 EE E4 EF 79 AC 58 CD 97
 37 0D 13 FA C1 A8 5C B9 E2 45 67 96 27 DA E5 56
 27 D1 BC 92 F1 A5 00 2E A3 54 5F 8F 05 B9 E7 EC
 69 05 4F 41 5E E2 14 8B 14 6E 01 02 52 6E 24 76
 7E B7 E9 4C B6 40 37 78 ED 6A 7E BF 1B D4 30 1A
 AA 1E 44 85 05 92 F0 AD D4 2B 2F 67 64 33 32 65
 15 6D 29 A3 B0 04 EC 70 89 A9 DB 31 62 B3 80 5F
 9E 92 EC CD CE 13 BD F5 CB 89 B7 77 25 3F BC 74
 16 2D 5F 4D CA 7D A8 BE 42 0C F1 C5 01 7F 5A A3
 61 CD A5 82 DB 39 6E 31 CB 11 C4 57 D8 18 3B 2B
 9C 28 6F 46 DC 34 87 CE 32 42 0B C8 59 41 8A 55
 73 00 48 7A 9E 4B F4 33 8D 23 9B E0 B5 B0 DD C7
 B0 EF 36 D9 A7 3A DB 2D 79 D4 B3 BF 0F 83 8E 15
 EB F3 AC E5 86 49 D6 71 E9 B5 F7 15 F1 B8 E1 0C
 25 0D 93 9E BE 2C C1 D8 8F 16 84 92 0F 00 56 76
 06 72 37 E3 9C DD 0F 5C 62 B5 ED CB CD 77 D5 71
 56 22 6A 55 87 0A EF 37 13 03 82 F4 13 74 CB 88
 52 46 9F 67 91 D6 AE C3 5D 6B A6 0B 53 54 88 72
 72 7C 75 70 F6 95 7C FE 0F 29 C9 11 F4 0B 53 D4
 BA 44 BF 5F 11 81 9D 48 D5 19 BE 61 5E 8A 88 F6
 69 6E 4D 63 0F AD 77 8C 35 9B EB 6D D2 33 DF 74
 9F 25 C0 44 08 A8 5D 22 C8 98 7C A1 7C 7C 4F C8
 41 17 CF 13 26 55 DF 91 63 D6 D8 3D C6 23 4A 6A
 2C 57 2D C2 4B 52 1C EE 87 F3 32 EF 07 73 C8 53
 0B FB 82 B4 B5 DB 63 70 EE 3D 4F 8F 83 2C 26 44
 FC 43 EC 01 A3 24 E7 5B 31 66 4E 19 CB EA FB BD
 A1 C3 20 D1 05 65 3F 11 BE 34 EF 8D BA EE FE 7F
 24 62 69 B9 1B 82 51 56 4D D7 6D 5F EB 34 B4 8D
 40 78 89 00 54 0A 17 F3 3E FA A1 18 06 B1 E3 39
 F5 F1 18 85 CC 47 35 F4 AF FD EE F2 0C 0B 6A 97
 DC 47 D1 AE F4 BD ED 85 4E 53 0C E2 27 5A 45 6D
 EE BC BF E1 32 1A 7A E2 3F C0 73 A9 93 9A 93 4B
 92 27 42 20 3F F6 91 FB 39 B4 50 AE 31 85 26 84
 B7 0B 45 BD 30 53 3C 3C 76 51 FA 22 AC E8 62 A5
 3F 1A 64 86 8D 1F 65 E3 44 16 96 01 2F 95 9A 9E
 95 CD 88 86 2E AA 6F 40 EE 3C 7A B9 10 05 5E 10
 65 3F 7A 57 B4 25 61 5D 30 F8 E6 B8 A3 0A 91 BC
 EF 14 17 B3 D4 C4 D9 17 BC 84 9A 62 8F 1D 56 D7
 47 F0 13 4C 56 AD 33 E5 B8 2E 55 1E BB 0E D3 9E
 1D 22 F9 F7 33 D3 A5 A8 B1 46 1F 67 ED 24 04 40
 02 E1 81 C1 8D AB 44 B7 A2 57 56 70 59 59 F8 E2
 E8 98 3C BC 1E 2B CA C7 48 A6 7F 78 FA A9 CD 24
 06 60 75 0B 29 8A A6 C7 31 95 5C 2C E3 5F 0F D8
 56 79 EE 85 46 2D 82 1F 41 3E 47 D5 35 21 A1 9D
 3C AF 07 E3 DC 0B 95 79 45 26 9C 55 62 3C 51 13
 19 61 0E C8 94 9F B1 0A B2 0D 9F 1F 4B B9 55 CE
 53 CB EA E2 D9 D8 8A EE 1E BD 8B 5F B5 92 1A 8A
 F3 E0 2A 3C 5F AD C0 0F 06 C7 22 B3 A1 68 A1 6A
 11 1E 66 05 CE 96 FD B9 E5 A9 E7 FD 76 0A 14 E5
 78 C8 80 8F F1 83 D2 50 D0 48 79 7D 62 62 2A 2A
 58 DB AD 10 90 70 C0 67 6E 4E F2 FE A4 4F 38 F3
 41 C0 17 A6 C8 45 F5 0D 77 A4 83 E7 AE 9E 0D 8C
 56 4B F8 60 3A A3 09 9E E0 DC 0F 67 88 F8 8E C3
 78 F4 7B 42 7B 79 D3 1B 38 A7 BE 7C CE E9 75 39
 2A 0F DD EA 02 09 FC AE 02 A9 AB 5A 45 F7 2E 9F
 49 C9 DE E9 75 FF B1 DD 00 B4 45 C2 EE 3C 17 F2
 E0 1A 23 06 7D ED 40 C0 04 96 35 D0 F3 66 53 80
 CF 32 61 41 75 53 0A A6 CA 3E 2F E8 79 B0 4D C9
 75 85 F1 9E F4 70 D6 8A 0F 0A 8C DC 2C A7 B7 EC
 26 2C 43 89 5B 9E B8 C3 28 55 D2 E3 46 55 66 9E
 85 FD E8 78 89 1D 53 52 C3 66 38 AC 86 7B CF 08
 50 34 47 8D 28 9A C3 59 8D 96 96 54 0D 26 4A 5B
 C8 D7 FB 0F 50 E2 78 3C 20 8C 92 91 A3 D8 80 D0
 2B 08 E3 08 09 ED BF AE 88 67 F4 0C 49 8E 15 57
 3C AB 2C 29 47 4F 00 2F EA 97 9C F9 ED 04 18 2F
 9E 5E EA AC E0 42 6C C1 1E 26 8B CE A4 02 CC 57
 5C 00 11 C6 B2 25 16 6B 11 E4 D4 3B F3 BE C9 EB
 EF C8 AF B3 15 57 04 47 85 30 44 24 2D 69 E9 D2
 91 A9 8E 5B 00 84 5A E8 8A 97 2C C0 2B 99 A5 AB
 DC A6 9D 78 91 4B 93 19 76 96 6B AF 14 75 2E A9
 C1 FB 4B 92 D8 D3 CA DC FE 9D 63 BA 17 58 3D AD
 74 8D F0 51 1F 7A 11 9F EA 92 3B 11 1F 9A A5 A1
 EF B8 B1 FB 0E 60 3B 03 F6 2A B2 C2 6D EC 1D 9B
 A1 B0 B0 6E 14 59 49 CA FF AC 1A 91 B2 84 AB A0
 E8 B5 07 FD 86 E9 D9 A4 5D E0 E0 88 90 B6 3C 91
 65 79 21 C0 71 0A 59 7D 21 C2 DE 88 15 40 D1 52
 98 05 38 EE 29 71 57 20 37 36 99 0A 0A B8 69 C3
 1C 86 29 59 81 55 68 BA 66 5F A2 0F D9 6B 72 82
 14 59 CE 48 E7 78 EA 3F FB A7 85 94 AC FF C6 2C
 E0 E9 8F 1D 97 5D 3D C2 95 86 D7 FB 75 0F 37 F1
 E0 D6 CD E8 41 41 EF 53 51 78 C0 CE 3E 5F 99 92
 16 03 A4 08 7C 85 0B F0 C7 F5 07 0E 78 39 09 24
 89 42 77 38 13 DB 4F 3B 48 1D AE A5 DE 32 46 4A
 A4 B1 EF 48 FE 8A E6 C5 A4 58 F2 3A A6 68 C7 E1
 32 D0 41 B0 D2 21 1D 6B DC 84 C6 53 28 BF A3 4F
 C3 8C CE 3A 4F 2F 4E BB 0D 98 75 74 87 DE CC 33
 1E 86 D9 F3 D0 12 31 40 18 B4 7A 7B 43 31 24 85
 CB BE A6 07 A4 9F 7A 74 46 A6 82 04 5F 50 69 45
 86 7F 27 C9 AC D2 C1 07 77 52 8D 28 00 A7 04 0B
 69 10 35 7F E4 7F 33 AF 1C AE 20 84 00 9B 78 D7
 80 2C 88 6C BC 94 AF 02 31 E5 9F F6 CB DE EA A0
 A3 BB 8C DA 56 58 AF 27 AF 24 D0 E4 02 6E 17 71
 11 62 64 3D 2D 50 30 4E 64 E8 5C 0B AC 77 CD 52
 A6 3A 27 06 45 51 22 DA 09 11 BC 0C 72 4C 29 2A
 73 AB 69 F5 43 D7 E1 42 12 49 30 1E E2 3D A2 C8
 2F 27 26 9D 58 41 B1 B5 51 BF 7F 79 29 EF 12 5F
 BB 32 6C 6C 0F 55 96 92 9F AC 13 A6 4F 08 47 EC
 B0 F5 77 24 E3 B1 42 BB D3 EB 16 52 87 D0 68 8B
 E7 7C AB 01 81 55 00 53 C8 EC 8F 88 F6 9C 18 12
 A6 C6 24 F4 19 00 61 7D 2C FE DA A2 23 E0 C5 D8
 E2 FF 5A 99 50 5C 74 19 2E 5A D3 18 FC EE 52 40
 62 CF 5C 4D F2 97 46 C9 03 5B 79 E6 00 DB F5 2C
 04 32 D1 EF C5 53 E5 96 53 AD CE 10 80 A0 F7 F9
 ED 71 E7 C7 FC F1 C7 5D 10 08 FF FC 06 A1 A8 D6
 96 87 BF 18 B4 F7 FD C5 30 86 0E 89 BB 6C FC E1
 B9 FC D1 C2 E9 31 8A 92 3A 39 47 DB E2 E6 A8 56
 A5 9E 82 80 EB 14 72 39 FA EF 3E 2D E8 D8 8A DC
 2A AB 52 56 59 73 8C A8 72 9C E0 90 AA AD 5F 79
 29 73 DF 4C 01 72 A8 3F 64 E7 7C F0 72 A0 6F D9
 9C 11 27 E4 2C E8 78 B6 0E A6 7F 7D 23 2E CE 35
 9B BA 8F 71 7C 0C F0 38 F9 62 64 8F B5 30 EA 51
 06 2A 6D 46 5A 16 03 55 32 4A 9B 79 70 82 62 B2
 03 03 9E 2F 3F F4 59 40 2F 87 01 75 D6 DD 03 FA
 9D 97 08 2A C4 54 D4 39 6F 86 15 08 AB 06 7C 78
 1D CA 32 0F 2B FB 91 D0 BE 6D D5 6B 54 EF 6D 83
 C6 FD 2C BA FF 54 05 19 BB 62 80 41 55 AE 3F C5
 E8 48 C3 D0 9B 43 44 D3 08 ED F5 59 62 00 1A 2B
 B5 C0 E4 7D 9D 69 22 CB F2 93 E7 D9 49 AD 56 F7
 F3 DD 93 28 D8 15 B9 5A 0F 4D 03 C1 BD 78 AC 8F
 C1 FD F8 06 C0 57 CA C5 3C CD 96 BC 53 49 54 CF
 35 B6 1C A9 4E 12 83 B4 87 29 DF A4 0A 68 9D 6E
 9C 30 3D F0 87 E3 87 7D 73 4B 49 BF 2C 66 B1 FD
 98 11 BD 5D 52 94 04 CF C7 39 60 A9 05 79 6B A3
 FC 93 DF C0 3F 69 F2 4B C5 FA CA 23 06 F3 D1 2C
 6E 63 11 88 D0 83 8E 43 13 24 2E 8A 2F 7F 18 1D
 77 3A BD 2F AC FF 32 C3 59 D0 ED 09 91 78 61 AC
 6E 4A 28 73 DE C5 E2 40 04 69 B6 BF 9F 0D AE D8
 62 54 0F 02 E5 E6 F9 02 F9 15 3B 6A 39 6F 38 12
 0B CE 07 F4 80 AC 05 45 6A C0 FC 80 62 BE AA C3
 39 AD FC 15 FA 84 FF 71 2F 29 6A 56 C1 18 2E 3A
 AE E6 4A CB 63 67 CD C5 D7 D3 00 5E 2B 9B F6 5C
 AB F8 51 F7 35 A0 09 E2 24 1C 5C 2B 52 7C C7 3D
 87 D8 3C 9F BB DC 4C 04 7A A6 ED EA 27 EE 67 D7
 6A 3D DF A3 AF 7D 50 2D C2 9C 50 84 74 8D 3A 52
 58 A5 FC E3 98 EA 78 61 31 19 C7 61 91 AE 97 E9
 44 27 84 09 79 91 60 70 94 C0 02 8E 5A 21 98 08
 01 5A 2E BD F8 7D 1F CC AA 42 E3 F8 6D 59 5F E3
 5B B8 F8 D6 E8 C9 86 4E 62 63 40 BC E0 46 3E D4
 F4 90 DB 54 FD 16 36 8D 00 C8 F3 37 24 14 0E 50
 F1 71 03 45 C5 C0 AA 9E 23 16 A5 22 E9 FB 2E 09
 AC EE 27 88 23 BF 34 C9 94 B4 34 C2 A2 56 FE 73
 86 21 90 71 44 9B E9 99 FF 8A C1 3D 53 59 5E 62
 13 68 DC D3 F8 6D F7 D2 67 1A 2D 2E F7 02 9A A0
 F1 21 45 B3 87 6D 4F F3 1C 31 09 A1 A7 71 19 E1
 68 E6 3A 75 27 4F 07 C2 D9 8E E6 29 CF FF AB 37
 B1 AE 22 1B EB 56 06 41 E3 C9 DA 7B F6 2D 83 61
 88 12 A0 FE 8F E3 A6 AB B3 91 AB 15 6D 26 F8 77
 5C 04 EF 50 00 7F EC 3D 3B 90 62 1F B3 19 EC 84
 E9 2F F0 08 E9 61 C7 FF 30 EF C4 48 9F 07 53 20
 6A C6 DB 9F 48 9B BD 90 7D 34 40 EC 58 E7 92 5A
 C0 22 27 FB 1E C2 7E 1B 87 4D 12 49 A0 EB 08 58
 42 A5 F6 39 72 18 52 CC 85 45 86 F0 31 51 A0 99
 12 CD 2F 90 06 6E 73 3F 89 8B 70 FF AD 18 CE 51
 AA B3 E5 A7 D8 82 C5 1C 91 0A 88 4F 10 76 38 77
 CC 57 DA EA 57 A1 FC E9 DC 08 D1 32 55 7B C2 60
 50 0E CA F2 2A 8E F2 44 88 CA 68 19 59 E5 16 1A
 B3 D5 18 81 F0 16 60 59 7C B2 95 CE E0 F1 E7 5B
 7B 25 0C 66 04 4B 9E 25 45 28 A7 38 DD F8 6D A6
 DA 49 1D C1 15 FF 07 E8 FF A9 29 67 92 77 01 43
 08 A2 D2 E3 8B 25 CB 42 66 2B AA F8 22 AD 48 03
 68 FF 55 42 52 E7 E2 90 80 E3 62 6F 1B E1 52 D6
 08 41 A6 DF C1 64 4B 5B 89 25 7E BA 38 73 C8 3C
 AE BE 1E D2 99 D5 28 9A EA 95 F5 A9 96 16 40 43
 93 22 65 A1 0D 4F 23 68 39 94 E4 15 83 CF 1C 6A
 0B AA DC 70 3E 02 E2 0C D9 DE C5 D3 68 AD 27 3E
 0F 5C 45 1F 64 E8 A3 78 F0 7B 4C E6 C6 5A 06 B6
 E6 1E B3 F3 46 2E 2A E7 06 73 5B DC C0 DC DB 3C
 8D BD E5 1F 91 3E AD A9 11 0A BA 4E 5D 6E 60 1F
 AE BF 04 62 67 79 08 AA 4F 6A D6 76 D5 12 63 5A
 16 B8 AC 37 A2 30 DB 6F EB F1 C0 6D 58 4A 16 91
 CB 27 31 74 63 5C 46 63 21 76 FD C3 DB F9 09 BF
 B9 02 88 02 AE F8 10 77 31 61 E2 9D D5 7D 94 F1
 CA 11 E4 A8 58 56 22 9D 8B DB 00 63 E5 FE 05 37
 CB 32 3C 0C C9 0A 9E 9E 75 E1 75 D3 17 98 EF B3
 FB 69 84 3A 03 52 D6 A2 79 1C 19 4A 85 E2 98 A4
 25 92 C6 97 D2 03 13 89 FF 05 B4 0B 32 19 40 FA
 9B 2A 81 60 26 95 50 1B DD D2 BB 95 F7 80 76 CA
 B6 02 46 DB CB 47 44 FE 72 C3 4D 24 FE 7C 97 A1
 DA 7A CA FC 6E FE BE 10 E2 E6 2A 9E B5 10 F1 68
 72 38 B3 8B 8A 28 23 D7 40 C3 6A 9D 62 70 7E D2
 53 BB 8A 98 BB 8E 4B A7 7B 3D AD 2A 48 BE 38 79
 AB 97 2A C3 20 2D 6F 6D 7B FB 55 5C D8 D3 F2 ED
 55 0B 71 35 68 31 8A 6A 02 11 1C 76 05 3A D4 91
 3B A9 FF 3E C8 CC CE 2C BC CB 1D 24 A5 C5 F8 54
 02 4D 94 75 9A FA 20 C0 38 AB FE FC B4 67 BA 7E
 54 02 67 7E 29 6A A0 96 A6 91 EB 8F 61 1F 2E 59
 F3 D2 56 D3 15 23 CA 0B C5 94 75 04 CE BE 16 02
 08 21 A1 E3 36 A7 80 6A 8A 4A 06 A3 8B 4E F9 83
 F0 02 9A 58 83 4B 4F 77 D9 D0 E1 A1 5D F4 62 AF
 2B 59 83 80 A3 11 8F 17 97 C4 C3 76 91 77 33 09
 3D 99 AF EE 2A 10 97 F5 FE 54 48 22 E1 2A FA 23
 3D 39 30 74 79 A6 74 49 24 E9 91 A6 53 E0 A1 45
 EE BE 60 1A 98 52 CB 37 6B BA 0F 71 DD 81 E5 26
 D7 73 EF 74 D3 B6 4D 51 4F 91 C4 9C 9C 6F EF C7
 EC 24 26 72 7F F7 71 99 18 A1 8B 40 4F E5 DE E6
 1F 23 63 F6 80 D0 1D E3 9B 4F 65 B0 C8 F0 8F 92
 FD A6 17 44 4B 21 4E 17 6A 96 60 CA 54 62 B6 8C
 82 60 5B D7 92 CC 0A 8F EA EA 88 B9 0A 84 28 63
 68 67 EC 21 F1 22 E8 C0 75 9B C0 E7 35 E9 62 2E
 B1 0B F1 B6 BB 1B 47 B5 4C 8D 0D B2 0C 9D 31 C1
 94 5E E4 7A 61 00 A8 24 C5 DF 17 BB 05 5E E0 93
 9D 64 4E 9B B2 64 DB 2D 50 17 1A 50 77 59 91 79
 0C 75 8D 14 27 36 0F 19 60 6D 0A B5 23 20 97 53
 9F E8 8D FB 5D 27 5F CD D5 49 5D 6A 1E 02 48 4E
 B5 EA D7 AC 05 47 6C 34 A1 83 02 4E EB C0 5A 9C
 F6 8F 48 B7 A3 98 44 07 EA 87 29 B0 2D 34 25 6C
 24 69 CB EE 6A 94 77 BF 6C CD C6 34 12 BA 50 19
 2B 80 DE E8 B8 44 4F FE AC 4A 8F 29 2A 9E 29 E7
 3A D7 FF 54 18 67 53 CF BF 5E 1C 5E 1A 66 63 75
 01 E6 26 1E B0 70 87 66 F3 62 8E DE 3C C5 B2 32
 0C 7F 1E DF A6 68 5A CF 0F 4D 30 DB C9 72 6C B7
 52 F4 55 18 F6 34 A2 3E 29 F8 A8 33 9E 83 B4 A4
 E9 89 57 DC 0C 1F 29 76 8C 60 E6 7D 5A 68 C9 55
 25 54 7F BC 5F CF B9 90 91 83 2B 12 90 04 F5 E5
 19 E1 D7 6E B0 D6 2C 3A 6F 3C 9E 01 3E 3D F6 F9
 CC 83 1D A0 EE 67 6F 0B 03 0C BD 80 C3 F0 79 60
 13 FA AB 0C BE 9E 73 FB FE B1 62 F0 C7 BA 6D 40
 AD CD 2E E8 23 75 EF ED 21 5D 78 49 63 D0 FB 6E
 AD 15 EA B9 2C 0D F8 7E 68 F0 08 E9 A0 48 B8 6A
 FC 81 A3 6C 1F AC 57 1C 01 38 D6 94 BC 3E 95 F5
 B2 6F B1 4C 7D 26 14 57 ED E9 90 7C 47 21 A0 4C
 FB 10 6C 76 2B 80 29 A2 B7 B9 C4 73 D6 27 AC 1D
 92 24 F6 93 BD FA 15 AA 5D 3D AC 78 D3 39 71 CA
 BC 42 E8 6A DC 01 DB 36 F0 09 2C AE 3D 5E 51 57
 C1 E9 61 18 E6 96 E2 0B 6A 7C F6 A8 00 AE C9 B8
 81 58 F7 1D 6F 9E 74 63 26 F7 50 88 6A 8D 6B EE
 95 17 9E 9C C3 7A 7F 63 3C F5 0C 2F B8 5F AE 2A
 9C 89 96 D2 53 60 9D 6E 7E D6 5B A0 46 BF 40 7F
 F3 07 C4 F5 99 0B 3D 11 BE 10 4E B0 93 F8 1B 7C
 E6 04 EA 0F 1F EE 73 BE 1C C4 2F D3 95 E9 DB 84
 F2 BC 98 0F 3C AA 54 67 86 5F 09 EA 99 A9 58 04
 96 57 F9 E1 B4 1E C0 C0 99 BE 3C 6A 4A 1C EC D6
 4E 8D 7A BE E4 55 EA F6 E9 D2 CF 05 03 FA F4 DF
 0C F6 AA B7 1C 37 4C A1 AE 12 1A 15 7F 94 48 5E
 E3 54 E5 83 FC 23 E3 5B D8 86 47 EE 82 B4 43 8F
 4A 8F 4A C9 1E F7 B2 38 00 8B 2C BA 86 15 9D 38
 12 D0 EF 92 62 D0 2B DE 19 62 D0 AC 24 32 81 C4
 2A B3 C1 3E 83 BA 07 0C B9 D8 E3 56 FF 6B 5D FB
 7C D1 0F CD 59 44 33 B4 9F FC EF C2 D1 C9 36 6D
 BD FA B5 76 41 2F 48 9C D6 33 2E 7F 14 5D BB 3F
 52 A1 11 80 D9 16 99 44 37 80 36 D1 ED 80 54 D2
 52 36 FC 5A 00 06 AE 73 7C BA DB CF 65 79 23 42
 58 75 72 63 D3 0D 98 0D A6 50 7F 19 65 F3 C4 71
 2E 19 E7 76 78 B4 90 75 31 44 6E 3C 40 47 F5 EB
 E5 B1 A1 83 39 1D A1 2A 02 55 F7 6F 59 5A B1 79
 A8 D0 63 1B C3 31 CC 2E B8 A6 48 B1 92 30 17 C3
 21 20 A0 29 96 02 41 89 61 51 97 77 4A 38 7C 62
 90 44 63 00 AE 65 CA F3 E7 31 CB 95 9D 66 59 11
 34 DB 77 7B 98 F0 47 6E EA AC 78 DB 5B 8E 98 1E
 9C 9A B1 01 73 33 55 E1 C2 B6 04 55 D9 45 8F 0C
 47 50 29 29 42 73 7C C2 DE 1A D9 E5 90 E6 00 52
 57 D1 46 DF 68 12 2C DB 81 F3 80 33 FD C3 95 0B
 B6 26 19 2A A0 E1 86 8F 42 42 B5 E7 60 5D 4A C5
 C3 AE 77 50 A8 03 DF 10 36 01 6D 23 C3 5F A8 D0
 BA E8 74 FB 03 03 33 DB 9D 5B 04 AF 85 8F 97 11
 1E AF 71 0C 13 D4 A3 42 8C 7C 3B BE 01 73 A4 E0
 0F 8D 45 B6 FC 9A CE 72 F1 41 8F 20 5E 1D 24 0F
 54 9E 13 CD 12 7E D8 62 11 20 C7 49 E0 6B DF 12
 65 92 85 CA 74 06 C0 B7 AC F9 24 D3 9D FB E4 CE
 B9 2D 1B 94 FF D4 57 5F 11 F3 C5 66 5F 2C F0 E5
 05 7C 87 D0 02 33 27 21 1A C7 A7 43 5E BF CE C0
 87 47 CA 2D 6B 37 40 7E C3 1E BD 23 D0 02 1F B8
 B4 39 A4 12 6A 38 4F 57 45 A9 C3 B0 8C 97 DD E9
 1E C5 85 9F C6 31 27 66 D7 F0 9E 59 9B 77 3E 60
 97 63 D2 61 35 E8 68 BC 47 DA 5D 8F B7 43 95 C6
 26 20 AD 31 17 D0 DE E5 B3 59 40 4A 05 62 4F 52
 2D AF 47 37 FA 45 6A 00 9A 63 AF 87 37 48 B3 46
 DE EF 09 E4 65 B8 45 63 CD 31 81 52 C4 FF BF BB
 2E F1 C2 45 A1 A6 E7 DB 9B D4 8B 1A 11 81 F0 AA
 36 5E 80 61 DE 0C 5D 7A BA A9 E4 58 21 16 1C 3E
 69 CA B2 94 E7 DE 33 69 42 79 34 75 CC 47 6D 61
 49 BD 05 78 F8 E1 C7 CD A2 89 AE 52 CA B2 B2 AB
 84 50 DF 6E 83 70 E4 8A 07 90 E2 7E DB C0 1E 3A
 A8 A1 1E B2 E4 F5 0A 21 28 FD C0 F2 A9 0A DF BB
 3B BB B7 F8 2B D2 AB 4A 25 8E 4D B8 30 AC DC 21
 2B 02 3D 0B 50 65 57 EA B0 23 70 69 A7 12 85 83
 A8 54 35 DD EF F4 B0 DE 3F A2 04 9F 47 9F 80 6A
 77 3E 56 D2 44 D9 2B 73 36 9C E6 DC CA D5 43 79
 E3 B2 FC 65 16 50 D9 95 0F 13 D8 CE F8 97 82 9E
 CF AB 69 56 BC AA 48 D3 47 26 94 5A 33 92 4B 69
 F1 20 1B 3F BF 1F 60 90 9C 60 73 EA 92 54 C6 31
 7C EF 43 C5 A9 B6 E2 5A 73 41 14 9B 54 0C 25 79
 08 F9 47 71 A3 2D 43 FC EE F6 9F 79 6B 63 4B 15
 2F 90 CE C5 CE A1 C2 73 F1 4B 06 80 BC 0B A8 0E
 54 6F C6 16 DF D4 DD 17 3A 49 AC BC 7A 88 CD 99
 1B B6 5E 0F 4A A9 77 08 27 CA 8E 35 E0 CF C6 1E
 82 30 15 1C AE A5 B2 BF AD 08 03 90 E4 C2 6A 67
 44 FE B7 12 BF D2 79 1E D7 4A 51 C0 9C CE A5 73
 8B E4 C7 A5 BC 5A 99 3C 76 A8 78 58 44 34 14 8A
 85 95 75 E2 5E DF B4 B4 CB A4 F5 73 E7 C9 FA 8A
 73 BC 7A 31 C4 C6 5C F7 2B E0 F8 DB 32 61 E1 22
 8D DF AF 17 26 A8 06 91 5A 12 06 12 41 7F B0 37
 E1 A5 15 B6 6C 53 8A B3 47 0F 55 9A EE 98 5A 29
 E8 38 DF 9A B2 80 7F 13 11 1D 62 0F A9 78 5A 12
 A4 68 24 13 5E A9 53 70 9C F5 61 85 AF 3C CC 3F
 51 24 23 80 C2 35 97 01 84 C1 E5 BD 13 D0 1A 82
 46 01 CF F3 6D 8E 1E 12 37 FF ED F9 A0 5E DE 42
 57 24 3B 11 06 CB AD 84 A2 59 97 83 FC F0 35 36
 A5 26 C4 9E 37 39 29 C1 2F D0 B6 82 39 79 8A 73
 58 84 14 7A 84 BE 9A 9B D8 13 E1 5F A2 97 8D BF
 DB 33 A7 D7 C8 4A 17 DF AB BE C5 E6 59 D6 57 DF
 FE 24 6D FC 54 99 B5 84 63 68 FD 51 94 FC 4D 11
 8B CB 9C 18 BC 5E 54 76 C3 52 EC A6 E0 83 3D F7
 69 30 2F 72 8B 67 EC 58 D3 65 1F 1B EC 1B 2F A3
 31 7F 90 E1 6F 7F 62 37 75 EE 21 46 17 53 9C 0C
 E2 2F 40 96 22 5B 25 D3 D0 C2 8F 70 AB 5A F1 FB
 31 DA 9D 2B 65 A8 0A 06 55 26 CA BE 50 2E C9 B9
 EB C2 F3 10 27 6A AB EF 93 B5 4C 30 C6 02 D5 B6
 DF A2 14 62 C3 6E 29 82 5C 70 73 05 1A 44 6C 54
 55 9C 0C 1A 43 C2 F5 30 23 55 58 D2 1B CD BF EB
 77 63 1E A1 25 F5 E9 2F 2C 0A 3A 08 5C 31 5F 52
 2F AA 52 9D 5C AA CC BA 7D 1D 53 ED C8 44 60 4F
 A7 C6 43 0D 64 B5 50 66 2B 6D 92 82 01 B8 9C 3A
 23 D3 43 72 B5 64 37 71 08 E8 92 69 D8 D4 62 D6
 01 F6 74 C5 6F 87 72 8A 25 E9 E3 2A 63 05 B6 BC
 40 CF 8F 6C 12 5C 5A 6F CC 59 CF 94 34 E4 74 36
 A6 FA D2 2F B7 C0 BA 78 18 32 EA 4F 3A 7D E4 0D
 2F 82 58 B2 E0 2A 25 1C 24 DC 2E 1E 42 BA 86 6D
 61 4C 82 DE 47 98 67 D4 EA 21 4B D1 E8 FF FB 53
 95 84 E9 6C CF C9 91 E1 60 DA D5 5B E1 45 0C B3
 B4 E0 E5 8A 1E D9 E8 FE 28 FE 8A 93 8D 6C FC C5
 D1 84 82 B2 99 33 6D 2D 2F D8 7D F9 21 9A DD EF
 C2 70 EF 6A E3 8C 92 18 66 0A B1 04 63 11 F7 1E
 0C C6 29 19 C2 40 42 88 00 38 8C 64 0D A0 79 EB
 91 54 21 92 4C 99 BC 73 8F A4 61 54 8C 9F E5 D5
 3D 5C 95 BB 1F DE 4C EE 02 AC 08 37 2D DF F6 C8
 48 22 BD 07 D6 01 7A 84 20 84 B4 30 B0 8B BB A0
 F9 3E B4 E7 4C 2E A8 D6 D4 2B 2A 44 F3 87 08 BA
 19 25 6E 11 8B 12 75 9F 2A 0F BF 80 40 91 83 FA
 91 43 A8 5C 53 A3 62 80 28 59 86 BE 25 1F A7 2E
 97 13 EE 8F 6D 63 D7 77 2F 9F 51 2F B5 E2 0B BC
 FE A4 37 86 93 90 F0 6A AF 90 E8 8A 9E 41 42 18
 63 67 D4 D2 81 11 D5 D6 B9 61 32 3F 10 06 2A 31
 4A 23 2F C9 75 9F EB 7F 10 2D 76 44 5F B3 7C 29
 E1 42 D8 D6 6A BB AA E3 15 89 25 62 A9 17 C1 E4
 5C C2 15 2B 44 4D B9 FF 56 69 11 36 AA 93 59 18
 3C C9 10 A3 87 18 37 91 0D B6 8A 78 66 6A D8 65
 AD 70 B0 47 73 AF 46 A2 B7 0F BF B2 66 72 D6 E1
 38 55 74 6B EA E8 50 CB 86 30 1B 61 4C F3 4C 64
 54 10 00 E1 C0 18 9F ED DF A2 BE EC 7D 7C 3F CE
 32 BD E4 9E 52 1A F9 16 42 3A 46 F8 8C 4C FB B1
 9A 8F 4F D1 A4 9E 9A 58 12 9A 5F 6E 77 E8 2C E9
 9E 48 0A B5 CE C2 4B 1C 04 F4 AA 92 DD B1 1C 22
 CE EF 67 E9 A5 1B D4 12 6B EC 51 38 2E 36 18 2D
 5C 46 1E 96 EA 59 6A 2C 4D 72 EF 77 65 4E D5 9F
 0C 61 9E 12 93 6D 50 D2 85 39 52 40 FB 27 B0 11
 C4 14 8F 82 0E 27 DD 93 52 6F 3D 8C CC 39 3C D6
 F2 6B 1B 18 9B 88 A4 AD C0 57 8C 88 67 02 CF EF
 F4 58 99 05 5D D9 1A 46 D6 53 81 68 C2 1A AC 84
 C7 5A 7E C6 5E F4 CD 3D D0 D3 F5 EC 29 4A 0E 25
 C8 14 FA E7 55 DB C6 2D 35 A2 E9 CC 5F E7 CF DB
 48 42 CF EB 9E 55 9F A2 A0 E6 B3 4D 90 2A C5 AE
 5A D6 D0 92 F1 F0 BB 50 30 F4 3B 3F 4B 22 14 BA
 07 20 E2 3D 66 E5 CD B0 A2 44 91 DA B9 1B 61 58
 2F 1F 8D F2 9A F6 6D 62 4A 63 07 8B C8 C5 C8 49
 F4 49 82 31 CD 80 A6 C9 1E D8 7D 23 90 72 51 A9
 31 41 88 DE 62 07 9E E9 AD 3F 22 7F 3E 16 CB 9D
 FD 40 B1 D3 10 77 7C 48 DB E5 B4 6C 9F D9 B9 42
 1E 83 B9 DE A6 5E 33 11 F2 91 FD 3A B9 56 3C 38
 6B 7C 13 4E 54 67 AE C7 B8 F6 48 B3 B1 FE 8A B4
 47 3E CC DD 5D C7 04 11 FD 01 BC AA 40 0F 11 52
 AD 8F CB B5 2F BA C4 C5 F7 39 C2 2F FE 05 B1 37
 80 48 5F 0B 36 3F 5C 92 67 F5 69 A4 8F 3F 5E A4
 BA 86 B9 C6 00 B0 C6 A9 68 F2 E6 92 CC F7 7D DE
 9B 06 78 C8 15 11 DF F2 98 A8 01 D2 71 D2 E6 02
 08 17 2C 7D 2E 21 2A F9 2D 81 72 5F 95 A3 13 C7
 81 5B 16 67 9C 16 F7 1F F3 CB 0C A1 0A 17 CA 85
 00 97 D6 D3 85 01 42 19 B1 71 5F 78 5B 3A 7F 0D
 D6 81 A7 75 8A DC 58 F5 02 37 4B 68 2B 4E 8B 43
 22 BE 01 40 8B 43 11 16 C2 C9 00 BC 85 69 43 3B
 FB E4 2F A7 2A CB 4F 1D 01 99 8B D7 91 95 4C 14
 9D 6D C3 FE 6D 2D 23 79 45 85 C8 25 38 27 66 05
 FD B0 E1 FD A2 A6 A3 DA DA DD EF 4C D5 24 0D 07
 78 F9 2A 81 B0 A3 17 23 C8 1F 4E C5 F0 E3 9D 4B
 96 BE F9 B8 57 F2 40 F0 B5 ED 03 12 BC 8A 82 26
 AA 48 3F 63 24 E0 EE 8A 2C FA 6A AC EF 04 D5 3D
 86 5C 38 68 07 83 AB F0 B7 76 AC E1 6E 98 5F 01
 5A 84 C2 68 3B 08 04 AC EB 2C F4 25 C0 FA 51 A0
 7E 78 9C 1F 85 80 A1 31 6D 17 6E 28 11 E7 3C 3F
 90 7D E9 2B 6E B0 E2 C1 8A 08 AC C1 1E 45 AF FB
 2C 49 96 45 C9 C0 FA F0 D8 2A 86 CF BD C3 15 BA
 4E 07 63 D0 9B 96 86 D1 84 CC 54 F1 19 9E 49 17
 3D 79 23 6B CE E3 30 D1 5F 6B 71 33 F9 9F 9D 03
 B4 19 27 14 1F 32 79 1B 54 12 C7 03 CF 84 04 4F
 FE AE A2 90 F9 0D 01 EE 98 7F 3B EB 18 D2 DF F1
 B8 D8 85 9E 6C E8 84 EA 81 28 3C DC E1 08 11 B8
 A5 67 A7 E3 36 03 88 98 09 AB 3D 6F A9 16 61 E4
 EC BC 67 30 84 42 80 35 10 E6 0B 3F 2E FB BA AF
 C5 4E 11 47 4F 56 8E B6 43 4D 60 38 61 B0 21 04
 44 84 7D 18 1B F9 46 96 4D 98 8E 71 5C 68 F1 43
 AB F9 87 B7 E2 48 60 B5 86 E8 6A 34 16 46 C7 B5
 23 F3 56 A4 09 82 2F 7E F8 95 AE 30 97 00 9F 6D
 7D 01 50 9C 6E 56 4A E2 B9 05 23 9C 3A DF C0 BA
 9F 8B FE E7 4C 03 09 CF 9D C2 49 EF DB AD D1 04
 BC C0 77 FB FB 5F E9 F0 8A 10 70 C7 5E E9 0F 03
 23 F3 F9 A3 A0 05 36 20 F1 F3 5D 0C 9C 0C 06 00
 74 8D FE D6 AF E2 CB A3 F7 3B 44 69 DD 29 71 02
 68 70 63 C2 0D 5B 35 17 F2 52 5B F0 60 9B 51 E6
 78 7C AB 79 E3 44 AF AC A0 A7 D1 89 93 77 F2 88
 2B 83 4C 42 AA E2 45 4A DB A3 EB 9C 0A E0 C8 E4
 06 FE FC 1C 6B 78 36 AE 78 9C E9 3B 15 CB 8A 13
 E4 42 5C E2 24 A7 98 29 1B 37 C6 6B 3F 25 FF AC
 4C 57 9C 17 CB C2 D4 77 99 DC 6F D0 A7 1F 93 43
 AA B5 78 37 76 93 46 A9 78 5C DC A4 14 5C 75 CB
 01 69 0A 2E E6 CD 40 1D 5D 5D C8 98 2B 34 26 64
 65 47 14 97 84 B9 A4 25 4F 24 60 39 27 6F C8 53
 B3 CF 22 A4 07 CB C6 D4 F0 06 19 61 C3 01 21 E8
 2A 7A DB 6C F1 57 A5 76 6A 90 6C 84 2C 2E 3C F9
 28 54 C1 BB F9 4C 54 05 95 B0 AC BA 64 19 52 0E
 72 D5 49 39 1F B2 83 1C 35 F3 0F 78 A3 DF 53 76
 D0 78 39 EC 2A 7E 84 5F 2B 2C C4 B2 A7 F1 1B 5D
 86 58 7A B4 74 5D BA 06 0F 19 2B 1D DE EF E0 5D
 A4 87 C4 C7 FA 7F CA 71 26 52 C5 DA 83 7E EC 73
 E2 77 FF BD 6F 64 F3 25 92 D5 26 D9 28 E4 32 B0
 94 BB E3 CC EA 48 F7 92 19 55 87 70 B9 62 F2 66
 9B 56 36 25 CF 02 9C F5 54 60 04 FF 7E 2A C3 6F
 63 84 C3 25 C3 34 6E 9A 6C C6 6E 0C 35 85 11 F4
 74 DD 70 F6 C6 A2 92 58 68 EF A0 74 BB 46 BE 9F
 34 18 9D 04 28 96 1A 45 CC A6 D0 6E 0A 53 2A 0E
 65 72 39 79 D0 67 E0 E4 48 A6 1D C6 C8 E9 F9 18
 EF 07 6E 3D 0C 49 C6 58 1A D3 28 2C AF 70 25 82
 7F 64 F6 4B CE EC 2E EF 5A 66 30 B8 42 6C E6 58
 4B 6A DB F5 B0 5D 04 21 CE 65 DF 47 21 63 18 9E
 C5 2E C5 7A 9D CD 29 A6 17 2C 48 29 C7 63 AA 3A
 BB 79 BF 5C 29 B3 E4 F7 E1 47 93 F5 7A D8 8C 76
 28 EE FE 96 27 49 8F F5 1D 3E 6D C2 6C D1 6B F9
 74 49 FE 21 7A BF F5 85 C8 26 A9 94 F0 6A F8 2A
 DA A3 A1 A0 5F F2 BE 10 66 58 BC 52 C5 42 2D 54
 14 27 42 A8 71 5A 42 FE 17 A4 C1 14 46 A4 69 8D
 26 3B 79 5A 62 93 82 32 12 CE 8B A7 CA E5 96 1C
 81 B9 D6 DD F8 90 CB E5 C2 0C 1B C0 D9 9E FA 61
 8F 2A EA 0A 84 D8 D9 21 C1 5D 9B 6A 0A E7 8B A9
 54 F4 56 19 F9 C1 B9 C9 92 6E D5 8A 9D B1 01 D5
 0C B4 2C FE B1 EA 66 C5 35 64 A4 39 33 39 B6 0A
 3E 61 7F 6F 65 F2 07 85 2F 8B 3D D2 6F 94 49 3A
 DF D7 E9 22 44 CE 93 0F C7 0D 67 4A EA 11 30 7C
 77 F6 72 01 FD 31 35 6E 41 C5 9E 39 D7 6E 92 AC
 29 C2 EA F5 24 F6 69 8E 96 B9 15 D7 0E CF DD D8
 E4 39 6D A6 42 47 44 C1 F1 BA 65 ED 23 FA F1 5A
 8F FF 57 60 29 E0 C6 33 0B 75 87 9A 5C 15 CF 2A
 63 01 CD D1 83 C4 51 0E EA A4 50 DD DA 23 6A 48
 B0 A6 D1 64 06 3F 55 8A 16 4C 66 25 81 DE 47 38
 5B 04 08 B4 0E CA 1D 86 7D 6D 36 31 25 CE 4F DC
 D8 75 73 DC 29 DC B4 E4 63 A6 2B CA 72 4A 4F 2F
 43 4F B0 B2 E6 15 16 7C 59 E2 46 BA 5F 05 61 53
 CD A8 D8 73 3D 88 96 DA 59 C6 BA BE 99 95 D6 61
 66 DB 6B 2B 1C D3 E4 BC F2 59 B0 75 5C F3 90 D7
 EA 5D 12 E8 82 B7 68 EA E3 EF 58 6E 40 DA 89 5D
 53 7C 47 EE 47 19 AB B3 20 25 23 AA 8E 2F 53 53
 63 9C 0D D6 A6 F9 0C 6B A0 6A D3 9A EB F4 05 A3
 DB E1 DB C2 FF D1 6D CD 46 A6 66 87 1C C6 C8 81
 7D 7B CA 95 3C 20 A4 08 60 5E 6A 95 B4 D1 E3 23
 83 04 BC 16 F7 81 E5 EC 37 70 4B 16 06 2F 4B 81
 B4 A5 5D 54 4A 64 5E 47 2E 51 3C 21 B7 19 F2 F7
 FC 0C 44 AA FC 27 66 51 B8 D2 08 78 A9 AB DD 64
 5B 5E 06 EF 04 A4 E4 21 25 17 E2 7A 25 1C 41 64
 AE 51 75 A9 7A BA 07 FB BF 28 FD E6 64 FE 9F 8F
 CD 29 EF 36 03 F6 4D EA 3E E3 15 DD 39 9F D9 8C
 24 D5 A7 27 D8 0D 1A 6B DD 92 96 B5 1B 82 BA E6
 9F 6E 61 83 CA A6 06 50 DA 80 CF 10 7E 91 AD 7D
 54 15 3C 58 1B C3 F5 AC 71 F6 F7 6A 46 F9 F2 1C
 FA BA C9 E9 02 CB 26 AD 4B 28 10 DF CF C9 7D 39
 B6 23 A5 E3 0C 11 07 2C 57 86 0B 5E BA AE 7F 52
 A4 F8 59 6B E2 50 86 25 E2 57 97 F7 A6 86 69 70
 14 52 65 B2 1E 96 68 4C 1F A4 D1 B6 F5 D3 ED E5
 A9 AF FA E8 73 F7 24 6F 89 BD A1 01 3B 2B A7 0C
 21 A1 FD 03 E3 47 EA 2A 4B F4 CE DA 06 E8 27 A8
 66 5D 5B 78 44 D0 B7 49 04 DC 21 54 03 3D AA 5E
 8F F4 6F 85 F7 E3 E3 F3 24 D7 D2 07 EC 12 29 29
 15 DC 93 80 D2 2D CA D2 44 1D DE D2 AB F2 8E F9
 4D 10 60 FD D4 A1 3D 62 C1 00 AF 46 0A 92 1C 28
 B3 0E 72 59 5A C0 0E 4B D8 33 2B 48 16 5E E3 88
 0D A5 B1 2C 28 E6 4C 80 0D 60 44 BF 28 B3 C1 7C
 71 3D CB C8 26 FB 46 76 27 59 33 D2 9B C8 F8 23
 27 5B 0B 48 01 27 FA 24 5B 16 C7 A8 28 BB 02 1C
 08 30 39 64 2A A8 02 0F 0A 4D 37 46 B3 EB DF AB
 7C 20 4B 95 E0 91 D1 67 05 69 4A 12 A0 34 38 7F
 46 68 03 22 BB 40 64 74 A4 66 73 08 7E 4B 42 EB
 72 5B 17 B8 50 86 40 B9 15 C2 40 D2 A6 67 6C FB
 2B B1 A0 31 18 A7 F1 2A F0 FD 1E AB E1 56 B1 F3
 DC 5C 55 5B 56 D7 07 13 31 A6 84 F9 36 A5 9E 72
 09 31 05 19 45 CF 9C C0 27 37 29 8E 5D 34 05 39
 A0 BB 75 22 F0 90 36 26 5C 89 E3 F5 85 87 22 07
 5F 2B 57 E9 FB 2A 01 D4 CA 2F 1A 4E FC C2 85 A5
 DF F9 6A D5 00 F8 74 A9 0E B6 AB F2 E3 7F 06 CC
 44 58 AB F6 3D 63 C7 0F 99 63 0F 01 1D DE 84 BD
 63 60 19 12 53 7D B7 4B 4D 56 C9 0D 15 C3 97 AB
 1A CE C4 BD F0 9E 72 80 BB 5B 21 DC E3 33 6B 7C
 2C 85 40 99 4B 93 A0 3D 02 89 AA DC 54 47 33 09
 D5 04 70 0E F3 B5 77 F5 49 C9 61 87 E5 6D 48 DE
 DC 92 AF 35 68 04 6D 6E D7 D6 FC FD 2A 63 52 0F
 A8 AB 05 8A 45 29 5A 77 5B 62 B1 F7 47 E1 1D 50
 B2 70 E2 85 C6 99 88 85 21 54 CF 29 F0 A2 3C B3
 BC A9 AA 8E E6 2F 6D 40 10 48 79 73 1F 0E 70 C9
 76 E4 26 F9 BA 77 7A A1 D5 6F AA 72 5D 12 32 3F
 E5 78 14 CF 32 37 7F 2A EB F9 D4 40 4D 55 8A 98
 59 4F C8 27 23 63 35 20 C9 C3 24 C2 5B 74 BD 29
 53 DE CF 64 19 E6 8F 9B 36 06 D2 DB 00 E9 9A 88
 62 3C EE 81 FC F4 FC FD 9F FA CF 9C 79 54 EE F0
 3E 7E CF 43 BE FF DB DD F6 BC 63 33 1D 35 75 5C
 20 CC 0F E2 C5 30 60 44 09 27 C0 CC 84 F8 FB E5
 57 8F 15 D8 49 2F A0 5B 95 01 E5 63 BF 11 40 C9
 06 1E F7 67 96 8E 90 C5 97 F1 89 9B 8C CE 99 C7
 06 E5 69 CA AB CF FD 4C D6 97 28 0C 7E E0 BF 5F
 21 A5 9B CD 10 67 7B 54 BD 84 7C 0E 81 7F 70 0B
 5C 52 D9 38 66 CF DD 69 EE F2 21 29 AF 6E A5 57
 10 31 86 6B 05 9A A9 BD A8 BB 8E 6A 57 DD 73 D1
 7F E4 C2 8C 94 B5 4D F4 58 2C 23 43 D5 6E 97 C2
 64 9C 94 99 C4 7F 00 76 35 D7 F8 30 DD 92 FE E9
 FB 24 02 C8 4A 4B 16 44 C8 90 0F 82 74 A0 92 A2
 65 49 40 5B 0F 39 69 94 26 01 1C 42 3B 11 64 DE
 7A 89 C6 16 C7 0C 89 DF 89 58 8F 31 B0 D0 4F 78
 9B 43 1F 15 77 DA B4 D6 55 FC 35 8C 25 D1 F1 67
 E6 AE 03 ED 1D 85 06 74 3F 9D 32 0B ED ED B2 CF
 6E AC 59 56 E3 AC 96 A8 5D CC 26 E9 DB DC F6 D8
 89 BE 99 30 B6 5D EB 77 9C 4F 11 E7 E1 8F D7 41
 78 B9 81 18 D6 89 26 1F EE 1D 0A E1 58 B2 30 DF
 07 E4 DE E8 99 E0 72 40 B5 63 88 17 87 55 D2 DB
 A1 FE 6B DA 53 45 0E 19 68 15 AD CC 8B 9B A5 ED
 04 74 69 9B 8F 45 C9 4D F6 48 F8 E1 0D DB EC D8
 42 74 CB 0A 18 92 E2 16 13 8F 30 F6 88 CC 61 7F
 97 4D 10 05 A6 99 A8 CC 68 0F AF E3 4D 91 4E 25
 C5 D9 A0 2E AE E6 73 BA 91 4B 3F 7A C1 8A 99 ED
 AD DB 36 E9 A0 80 20 A6 5D 0F C0 23 10 6F A4 C8
 4D 9F B9 D8 78 B6 EB FD 7A 23 31 5A 79 D2 63 B0
 10 7C 59 8D A9 FE 14 EF DD AC BD BD 33 20 E3 37
 1A 9D 79 F9 29 7E 61 DF CA B3 3E 28 13 BF FA CB
 1A 8C 65 96 CE 67 6D D6 EC 49 60 BC F4 34 77 FC
 5C 35 65 20 A9 C2 AA B8 9B 88 41 C1 3B B7 BA 63
 72 AE 0C 09 F8 B0 67 B8 12 64 A9 E2 E4 6B D8 EB
 51 3C 6C E1 73 E7 EF EF 3F F4 D0 A2 D9 5C 29 2C
 A1 CE 4D CE BE 43 13 DE F5 88 A8 BC 00 50 AD 23
 B3 7C A8 E8 16 34 F1 C4 26 C8 B3 B8 16 03 27 F8
 E9 5F AA C2 8F 10 88 76 C2 0E 6B 04 95 44 FA 05
 0B 73 1C 21 AF 35 4B 11 6C BD 10 28 27 2C 7A F4
 46 A6 01 D8 07 D4 CA 42 5B CA 45 AD 70 A5 68 53
 81 CE 61 F8 CD 19 CB C6 B6 B8 E1 A5 63 18 F6 88
 ED 24 B1 E1 3E EF D4 7C CB 3C 39 61 17 64 53 06
 33 68 EC 7D DF 24 1A 76 62 06 5B 66 43 E3 ED DF
 51 EF 54 B9 73 9E 8A 65 4C EB 57 BA C1 6D 31 CC
 AD 82 55 E1 01 9D C4 6D 17 32 3C C5 E7 09 AD 30
 8B 23 F2 1F 14 F9 AE E3 CC 4A 4B 20 E5 71 48 BB
 3F 25 87 04 04 92 90 15 A4 D4 DD B9 F7 E4 12 1A
 B0 98 83 8C 6F 30 04 6E 6A D4 3B 4D 5C 6A BB C5
 09 96 9E 2D 10 E0 EE EB 79 23 86 B4 0F 59 8E F3
 48 58 63 15 35 8B 02 C5 82 5A 89 07 57 C3 0D D4
 87 43 16 16 80 AF B2 CC 06 24 04 EC 38 8E DB 84
 48 44 4C 46 41 ED 83 B3 85 4B 1D 4C 14 A6 56 08
 1B C6 68 DF 50 23 50 A3 8D E7 77 62 19 88 E1 9C
 25 9D 3B 1E 42 83 AB 72 21 CD 9E 0E 53 DA 42 ED
 B9 19 46 94 68 1C BF B9 C7 DA 59 F8 84 7B 5E 7F
 20 FE 8F 9C B0 3D 36 AB 22 9F EE 45 6E 36 B0 48
 38 13 5D 65 5B 58 CC 4C 19 E2 87 FE 0F 26 D1 A9
 3C 07 67 FD 21 B7 31 E1 6A 39 22 4E 41 45 C3 0E
 B2 A1 03 83 A0 06 C6 B9 51 3E BB 7E 04 D3 06 6A
 C6 FA 62 E6 73 1B 91 45 76 1B 83 AB 0B 56 B3 E0
 14 22 66 1C AC A8 51 91 9D 99 6A 33 07 51 B5 D0
 A3 58 86 FF C2 1A C4 4C EF CE 42 DD 2E AB 20 26
 98 80 FD 98 76 AC 20 CE 6C BF 35 07 8E 39 08 9C
 B7 F8 0F 1B 7E AC DA E4 5F C3 5E C4 64 B6 95 34
 D6 A2 FD FE F7 E8 A9 F1 DC A7 46 09 FB 54 59 43
 E4 94 B0 03 19 BC 22 4D 88 D4 8E 2A BC C3 56 63
 02 EF 1A F5 D7 4B 1F E7 3C AC 7E E0 75 76 47 DF
 03 17 9D 5F 0C E9 79 34 6E FF 95 C2 E7 56 4D BE
 ED F3 4C F5 EC B9 CC B6 B0 22 E1 83 62 72 ED 29
 D5 70 9B 74 CA D0 60 96 73 0E B3 A2 67 BD 8A 55
 BD F1 1C 1D B7 39 ED A7 F0 EA CE 94 DA 45 9D 37
 56 CC 58 BC 4E 09 FF E9 D6 42 EA 7D CD 61 8A 97
 1A 60 A0 66 E3 FC 5F C1 E9 13 E8 65 AF 65 C4 99
 8C 20 6F F0 B5 A3 E1 1A 1F EE 98 92 A6 8C 2B D1
 63 B5 AD D8 E6 52 BC 2A FD 44 C8 BD 75 75 0F 02
 41 A7 1A 1C 67 87 73 49 A0 84 CD D1 52 B2 7F 6A
 00 E2 79 23 A3 88 A1 9A 16 88 6A A4 F7 44 74 53
 99 73 FB 23 1F FC A5 23 8C FB 74 78 75 52 B4 18
 56 82 7E A0 32 6B D8 9B 85 83 30 E2 9A EB 17 99
 84 1E 44 1E 06 72 A6 B4 1C 26 9A 48 B9 23 32 FF
 2F 6B 5C A7 A3 3E F7 B8 39 4F 4B E0 99 31 FE 3C
 EB A0 6A 07 C6 6F 28 EB 83 F9 12 29 BC A3 3A 88
 43 0C F3 01 B0 D8 E6 6E 87 E1 43 2B 69 BA 98 46
 D6 6C 1B D7 FD D5 47 38 69 44 97 E4 45 8F 31 C9
 12 40 62 7F 8B EF D0 97 DA B4 55 81 B8 38 6B B2
 C0 F6 24 7B 3D A4 6A DC 73 40 0A E0 DD 24 9B AD
 70 E4 FD 96 C1 5D 4B 33 E6 77 12 E9 24 04 9F 34
 18 78 E1 62 01 28 AB 95 B7 F3 E5 CD 8B AC 66 0B
 32 EE A5 94 C5 21 AD 3B AC ED 90 00 0C 22 43 F7
 01 36 5D E1 AB C2 B9 C4 C5 0A 79 73 AD B5 50 C9
 06 5E F8 64 B0 A5 8A 7A 15 EB 84 E5 B6 57 A9 09
 15 9B 52 A6 DE 71 7A 6B C6 C0 32 61 E9 4F D3 04
 8A 1D F2 3F 23 29 9D 50 9F 93 6C 94 C1 40 90 8C
 22 C6 DD E1 4C B2 2A 78 73 E9 18 93 A2 41 48 E4
 75 89 BA 10 99 7F C8 74 4E D1 AF BA 65 5D 4B B8
 37 0D 9C C4 F7 E0 57 76 D8 D6 CF B9 28 8E 74 00
 D3 AF 8A D5 12 35 FB 95 DE FE D3 93 81 9B 3D 74
 DB 1E 79 F4 68 69 5C 5D F8 50 04 4E 39 F6 71 08
 D9 75 1D AF C4 C9 C3 02 F8 D9 A2 9A B7 B0 40 02
 A7 1B 54 59 9F CE 2B C1 D9 27 5C B8 E8 02 06 CA
 E7 C6 8D 54 42 0F 00 DB E3 00 7F 28 DE 29 4E C6
 CD 19 EA 6D 75 0E 1F 68 9F 5C 03 34 11 EC 3F D2
 17 95 06 E7 8D 48 B5 C1 93 82 9E 61 86 6E 97 44
 81 77 F7 A1 AE 12 64 1D 2D 1A 7C 95 F5 26 B1 FE
 88 0F DF 52 20 84 94 3D 36 5F C7 31 44 87 D8 6F
 17 75 58 2A D5 97 AB 50 FE B3 56 C6 0A C6 11 FB
 EB 02 FA 84 49 84 ED 39 44 85 68 E1 4E D7 FF 18
 2B 61 51 5C BD FB 48 7B 12 6D E8 F0 29 43 90 D1
 E4 80 30 6F A9 64 A2 12 9E 21 88 A5 51 9D 2B AA
 23 C6 D6 57 76 CE C0 0B 6F F2 A9 61 E0 32 51 B7
 94 45 D6 14 05 BD 5F 45 C2 D0 62 F7 8B CC D6 2B
 2E A3 7E 01 29 6E 84 E4 63 43 4A 11 E8 91 7C 45
 FF C5 82 D2 74 82 AA 8F 54 1C C5 A9 05 A4 EE 6D
 D5 3C D1 E5 97 B4 CA 91 EE 35 9E 84 1A 11 09 59
 D2 D9 60 DF 75 F0 DF FE 8F 60 FD EB 52 0C 21 1C
 71 32 70 DE 35 89 22 BC F8 02 30 4A 67 EF FD A7
 58 B8 98 FD F1 51 86 11 C3 8A 72 32 C9 91 C0 05
 70 A0 09 49 A8 31 3E B7 16 EA 24 55 C2 E7 9A 75
 98 FE D3 9A 3B BB 03 6E B2 B7 98 7E 54 17 5B 4E
 4E 26 AA B4 28 05 50 58 4C 57 59 7C EC D4 33 A9
 3D 9E 9C 3B 10 EE 35 DB 5C B5 E0 B5 87 6F 87 00
 B5 0C 3A 3F B3 E1 BD 83 61 98 81 5D A0 D7 84 C1
 D3 40 90 E1 99 D8 3B 5A 37 5B DB 87 95 FB 97 4B
 9A B4 2F F7 44 10 70 E2 83 48 EE 37 A0 8D AE 4E
 27 99 71 E5 60 30 1C 0B 23 12 DA 30 C2 C7 07 9F
 34 9A 57 13 B7 E5 37 20 B6 6E D1 0E CF 99 67 95
 1D 73 E9 9C 7B 82 10 0B DD B7 61 F9 3B B5 A6 06
 4B B3 B0 43 93 19 EB 6B FD B2 6B CF D9 E4 9A 2A
 9A 93 70 99 DC BE 5A 13 57 4A 01 C8 EA D8 C3 7C
 6F 01 79 AA 08 43 E3 AE FB D1 9F B7 01 CD 50 44
 47 0D E7 22 16 3C C0 F3 B5 46 41 B7 70 7D 6D 81
 B4 7C 8D FF 57 4A DD D6 68 EF 65 F0 67 81 94 5C
 C5 9E 87 54 92 BE 27 E3 37 D4 FD FB 0E 77 87 39
 C5 CE 4F 4C 60 72 45 93 75 55 39 52 C9 6F AE F1
 5B FD D1 1C 07 81 AA 84 6E 32 40 AA 14 3C 3E 92
 EC 1C 87 41 7A 17 2B 7C 07 45 CE 76 EC 1D 19 4B
 98 9D C8 E6 52 3C 1C 40 6F 07 AC 94 33 22 33 E9
 ED C5 09 2D 27 BB 47 B4 5F FA F9 F9 60 B3 03 FA
 C4 1C 1D 53 96 28 72 CA 26 79 55 29 E4 76 0D 9C
 AB 2E AD CA 05 65 00 10 60 97 47 C8 61 42 0B BA
 6C 9C 82 8E 1E 16 CA 83 6D B5 EB DA A5 03 6E BF
 5C 3B 34 67 B7 72 67 8D B0 0A 21 AC 88 3F 48 8E
 BB 07 38 20 76 BF AC C0 23 5C 5C D2 FD 1C E0 D7
 53 D9 D0 0C FE 93 00 44 4A 5A 49 88 78 3B B1 5A
 35 20 82 4F 1C 0D 34 EC 13 CF 24 83 AC 95 03 11
 D4 69 7D 35 4F 0E B9 67 99 8F 87 7D 9D 3A 67 11
 C7 B3 CB 29 D9 80 86 AF B2 62 D9 04 F0 EC 73 1C
 E3 64 32 4E 4E B0 2F 28 D0 D8 A3 90 E2 6B 08 4A
 65 83 68 6D 67 F2 AD 1E 0C 90 6A 01 CC 16 72 97
 95 4F 6C FF 50 2F CE 7D 56 CB C8 D1 56 37 A8 8D
 49 89 4F C4 25 34 48 31 4E DC 69 96 83 C0 17 88
 BE B9 D0 DB 9F 29 5A 54 A6 83 6B BB F2 ED 32 74
 FF 98 95 0C 27 AC 54 93 C2 7A DB 22 45 1D 1D F2
 6D 0C 9E 96 12 8F 49 94 A9 C4 13 B4 01 EA 9A 72
 C0 75 EA ED 8E BA B1 2C 01 5E 05 E5 57 1C AA 08
 4F 90 19 36 93 2F 69 B3 29 DA F1 DB 33 D1 A3 C2
 2D EE B3 44 92 AE E7 2E E7 C1 33 19 AE 0C BD A7
 09 CB 7A 4F CE 41 79 BE B0 55 82 AB 87 1C 91 26
 1D 79 C2 3B F6 54 21 A5 C5 1E E1 4A E7 0A 07 79
 A9 CD A5 95 E1 09 23 34 85 5C 10 32 E8 DF 52 CC
 D5 F7 64 E3 82 0F 52 4B E2 A3 EB C6 2D 7D 64 28
 84 4C 3E C8 51 A1 0F 7B 61 48 B2 3A 6E 15 D7 87
 BF 0D 41 62 E2 6A 56 32 4B C6 CA 57 2A 18 48 B8
 3B B1 B8 35 A0 D4 30 66 25 02 82 CB 81 74 2B BD
 5A A1 BE AF F0 0D DF 90 54 BC 2B 31 1E 90 D0 25
 E3 85 E0 6E EB 1A E5 34 DD 1D 6F 09 25 2B 1A 91
 03 D4 55 18 FC 83 72 A4 89 BD 63 8D 66 0D 37 68
 09 55 44 97 A5 F5 F8 CA 7D 9C A2 6F 98 35 32 54
 15 6C 79 6E 50 70 C9 0F 4C 6E 13 CE 1C 24 2F 37
 94 C0 C3 9E 83 16 42 12 F2 D1 26 74 2A 21 44 D9
 36 66 74 63 82 BC 4A BF F8 E9 00 CF 79 32 9D 7D
 7E A3 95 31 6F BB 10 35 67 2B 30 B8 CC 28 75 30
 D9 D1 3C 69 4B 92 EE 56 D3 76 E9 10 8A B7 D7 AD
 6F 27 83 A5 FE F0 70 35 76 FD 3E FD 81 0B 68 2B
 8C C6 A3 14 4F 9D 92 64 B9 7A EE 59 06 69 BC 6D
 E3 6B 54 A6 63 12 6D 37 CC C9 50 BE AA 9F 1C E2
 A6 40 1A 2E 75 13 E4 C4 4D C9 4D D2 91 62 A2 AB
 35 2B 71 2B D3 CA BD 67 D2 6F 90 FA 1F 72 35 B8
 71 C9 BA 5F 9E A2 BF 70 68 41 43 C8 70 24 75 C8
 1B B0 69 E9 AC C9 0C 92 EB 0E 7B 7E 44 71 BC 43
 3F 01 00 93 CC 89 64 D4 98 18 AD D8 AB D3 C0 C9
 23 30 90 15 EB 4F F2 7D C2 8D 68 41 08 1B 5A 4D
 3B 54 D1 5E B5 F1 AC 1D 7B AE E8 E3 1F 9F 8E 31
 EC 9B 1A 22 D1 65 F3 F0 A1 DA 52 AE 25 D2 23 41
 D6 91 1C 0E 85 6F 73 CA 5F 63 A6 EA EF 44 1C FC
 7F 39 E8 22 C6 4B 67 0E 54 16 41 06 E3 48 C9 07
 04 8A A3 31 A2 16 6D CF 3E 0D E3 2B AF FF ED E4
 0D 57 1F 1F 57 05 C9 BA DE CD D2 81 0F D3 AA 05
 A1 CF 84 12 54 87 A6 F5 4F 2E 42 1F 99 FB DE 48
 6B EA A3 16 88 FF 1E 34 CE 44 7C 8A 8F 3F 62 E4
 B7 95 B9 D2 87 C0 09 F1 CC 43 9D 5E 9D F2 70 00
 77 A3 E1 79 E5 8C 7B 09 8F 42 94 8E 0A 7B 69 9B
 4B 4A 30 C5 59 80 B8 BD 4B 8C 95 5A 12 76 EF 24
 13 D0 DC 7C 7B 67 01 BC 1C C2 C0 4C 9A 52 2E 64
 89 1A CC C0 AB DD 46 15 3F 34 3D 4C DE 57 72 60
 2F 59 A1 46 51 CF ED 97 FF 96 51 C7 4E C3 D7 51
 00 17 84 D0 E9 39 51 77 85 6F 77 02 76 26 24 41
 D8 F0 37 48 D6 B4 4B 12 DB 08 9A 43 52 18 3D 59
 C7 E3 DD 30 3D E7 74 1C C8 5E 07 DF 68 61 3F 2C
 C8 C4 C4 EC 5A 87 B2 CB 57 7A E9 E2 4C D1 C6 BA
 AD 9D 87 01 D1 7F 68 89 70 87 9F 26 C2 85 06 0C
 5A 0C 43 3B B4 7D 20 7B 6F 84 43 D7 8B 18 C2 40
 CF C3 A7 09 0D 0D 86 9B DE F0 DF 8E 41 10 4A 57
 C5 2C 0E A4 8C 7B E7 E6 5F 9F 63 51 15 A3 F5 7D
 3A 79 17 71 2A 88 78 B1 2B 50 8B A2 48 79 16 9F
 1F 8F DD C3 38 4C BE 14 E7 1E A5 58 83 64 06 52
 A1 A6 E1 26 25 03 41 3A 85 2A 11 41 5D 52 28 06
 E4 4F BD CA 2C BA FB 1C 26 9A E5 FF F2 C4 72 C8
 61 56 CE E7 0C 2C 46 98 38 42 23 ED 61 B5 5D D0
 72 A4 EE EC CF 23 83 80 01 56 58 4F 74 31 82 4F
 2A 4F 69 37 31 03 C4 CD 50 C1 C2 EE 21 8A 59 C9
 10 41 BB 16 96 57 51 E6 CC 54 31 72 85 07 D5 70
 3A A5 98 23 9E 6E 8B C1 EC 1A 25 CD AC B9 C6 C4
 CE C6 1A 12 0D C1 66 B4 54 94 3D 61 B2 4F 39 01
 95 10 FA 99 7F EC 82 96 E8 F4 6A 66 79 72 6F 74
 FC A0 F8 EC 93 32 C1 F3 48 0E 63 A7 06 FF 8B 6B
 ED 3A 8B F0 BC A5 8F E2 C7 68 FB 85 A1 5D EE D7
 60 CA 93 F7 10 3E 83 13 E1 AE 04 A3 12 C9 9A C6
 CC CE 0D 18 64 72 54 D8 1E A2 2C 3A 00 E1 12 A8
 7D C6 11 DE 1B 58 F3 A1 95 9E BA CA 4B 13 AF D5
 DD 9C 0C F5 47 D2 D1 D2 6E 75 A8 AB F7 49 DD BC
 61 FE 58 2B 6F C7 DC D8 27 3A 5B B4 25 F3 04 29
 29 A7 DB 86 97 08 F6 06 AF 77 1E 5E A0 70 1B F7
 C1 DE F2 59 39 D3 A2 6C F3 84 75 E8 80 3B 0A A7
 2F 0F 0F C3 05 54 87 2C 86 4E 0D E0 D8 2F 89 D4
 AA E0 FF 68 2A 5E 79 07 82 34 8B B9 52 6D 04 E3
 7A 93 B8 2E 5C D2 15 6A 22 58 F5 A6 10 02 FD F0
 88 AA 1E 93 F7 B3 E5 74 C8 2C 8D 0C 14 6C CA 60
 C1 5B A4 2C 7F A2 25 F8 F3 D7 FD CE 7E 4F 2A 8D
 DA CC B0 10 AE 97 9D A2 A8 87 98 AB EA EF 8D 2B
 6F 8C FD F4 76 69 0B 45 B5 AC A0 21 92 BB 50 C0
 21 63 1B EE 75 4B E1 CC C5 7D 3C 33 BD 7D A8 36
 A5 32 C3 7A 0B E7 9F 1E 47 EF E4 5A B6 83 1C 72
 DF FB 5E 5F 77 CD 87 98 D8 58 49 2B 43 00 5A C9
 DB 0D D1 91 15 53 7E 13 61 99 0F 4D 73 70 F6 AC
 A6 31 6F 61 C4 59 E5 07 B1 27 04 9A E2 16 01 7C
 3B 3D 43 F9 C0 77 1E D0 D4 A2 7A C2 F1 C4 1A F6
 F5 2B 41 DE 24 AB 89 90 CE 0D B7 A2 59 57 88 5E
 33 AD 77 75 6D 59 C8 58 E9 60 FC 42 8E 5E C9 2C
 D5 F9 14 5A 4D B7 76 71 71 F4 4A 17 E0 69 AF F7
 22 25 7A F9 51 4C 7E 44 6A 40 78 A9 4D 25 23 51
 D4 2F 67 06 55 11 11 1C F6 87 72 8D E9 37 2E 02
 50 48 05 4D C8 13 67 30 DD 8A 36 EC 39 63 C4 3E
 4F 07 95 EF AE 1E 6F F0 B8 CC F3 FF 01 84 A4 FD
 20 69 CB F3 D3 3E 2A 9A 70 3E 76 DE 71 DD 2B 7A
 68 5F 18 CA 2B 7E 0A 99 58 28 E5 DF 69 35 37 37
 7C D5 9C C3 46 7B 73 85 C1 95 43 BE C0 04 EC 45
 5A 66 06 6C 68 0E 2E 9A 17 E8 27 22 F6 23 47 ED
 22 BA 28 8B C3 2D 26 08 27 60 DC B5 67 E4 F6 87
 9C 4A 14 37 CA ED 09 A7 74 96 BA 34 A7 CB CE 33
 37 2F 78 07 BA E0 71 35 2C 56 12 6C 62 B6 B0 83
 31 8D 1A 79 5D 43 BE FB 96 74 6B 29 ED 90 13 B5
 D2 EF 14 7D 0F 72 BE DB D8 DF C3 99 36 EE AE 6A
 C3 38 3A 44 44 60 92 E3 98 A7 E6 6F 89 7E 79 D6
 CB F2 1A 0B F5 52 58 D8 56 F9 4F E7 8F 9F B2 CC
 FA C0 E5 C7 C2 8D 6F A8 D3 3A 11 F4 D7 D9 9D 23
 51 F6 82 77 8B 08 6B 53 6A 76 AF BF 80 5B 59 95
 7D AE 1E B7 29 F4 38 84 CD 0D BF 71 5E BD DF 90
 BC 1F 47 99 36 79 03 27 DA 15 BA 74 6F 2D C0 3F
 5B 73 34 8B A4 5B 12 EF DF DB 82 C7 9F B8 84 1A
 EC AD 29 5A EE E7 7A 7A D1 AA 7F 9A 82 07 B3 99
 AD AA 6F 86 88 48 59 4F 80 B8 A8 82 B7 4A A2 5D
 38 9E 0C 16 9A 04 E8 3C 12 FB 35 4E 84 47 13 B3
 39 74 1F 0F 9D A5 09 72 09 D3 F3 CD CD 9E 2A 71
 6B 25 59 6D 42 5D E1 CE 25 1F 63 B3 B0 B5 85 55
 D5 45 E3 C3 E2 C2 A9 93 BF 8F F2 D6 22 26 DE 38
 F2 C9 8C 9F 6D 27 D8 A2 A8 A9 21 8A 2B 65 78 DD
 DF DE 26 65 0B E2 84 FF 16 AB F3 A4 7C FB 65 50
 34 C1 33 97 2E 79 31 3D 5C 3A 72 A0 39 31 8D 29
 C4 24 6B 08 26 5A 84 05 F9 24 AE F2 7C 24 D4 ED
 D9 92 7C E5 2D 07 24 F6 2B 11 38 BD 6B E6 5E B6
 95 66 11 36 88 B2 79 57 38 0D 35 41 27 A3 CC E3
 DB 67 AD 8E F9 79 D4 62 90 D5 23 06 C9 F4 9C 37
 5C 9E DF 28 29 A1 E3 F3 A0 AB 99 B9 1B 4C 51 2A
 31 72 E8 A0 52 F2 0F 68 4D 70 C1 CB 30 00 CD AA
 84 F1 AA 34 F1 60 4D 49 0C 5D A5 0D 55 ED 04 06
 BD 29 EF B0 28 A6 3B 2B 8D 47 73 60 D4 E3 7E A4
 02 70 58 3F 32 DE 5E 09 02 57 9E EF B5 5F 46 60
 6E 68 76 84 66 4F 33 36 A4 09 FC 7D 90 05 5A 0C
 BB 90 4E FB 23 E1 85 B4 F3 02 7C 02 A2 31 37 BF
 39 6D 6D 39 68 B8 09 35 C8 6C 55 6D B5 5D C1 1B
 F3 CA FE B7 00 59 6A 45 43 2C 16 3F 46 66 F2 4E
 3D 05 E4 23 71 D1 1E F9 6C A0 2D 13 60 67 C9 FD
 09 A4 5D 89 58 F2 39 BA AF D6 AE 6A FB EC 72 06
 20 CC 3C 66 28 CD 06 01 5C AD 47 54 1F 2E 95 67
 0B 53 61 40 8A 5B 94 12 0A 9C 4F 01 26 79 E7 DA
 00 CE F7 53 CF 1E 00 F1 03 7D 76 BF DB 62 FF CD
 E8 59 D9 9A 81 CA E1 B7 76 5D 6D 3D CF 01 E8 BB
 FD D5 89 07 22 6F 20 66 F2 2E F6 D0 E8 D7 C1 39
 53 D1 78 C3 50 BB 29 8B 47 ED 6D 31 16 51 D5 24
 BE 51 FB 63 66 43 19 89 33 80 5C 3C 81 86 BB EC
 B9 5C 0D 89 2C 2A B9 89 46 FA B6 D8 23 B5 13 CA
 99 13 5E 89 E2 0C 6A A6 A8 DE 5F 8E CA A2 9E 6F
 44 B6 66 FC 26 BC AA 20 E8 27 CA 61 29 1B 93 FB
 4B FE E0 F4 49 9F 3C 45 61 E9 2C 68 C2 DC AA E1
 6A E0 A2 61 E3 FD A0 FC AB DE D7 3A BB 6F 70 9A
 77 75 B2 CF 95 88 14 37 8A 24 55 66 BC 5E 23 1C
 2C F3 90 7A 25 67 9F 5B 45 4C 87 15 38 64 F8 31
 C6 E4 B5 B3 EB 32 A2 9B 08 57 F7 0C 94 A8 39 DC
 D5 D7 D3 06 ED 51 9C 49 3D 2B BB 44 66 AC 3C D1
 D2 D4 D6 E4 B5 8F 8C 6A 20 78 34 C3 13 2A 48 AE
 F5 E6 C8 12 40 3E B7 7E 5B 02 61 B4 E9 1D CF 45
 BE 01 65 66 82 F8 80 DA B4 B7 8B 5D 83 AC 27 A9
 2B 52 E6 09 6D 71 D8 07 94 8F 10 9C 16 D5 BF 04
 FB E4 0D 52 01 F9 96 42 E4 E4 F6 94 4B A7 8F 49
 81 D4 05 2A 6B 58 82 71 F3 DE 81 11 59 F6 D2 99
 15 45 CD 17 41 7E 00 BB 45 12 86 37 53 F3 2B 5E
 39 BB EC 4C 28 EF DE 2D 9D 47 F9 24 4A C8 7C 63
 68 3D 14 1C 94 EC 60 D7 B4 3A AF 55 44 35 85 0B
 B4 D8 74 E1 7F 03 D1 32 03 C6 E8 6C 2F B0 22 7B
 FD 53 88 2D C2 B1 4D 01 42 BB 42 0F 0E A2 ED 77
 1F B4 F1 AD 5D F6 4B AD BE A7 79 3C 40 B6 B8 2A
 BB 46 CD 09 9B F4 C4 D9 E1 80 18 C5 09 5C 67 4B
 E6 21 82 EC 01 C4 3B 2F 66 51 F1 DD 97 87 33 B6
 C3 0D D3 82 DE F1 82 F1 0A F4 9B E9 05 E0 92 F5
 67 E3 0A 65 35 A9 F7 C6 72 B1 ED DD F9 B2 9E E5
 7B 3B C5 95 BF A0 FF D0 83 11 F8 35 52 9F 46 39
 3F 22 CE C4 48 91 8A EB 5B 9C AB 64 DC BD 8D F3
 E7 D9 0D E2 E8 53 9F 79 72 2C 11 69 F6 AF 6C 5D
 6B 55 1D 84 62 A8 A0 63 F7 AE FF 6E A1 E3 9F 62
 B4 18 EB DA 97 45 C0 A6 19 00 AD 4E B0 17 3B 7A
 BE 1A 29 43 41 36 CC E7 AB 92 67 5C 1B 94 D9 12
 B9 7A BA 98 3D 6E 85 74 A8 54 EA 16 E4 EB B3 E4
 3C 73 5C 95 B0 FC AE 36 91 75 E0 12 40 17 27 CB
 09 42 2B 29 67 BD ED 72 E7 EB A6 2E 9E 1C 7D 91
 EA D8 3B 9B FA ED 32 59 70 A6 89 C0 7A C7 73 38
 A9 F6 2E B9 67 76 31 76 AE 21 72 03 32 0B 23 12
 75 1D D3 7A 97 AB E9 C2 0E 12 B9 CD C5 4D 99 A4
 1D C6 8C 43 6C 7B F8 34 1F B8 3E 6C 8A 79 5A 79
 ED 03 F7 C1 42 7F 97 E1 F5 D0 7E 74 1F 14 2A 03
 BC 91 AE 1D F0 25 03 A4 0E F7 74 7C 1A DF 7D 0D
 A0 AD 87 3B 3E 27 1F 5E 5D 0F D4 1B C7 57 FA 50
 79 C2 C8 63 81 6D DD 4D 2C F0 05 5A FB 80 53 BF
 17 CC 01 80 45 DE DC FB 9D 55 4B 8E 56 4B 7A 1E
 7D 60 D9 35 A4 5E 46 B7 3A 0D 16 1E A9 44 78 07
 F9 68 47 65 7A 37 66 A4 1D 02 A2 AC 56 57 CF FF
 70 FB 4E 3F D9 EB C9 6C 20 0C DA 9F E7 18 40 66
 D8 FB 90 F4 A8 23 FA C0 96 AB A3 A4 5A CB 7A D6
 E7 32 22 C3 9A 46 FB BD 2D F9 D3 B5 D8 70 32 70
 E4 59 1C 20 FD EB 63 A4 C4 36 E5 0E F6 39 42 25
 43 D6 B7 A0 EA C8 CC 85 9A 58 20 C8 98 0D A0 9A
 1B 65 81 D8 19 6E 06 99 4F FC 0C 8D C6 CA 78 0D
 0C 90 73 9E 37 3D 98 B9 1A 60 EB C5 00 34 0A 20
 C0 1B B5 BC 76 06 8D D3 C3 85 73 48 78 46 D7 F2
 12 24 9C 02 77 00 68 86 7D F8 F9 58 55 D0 DA A3
 98 E3 75 31 88 A8 1E 98 EC A3 BE 53 EA 73 C2 C8
 B7 B1 36 7E 56 F8 2F BD 9B 9D C6 DD F2 E7 86 04
 9C C3 B5 D5 FC 3D 74 45 71 AE BD F1 0D 21 42 68
 BF 7F CA 87 08 5E A9 8F CD 2F E4 F2 31 53 35 DC
 50 40 65 1A CC 6E 91 E6 C6 55 10 3B 37 FA 96 B3
 E1 C1 16 82 82 E4 82 C5 76 A9 DD A2 1E DB 98 BD
 64 F8 06 AE 34 1F 8D 2B B5 7F 68 BE BD 67 F0 C3
 D7 B7 B0 6D 7A EA 26 F7 99 C2 03 BB E8 DA CB 27
 F0 E9 A9 FA 16 0A 9A 52 28 FE F1 37 07 BE F4 A7
 F2 5C C9 76 93 95 2F EF FF 8B BE 9A D4 95 83 0B
 A4 04 9B ED 00 84 98 FA 46 31 E0 56 D8 0C 9D C5
 45 BC 52 45 C0 E8 2B BA 27 1C 6B AB 96 E0 8E 54
 7B 8A 8E 50 5D 4A 07 E8 BB 08 82 AF 1F 5D 8D B7
 BC FB 84 F0 67 E9 4A F3 57 A2 9A AE 5E 61 70 82
 A9 A6 51 80 E3 AD 24 DC E0 B9 0B 1F E5 EB 3B E6
 C2 20 14 F7 58 35 BF AC 8F 17 94 9E 5D 4E 56 45
 46 D0 2A 02 38 E4 C9 6F 72 9C A4 9E B6 81 77 71
 02 4D 1B F5 2A B4 42 AE DE 2B EF 03 B6 4D BC D1
 49 03 6A DE 9E CC 2E 3E 65 93 C3 1B E8 35 9B 9F
 94 74 AB E3 9F 3B 81 0F A2 4A 22 4B 70 CE EA E6
 64 13 1C 17 C0 C2 2C E8 7D 56 A9 14 1C 09 01 42
 E5 BA 1B 3F 67 85 B6 2B 95 C8 D7 DA 99 0B 3B 80
 2A 26 A5 91 6B CD 9D FA B6 19 80 EC EE 8D FA E4
 38 2E 54 2D 2F B2 B6 AD B5 84 47 4F 3D AA C9 38
 9A D0 00 53 F7 07 82 B2 07 7C 53 3D 68 B7 7E 26
 A9 51 8D 06 05 4C 9F 6A E6 0B D8 8F D3 37 0F 3B
 DB E8 36 43 6E 3B 40 DD 29 71 D8 F9 55 AE E1 48
 7F 05 11 0A 33 76 22 74 DF 51 74 11 5B 57 FD B1
 0D 57 A8 E7 9D 4B EA 73 BC 96 1C F2 28 5C C8 5F
 F1 8D 1D 53 E2 38 B0 E0 B6 71 43 22 33 D7 B6 2A
 FB FD 1E 11 D0 EE 64 31 2D E9 70 D3 89 CC 70 9B
 FF 9F FD 32 A3 A4 B8 A5 A8 8F 73 75 A9 D1 B8 83
 13 E6 DF 09 6C 13 C9 11 F1 51 0E DD 8F 2A 69 C5
 08 5C 5F C3 98 18 84 48 48 A2 E0 16 5B C8 8D 39
 57 AA DB 5E D5 1F 5E 55 63 1F F1 1D 79 43 1D AF
 8D CA BB A3 4F E9 2A 2B 37 CA BF 69 A9 8D B2 38
 22 B7 EF AC E3 F5 D4 14 EC 52 3A DB 9E 82 09 AE
 44 54 C8 2B 1E 45 BD C7 51 41 C4 68 B8 69 07 27
 7B BF 2D 67 06 96 9D DD 8E 72 AA 2B 78 AC 56 90
 42 D0 0D 73 AE 21 6F A6 BB 16 AF AD 52 D4 01 E1
 00 07 44 7C E9 CF D6 B6 0A 0E 93 9D 39 8A A5 60
 1D C3 71 41 C1 04 5B 2D 8D 56 86 13 FC 34 AD 27
 0B 82 D9 C6 CD 29 90 10 09 CC E7 B0 06 2E C3 EE
 07 AF EE 78 BF 1B 07 21 A9 6B 04 12 CD 09 AB 1D
 B7 76 F7 06 77 7D BA D9 28 A8 D9 B4 20 B6 A6 B9
 E6 90 CB 0E 4A FA C0 F8 EB 7A 85 8D 56 FB EA C6
 09 67 DD 92 70 A2 B1 CD 91 43 CD 50 D0 80 B9 11
 81 30 27 5B 25 F6 81 AA B9 18 90 17 7C 05 B9 75
 16 84 16 E0 8F BF 6D ED B3 C7 96 2C 9D 2A BC 74
 37 86 5D 83 DB 68 1F 24 55 3E CC 70 4B F5 9A CC
 51 60 D4 0B D3 BB 20 D9 9C E7 C8 C5 5C BE 82 8C
 CA 53 8F 52 DD 62 AF 9C AA 25 E8 85 22 E3 E7 F5
 1B 86 62 14 54 04 1E D9 C6 CD 59 81 D7 45 37 6F
 07 88 0A 2B AC 46 17 76 13 C6 52 2C 2B A0 62 C3
 6D 15 EF A5 68 1D 4B BB 97 2A EF 01 1D 56 AD 1F
 6A 78 4B A2 C3 47 D1 5A B8 E6 F8 F8 99 A2 2B 7D
 BB 8A E9 0B 22 A9 8B B5 41 0B 0E 24 73 61 68 6E
 E8 05 7A F0 B1 D2 F9 4E 30 36 18 44 5D DF DB 5A
 CE F7 1F 18 E0 7F 48 6C 30 F6 62 3B CF BC 4C 35
 7F DB E4 46 6E 45 53 91 18 4A B0 DC 4D 14 CB 34
 52 41 64 20 7A CC A5 85 50 E2 69 36 84 80 52 56
 E1 6D EF 54 1B FD 08 81 EB 45 E3 98 D9 C2 C6 A0
 BC EC 8E 7A 40 E9 4A 00 74 54 DC DD F2 85 81 C1
 55 2F 59 2C 42 21 19 F9 27 A7 C2 D9 8F 90 BA 1F
 DA 92 5C AA 52 C7 65 80 17 DD 5F 6F C4 FF 37 25
 00 7E 8D 19 AC E7 E5 2C D4 8C C9 C0 C8 EC DF F0
 4F D5 61 13 7C 5F 62 41 22 BC 0E FA 1D 6E 92 8E
 0F FC 68 16 37 64 CF 72 C8 A9 2D D0 DC 9E B3 91
 FB F9 77 2D 47 AD B8 33 E2 5D 37 93 94 1E D5 9A
 F4 FD 22 AD 73 06 AD 2D 04 03 B0 93 8C 15 A9 F5
 28 E7 96 18 38 AE 67 78 DF 4E 24 5D 5B DB 3B 84
 80 C0 8F C3 18 17 63 1A 1D D6 B0 B1 33 EE 23 3A
 0C 10 B0 BC 27 4D 14 9C C0 D1 D2 F0 4D 06 A1 44
 47 56 38 A7 92 C4 81 39 F3 1F C8 A0 FF AC 40 63
 E0 99 3D 31 48 BB 15 4B E2 B4 21 D6 BE 29 7E F9
 F9 C5 52 07 CD C1 5B FC 14 8A 52 2E 05 F9 DC 1A
 CD CB DE F8 5D A8 A2 87 94 28 9E 6F 32 28 63 64
 22 4B FE B3 07 4A 40 A0 EC 2E 62 15 E0 A9 42 19
 8D AB 2F 37 37 F4 0C 79 6E DE 4D C4 C0 7E AF 7C
 7F E5 75 25 51 BE 09 7E 6B B9 82 F6 0B E2 B2 DF
 3E BD 86 DD 8B 8E D4 5B B5 2E 8A 48 BB 2B E8 D7
 EE 74 07 E4 BA 0E B4 E4 39 F2 B7 5B 01 B9 40 50
 FB 9C FD 4A C8 BF A1 BA 16 51 EE 10 C3 1C 88 DD
 2C B3 BA 8A EB 0D 38 8A 9C 8A 88 8B CC 9E 9F A1
 60 6B 32 39 97 6B F3 EF 60 6D B7 11 8C 63 69 85
 A9 D2 17 20 23 14 8C AC E0 62 7E 78 66 5F AA 42
 E1 C5 BE 95 55 60 D8 B5 CC 89 EF 3F CE 5D 9F 1E
 88 A2 AB ED E0 41 80 82 DD D5 61 2F 82 35 6A 93
 7E D2 C2 81 77 07 DC 94 81 C9 1E 16 B6 88 2B C0
 D7 43 BB B4 0B E9 B3 F4 6F A6 4B 20 C8 4A 0D D7
 03 FF A5 03 44 54 F9 E0 33 84 91 25 24 46 B2 06
 CA 47 09 9E 2B 6F 00 37 75 B8 BE 3E CF 11 B5 B8
 B4 9E 32 0C 48 58 2F C0 90 4C 84 EE 00 B1 5E 48
 39 CA 4B 17 49 A1 0D 13 E1 6A C4 9A B6 D0 08 F9
 3C B5 D0 26 5B 9D 85 92 51 E0 A7 82 68 E4 0C 76
 DC 77 27 F7 53 D3 18 8C 85 5B 59 86 B1 91 95 AE
 E0 25 70 AB 2E 5F 20 3F E1 EA 08 EB 3C 64 50 81
 B6 E2 F6 8E 7D 47 E3 A4 A2 2A C6 01 F1 8B 90 32
 C4 DA DB 5C BD F5 55 44 93 96 1A DC 49 97 47 1F
 69 BE 06 DA BF 5E 1D B7 D0 F0 AA D3 4F EA 01 6A
 37 0D 42 E1 A4 57 F3 F8 48 9D DC 72 12 76 1C 82
 C8 97 2A 79 2A E2 B2 00 34 5F C8 64 39 4C A3 6A
 48 24 B4 4E 2C 62 E0 FF 00 5C 2E 96 FA 1A F4 42
 99 A1 7E 16 23 DE 65 D1 66 C9 5B 59 45 D3 48 EA
 8A D3 BE 40 5E 40 9B C1 7C 81 F5 E5 32 05 DA 4C
 BC 5A A2 90 BA 05 1D 86 E4 2C B8 F0 ED 71 E3 66
 BA 1A 01 C7 E5 46 32 99 48 AB 6A 9F 4B A4 C6 D3
 89 AE 0D 12 F8 F8 BF 7D A0 7C A8 7F 24 27 5F 38
 AA C8 19 8E E1 1A 27 12 A8 8F 8F 9B CC 07 CB BD
 69 06 0D 6C 60 D4 C8 FD 00 20 7B BB 47 BD 72 FC
 EF F4 30 CD D1 F5 88 BA 36 88 20 AB 79 76 6D DA
 0C D8 57 B1 1F D6 C6 22 1C 89 40 12 EE 40 37 DF
 F9 42 8B 27 FE 53 69 4F 7A 57 A1 C4 40 0B 2C DD
 2E 5E 80 1D CE EB 0E C8 5D 9C E4 1C C7 BA 40 EA
 CC 94 45 23 2C B1 48 0F 4D D4 C4 A1 2B CF AB 52
 32 21 42 96 42 A8 95 9D 10 4F 93 B5 17 29 A2 DF
 F6 67 4B F6 44 7D F0 7C 67 3C 2F CE 62 FE 33 CF
 C1 22 99 CD 6E 3D 53 72 C5 12 3F 66 72 B4 DF EF
 DB 33 0C 09 54 D5 58 A3 D8 FF 12 18 1E B6 01 30
 AB 8E A5 3C 72 25 C5 2B DD B0 2E 09 8B 8E 9F EE
 66 5E E5 B4 C1 81 9F C4 89 C0 75 54 31 33 59 8C
 66 B7 00 05 4A FB 68 52 9D C7 D7 E1 5F 23 63 A3
 12 99 9C 87 5C 6C 04 C9 0B AF 31 90 F7 36 B7 49
 B2 E6 B9 BE F1 62 49 0B D0 6C 73 02 D0 31 A7 8F
 92 A5 C8 EF 57 89 48 86 2D DB 34 4D C8 23 3A F3
 54 37 3A 7D B7 C6 08 A6 CB D7 53 E7 B9 EF 30 2F
 47 6C B0 76 A3 D1 6F 70 57 B3 E3 37 6B A5 30 F1
 15 47 76 AF 28 B9 E8 6F CD 43 CB 7B 0C A8 B3 0C
 1F BC 13 B5 BE 36 BB 2E D2 67 49 C4 21 56 BD 83
 F1 5A 5F 6F C2 BF 07 BD D1 18 7D DC E7 F6 5F 32
 E4 9F 9A 99 8A 8F BD A1 28 4C 83 7C DC 15 77 69
 7E C1 D5 3A 34 FB 1D 90 AB 30 7A B9 C4 A1 52 8A
 8F BE 13 75 0F 83 05 77 94 3E 66 4A 01 68 3C 34
 18 8B CC 05 A7 B8 83 F2 26 F9 CF FE 29 16 20 91
 46 D7 C3 69 B9 34 ED 11 9E 6C 04 0F 9C F5 78 CC
 DA A1 CF 72 55 ED 47 05 94 E0 18 E8 3E 60 96 74
 57 57 27 35 82 A6 85 E9 6F A0 57 C0 86 D7 62 EC
 B7 63 E5 E6 B4 1B 94 44 F2 8D 65 C0 99 90 CE 12
 82 12 C6 4E 9F 45 06 DD B0 F6 F7 38 37 8E 74 77
 10 4C E6 E6 F9 33 AB 0B FA D7 2C CC F3 66 D7 BF
 F5 46 37 DA DE 7E B7 E4 76 C8 C9 21 8C AB 91 1E
 FE C1 0C 6A 8E 2C B6 59 6E B8 88 03 6F EB 62 35
 46 3B 85 C1 EE 97 FE 30 C1 D4 17 F9 91 D0 0B 74
 BA BB 26 96 A7 57 09 43 B1 C8 A0 91 0F 5A A0 EB
 45 55 2D A4 5A 4D 92 01 73 DB 76 7C 39 7D 9C 77
 25 C6 A3 30 39 88 BE E9 99 6C 04 9A CA 0C D5 41
 24 9D 95 17 75 1F 28 20 2F A6 46 30 F1 5C 00 02
 48 D5 2D 03 A0 CE 0C 65 F6 FD 8B 74 84 0F 07 1E
 77 1C 1E 6D E6 F2 00 93 08 DA 07 EB 5E 93 09 F3
 03 A5 85 4F 60 8D 90 02 55 8F 0F 2E 0F 75 56 74
 A2 43 6D 15 4F 77 FA 51 01 7D 86 75 88 9D A1 B7
 6A 85 9A F2 8B 96 B3 F1 71 0C 34 40 01 F4 ED 13
 E3 70 46 47 84 82 27 7E 76 9B 8C 16 6F DA 1A C5
 F7 DE BF CC 78 F2 E8 8E 66 6D BF 02 B1 45 B6 C7
 DB 6A 21 CF 01 BA 43 96 02 91 7E 8A 00 34 11 A5
 9C 88 56 8B 2A B8 5C FD 98 75 2D 89 68 7B 04 1D
 8A 73 F7 28 7B 95 6C BE 08 FC 9A 29 FC AF 3E C1
 C8 2E E6 37 DB E1 E8 16 B7 A9 18 9E 95 C3 3B 0D
 CB DD 02 87 95 56 43 40 B4 44 79 3B B8 5E 47 E4
 B1 92 FF D3 EA C8 E2 2D 5D 45 C4 6B 8D 0E BB D3
 ED 78 18 79 8F F7 79 CB C7 CE D1 F2 F7 A9 53 36
 67 09 69 32 07 CD A6 30 40 D8 6A 53 AE FE 0C C0
 8C 80 63 F7 77 76 13 43 B1 54 72 20 40 3E 27 4E
 A1 F1 5E D6 43 58 9E 92 49 0A 0F 5A 2D 03 4B B6
 10 E9 15 D5 B3 BD 00 66 E6 C1 1B 54 54 28 37 52
 59 E0 05 06 81 42 A4 C9 F5 98 43 46 2A 0F DE DA
 A1 1B 52 EE D9 D3 8F EA B0 AA EA 27 29 49 24 1F
 37 68 A3 6E 9C 70 C4 C7 16 12 C5 15 7E 8F 79 EC
 9B B1 F3 7C 91 2D FA 1C 2C CC 93 36 6B 63 AA 6C
 A3 07 A6 9A FF C7 98 66 AE 96 2B 83 31 08 9E 11
 39 5E 68 A8 19 09 4A CC 8E 46 E8 26 01 DC 02 E0
 92 0B FE F5 B1 98 D0 D8 75 64 46 48 70 CC 12 3D
 88 56 BA A6 FF 31 A2 FE 2F A4 08 15 4A 75 A1 12
 D5 11 9E 2D 3B 40 D6 8C 35 30 43 D9 DB AB 39 2D
 C5 01 25 E0 BF 57 8C C9 C3 6C 9E 02 90 DE EB 60
 99 E3 7D 59 0B 8D C9 22 96 01 10 CE FB C3 BC 38
 31 61 1E 64 C9 08 ED AD CC FF 0C 35 CE 34 EE 6A
 EA 0C B7 87 A5 C4 43 3C 25 D9 5B BA 9D DE 87 F1
 6A A1 A1 2E BD 17 8E 70 9C EE 56 13 E7 29 1C A2
 37 DC 65 9B 70 3F CF 01 42 79 AC 1C 38 3A C8 E4
 49 CD 96 AF 00 E9 33 2E 31 7D 6E B0 36 86 01 5B
 97 D6 16 3A 4F 9D 7E 04 1F 56 C4 EF 0B 07 70 3C
 B1 D2 85 D8 8C B8 E0 88 3B A8 C2 01 8F 83 98 80
 5F EF 31 3A DF 5F 2D 5C 23 BC 06 0C 48 4D 26 34
 45 C4 F4 6B 90 9D 2C A3 EF 6D 74 44 BC 86 E4 37
 16 6F D0 9B 45 94 CE 6F FC BA 1B 4C A9 54 F1 BF
 13 02 63 52 3C A1 AA 74 A3 57 9E 3B B1 7D CA 44
 BF F0 39 55 77 B5 D0 B7 31 44 E2 A7 97 53 4B 2C
 43 50 3B 95 19 A7 3C C0 53 A3 69 3B C8 FF E5 57
 04 EA ED 0B 2B 48 12 3C 2B 04 EA 09 C3 BA 58 36
 38 3C 93 92 59 36 2D F3 FC A3 E6 3D 58 3E C2 60
 A0 4F D5 BD 6E 17 48 63 8B 17 96 46 10 A8 F2 99
 08 7A BA 68 D4 3B F3 DB AB 50 9D 3C 40 2A F8 C5
 A7 DC 56 F6 22 17 28 CE 08 21 A6 88 84 B5 A9 41
 F8 42 9B DA 40 B6 21 45 06 49 F1 15 84 78 CF 34
 EB 03 34 09 D2 58 71 09 04 84 1A 8D 3F 62 0D BD
 EE 21 B5 6C FD BC D6 42 13 99 CD 8A A8 1B 15 93
 5E 7B 73 67 49 BF 3A C5 CE 48 BB 42 A0 EB 56 C7
 01 9E F8 93 05 7E 6E 4C F4 EA 21 18 C2 F9 8C 4C
 E9 27 51 92 DA B5 41 32 AA 5A A3 5C B8 FE 61 A6
 5F 26 A2 1E C7 66 F1 C2 C9 4E 22 66 37 66 E2 58
 9C 9E 0D 34 AB 4B 21 91 A5 8D 10 27 9C F9 55 E9
 06 A8 7B C7 30 AD 0F 66 0C AF 2E 72 AF A3 F2 79
 CD 7F 4C 1C B3 D1 D2 43 CE 67 92 94 7C 60 DC DE
 9E 8A 6F E1 B7 FB 29 F3 F8 EE 76 1A 9E ED F2 5F
 A3 B9 29 2F 85 9A 48 B4 5E F4 C9 3B 8B 04 89 1A
 90 99 91 25 90 2B FE DF 41 B3 31 B1 AB 10 1E 35
 B0 52 74 BB 1C B3 49 5E 9B F3 61 38 29 89 A5 65
 ED CC 7A 43 57 2D 8C 47 77 6B 6B C2 3E AF 52 90
 94 5C B2 4B FB BE 37 87 F1 E3 01 27 90 80 9E 1A
 EF 1F A9 1A 4C CA 23 0A CA 72 72 47 33 4E B6 FE
 E8 0C 19 9B D1 97 C9 F6 09 98 72 69 18 CE 9F FD
 A1 95 64 77 68 B0 D5 4A E6 45 1B 21 43 B8 67 FA
 87 38 18 55 77 B0 B4 C8 DA DC FF BC 96 75 79 9C
 3D B9 E9 BA 72 75 99 DA 31 F3 47 45 68 2A 79 C1
 F0 1A 5F 53 BA 1E A0 A1 8A 03 6B 59 BC 22 0D 58
 2A B6 44 29 58 2D F6 9D B6 A8 5C BF 0C 8F AA F1
 99 39 F1 E1 F4 B8 31 35 D4 E9 C0 4C 08 AD A1 4A
 21 0D 64 2E 95 CA 4B 56 F4 86 9D 1C 55 7C 44 4D
 9D 34 B4 D1 39 5F 50 A3 8F 02 1B 6A 48 88 DA FC
 35 C9 48 12 B9 D9 18 11 74 0E CC E6 FA 51 6A 4F
 4D 8A 9B 4E D1 7B FA 47 31 45 E5 BC 26 93 F1 43
 A4 19 4C A1 D2 14 C2 BC D9 35 01 77 08 91 10 33
 06 66 98 52 52 CC 2E 1E 4D 22 B4 AB 28 01 3A FC
 E3 66 01 AE 1E 55 F0 C2 96 63 FB 01 7E 92 A1 E1
 9B CD C3 CB 33 B3 2E F6 93 19 B5 06 EB 2B 5D CA
 0B 52 E7 CC F5 3A A9 69 0F 9C 72 0B 45 A0 57 4E
 8F 79 7F 75 A7 2F DB E0 F3 FF 2B 9E 4D D6 99 06
 69 69 7A B0 C3 F5 9B 28 74 ED 3A 8C FA 3D 39 FB
 DE 69 18 96 7C 1A 16 25 08 19 45 5F AC 37 7F FA
 D4 3E F3 69 08 8D F0 92 A9 CF 35 61 BC 16 E8 90
 50 19 24 10 62 91 9F A5 A2 15 A0 60 F8 4A E9 8C
 EE B0 13 58 1C B4 9F 24 70 F3 56 7D 47 43 B4 96
 68 50 91 9C 7E AD B2 6C FC 03 28 F4 F7 32 DB EB
 4A 7B 3E 99 E2 47 DA 39 81 DB BC 28 5F CB 6E FD
 D2 F5 D1 B8 40 DF 78 6E 93 5E F1 51 0B 78 E0 36
 11 F1 3A 29 25 00 80 90 DE EE D4 5E AF 63 4C 9B
 30 EF 46 49 39 62 BC D1 99 F7 E3 AE D0 C6 AE 43
 2C A2 56 18 09 31 91 4F EB 2C D5 6B 19 E2 9B BF
 69 4C 79 3F 7A FA AE 0C 34 AE 44 B2 6B B0 32 75
 00 4C 9B CE D1 81 A3 14 DA 40 96 E1 25 E4 36 AB
 7A 23 9F 2A 1B 73 DA 82 C6 5B 10 D0 56 2A 57 21
 19 C8 5B B9 38 D5 85 00 2C F1 22 A2 25 84 2F BA
 A6 31 BA 8C AC DF B0 CC C5 74 E6 0D 01 E3 2E 5B
 D4 E8 5C 5B FE B6 A2 A7 53 08 86 8F 73 93 A9 C0
 97 1A 1D FA DB BA 13 FC 61 30 9F 30 29 51 0A 54
 93 E7 82 F1 1F DF 06 E6 62 7B 6E 3F 5E 7A 19 1D
 8D 90 2A 1E 6D 65 7D 87 CB 2E 52 4D AF AA C7 FB
 67 D2 23 06 94 CA 68 90 48 4E CE 73 B1 73 E8 9E
 3E 63 DC 62 14 A4 22 61 6D 43 83 FC 97 A3 14 7D
 37 D8 CC 2B B5 2F E9 D8 40 97 E8 F0 C5 96 CC D8
 4C 58 C5 43 10 0B BF 7A 3C AD 6D C4 39 CC E1 64
 5B 5F D6 42 D0 05 CC 35 73 4D 79 53 56 B4 86 9F
 3A AB AE 2E 67 0F 09 B0 F5 F1 86 B7 93 1C 26 67
 15 4D 76 32 0C 75 51 76 FC 54 02 A4 1A 10 9C 91
 EA EC FA C4 07 98 CD E1 21 56 65 3C DB F8 B3 C0
 16 FD F3 0F 30 D3 F0 16 26 B5 CD 78 09 86 11 4E
 44 36 A7 48 C2 A3 53 1A 05 8D 32 CB E7 02 62 60
 3C 2F D1 EC F6 6D 31 7F 6C 4E 00 98 5D FE D5 12
 A1 FC 85 C0 B6 FF 81 FC 95 10 03 05 8E 24 C3 E3
 7E 11 EE 1D AB 15 4E 02 50 83 24 8A 86 FE FF 55
 ED 34 B6 D9 ED E4 1C DE 9C E9 EC AE 8B CB AE B6
 C6 5B 75 48 E8 52 AF B2 6A A5 70 61 9F A0 4B 4F
 23 95 CF 34 4F 5C EE B1 AD EB 69 26 41 23 9A 51
 E7 61 92 1A A4 85 1B 96 65 BF F2 5C 75 DE C6 68
 6F DC 89 33 4B 1C D6 62 84 9F 40 D1 6C 7B CC 55
 7A 08 5E B7 FD 7A A4 D2 91 EB 6D 09 F1 D6 63 B1
 CC 87 7D 1A CB 7C D0 32 F7 63 E3 5D 41 FE 02 45
 DD 8F 16 EC 8B E7 F6 2B 2C 10 79 C9 9F A1 A4 D9
 8F 8F B2 91 06 A9 AA 27 BD 35 46 AE 52 40 C9 74
 43 32 10 D9 64 4B B4 FE E3 E9 8E 96 3D 26 EE 2F
 3B 4F 6A 89 A9 10 B2 A9 51 D2 D4 D7 4E 28 DC 3B
 CF 08 E4 75 0B BC AE CA 29 B9 79 B8 B6 07 92 4B
 EB 28 94 8F 0B B0 F1 34 E7 FA 68 21 F7 8E A9 26
 92 F7 C0 01 35 13 D9 80 97 D6 6A 97 F1 EB 45 09
 F8 D9 B3 86 11 96 60 B1 E1 54 09 CC DB 8D A8 59
 DF D1 E6 6D CD CA 29 A3 08 D5 12 1D 73 1D 6C 16
 C2 AC BA 54 75 2C 4F BA 62 BD D1 15 DB 11 93 02
 C7 2E C3 7E FB AF C9 CB A1 C4 28 57 9A 47 DD 18
 4A 8D 8C 5F 68 54 35 52 FE D7 B0 BF 9A 5C 59 79
 70 E1 E8 0A C2 DC 41 BB 96 3E C0 1D 33 DC FC 1D
 19 F4 6D 4B C9 6B 14 26 D5 46 8B A4 C6 84 AF 11
 75 C3 E9 24 7B B3 9C 65 FE 9A 9D BA AC 48 E5 5E
 8E AE B1 D4 B7 83 F4 31 D3 44 69 31 EE A3 E2 F3
 E2 33 F1 FF 3D EB 86 D4 2F 94 7A B4 69 FE A8 DF
 63 1B 3A B2 BA 13 18 34 0C E7 7D 89 F8 44 E7 A7
 EA 56 92 F9 4B A4 88 BD 98 4B 89 3E 5F AF 6D 83
 0C 80 A7 83 D8 81 2C 0D 9E 23 8F E6 46 F6 39 8A
 DC C4 C0 32 51 47 E1 D8 05 9F 98 46 F5 84 89 4A
 C8 5E 39 68 12 7D 80 FF 5E C5 4A BB 65 84 32 BC
 96 FA DA 20 1B 15 73 F2 F8 85 62 0A 94 AC 9E 6B
 A0 A3 63 8A 1E 89 16 BA 7B 53 A8 18 EB 93 C7 59
 3F 96 BA DA FE 92 5D 60 25 6D 01 8A 7C 8C FF 51
 FC 6E 4D 31 CD 4D DF AC 43 58 85 77 65 63 08 6A
 10 E1 91 BE 61 9A 44 FA F9 76 9D 54 B8 5C E4 51
 A1 2C 6C 08 B3 09 50 7E 1E C2 D1 AD 07 C0 B8 98
 F9 E2 FE 2F 9F AE 30 0F D8 79 9F D5 AA 19 14 D5
 6C BA 40 BA DC 03 80 E5 71 1F F5 14 CA 44 7D E1
 A8 91 13 A9 90 F2 87 C3 A3 5E 97 BB F5 74 0D 51
 85 54 84 26 0A 25 33 52 AB FC 67 29 D6 8F 65 26
 A8 33 BB 5D 76 F0 8D 8C 94 8A 88 9F BF B4 C5 B4
 47 A8 F6 4D 07 A3 72 8C 80 E2 15 D7 5D CE 49 C7
 99 96 CF 36 29 87 90 28 D2 71 89 86 DA B9 3B 41
 D4 5F 21 A4 60 EB 00 23 DA 0E 7D 2D C0 74 E4 40
 BF 2E 12 79 3F A2 E0 EC 3E 79 50 74 35 E0 DA F2
 B4 BA 46 44 25 55 DB 46 0F 11 CA 72 CD 8C 18 EF
 EA 79 75 EF 5D 6F 68 F6 92 B7 F2 E3 1B 10 D1 59
 40 7B 97 DD 31 6D EC 8B BB C9 A6 F5 6D A4 BA E0
 62 A7 7B 80 81 F7 46 DA 98 BF 30 69 DD 5D 19 25
 96 B2 53 78 43 D3 F5 F0 15 9E CA 90 EF FB 8C 6A
 A8 FF A0 14 56 4E 57 1D B6 2D F8 5C BB DA 4B D9
 D4 15 10 C8 05 D7 1D 48 3D B1 A8 4C B6 07 FD E5
 58 68 67 88 DD 8A 25 D1 EB 42 20 57 0D 02 73 20
 BF DE 64 B0 BB 64 E7 C7 11 01 FE CE 8D 73 71 D2
 8C 3B 79 FA CB 7D 5D 10 55 B1 66 D1 37 B9 A5 16
 BF F0 6A 1E ED 3D 73 50 90 D4 E1 24 81 49 91 4B
 9A 8F C2 4A 40 1C 7D BC DB 97 09 6F 41 27 27 EB
 A9 ED 8C 42 9D 5E 96 C1 00 AB 08 C0 8E 93 0B B2
 5D 92 CD 18 EA 63 38 39 8D E2 0D 2F 29 21 88 AD
 1A 46 58 E7 A6 58 DA E1 5F DE 85 28 EA A6 F5 4E
 9E 85 DA FD 12 40 91 C5 E5 B7 3A 1F A2 91 FC 68
 CF 26 11 91 0A DA 48 9D 74 9B A3 E2 76 1B B7 55
 2C 9A FB 01 EE 84 63 DD E9 47 46 8C BA 24 63 DE
 63 63 9F 8F 82 D8 3F 19 17 C7 CF BB FE F7 58 44
 D9 9A 0F A6 4F E0 7B EA 2E C8 50 5F F2 02 E4 E0
 2E C4 21 EC 66 F6 DF 74 2F CC 44 16 7F DA 39 2E
 91 D2 30 D4 5E 86 09 74 25 15 8F C9 CE C2 63 2C
 C3 0A F2 3F 49 C5 BB D5 F5 17 FA 1D 96 D4 2A 58
 DB 41 A1 27 81 DE 54 51 3E BA 44 03 20 C2 AE 82
 E0 5A CA 3A 1C 76 E7 FD 5B 7B 71 AE 9F 5C 2F 9A
 A1 0F 05 7D C2 DF 16 CC 1A EB AF AB 70 2E 40 4B
 83 E8 D3 50 4D 71 2D 77 B1 DE 35 44 35 48 B5 87
 FA 59 30 A8 B2 2B CE 40 2C F3 CA BD C3 6B 98 76
 D7 64 C0 7E 8C B9 FA 84 8C 9B A0 86 5A 00 24 68
 01 1C 52 38 BB 52 43 A0 24 53 AB 55 5E C4 A9 9D
 91 E9 CE 33 B5 87 10 16 3D 1E 92 EE B2 46 93 8B
 A9 58 84 A8 6C 40 4C 29 77 D5 94 8D 63 F5 8B 74
 F7 F1 7C 49 87 97 02 AF 4F 3F 98 83 7B D6 73 0D
 4D C1 CB B0 AC 9D C8 79 ED 9F C0 75 14 F3 E0 E3
 86 98 74 EF A0 31 D4 09 A0 DF 57 96 06 56 0F C9
 2F 8C BD 12 0B 4B 0F 73 E1 DB 96 B5 96 12 72 C9
 1B 68 C2 09 CE ED B4 0C 40 AB 3A 0F B3 67 33 31
 0A 2D 50 C5 42 C1 2F D5 2A ED 20 D1 75 6A DB A6
 5F 39 00 56 21 77 FC 47 F9 29 88 83 0D 20 3B A6
 F8 84 8B 9D 92 8C BA 03 C7 2D EA 28 5E 7C 81 55
 48 45 76 7C AF 6E F6 AC 52 25 5D F1 70 CA 05 DF
 8A 55 83 EC 1F 2D 11 89 32 A7 90 FF 34 37 3E 49
 E3 86 4E CD 6C F8 2F 95 B1 83 8E 65 05 B7 30 EE
 A4 C7 BB 6A 91 BD 38 BF 1C 07 F8 48 99 AD 34 F0
 8C D1 FE 7E 01 15 DD 61 50 0A 5E 84 86 D1 83 10
 54 A7 1B 31 FE E7 8B C3 C7 D8 8A 45 A9 F0 29 E3
 A6 5A F9 68 37 85 29 76 76 DA 39 CF 84 CB 60 75
 6F 3E 49 B7 9F FB A2 84 BE 4B 9A 3E 76 4A C5 A7
 FB C6 12 99 9E 78 6D E9 EF ED 82 D7 5C 41 9D 05
 1E E5 18 1C 1F 1A 4E F2 3D 4F 80 FA 32 EB 6D BC
 90 51 E4 09 17 A4 B4 48 AA 5A E0 1E 8F 22 91 A5
 B3 D8 0A 4E E8 DF 83 33 BA 29 A3 75 62 D5 AA 7A
 E2 56 C6 9C A3 67 CF 61 34 32 8B 81 8B 05 E9 15
 61 83 BF E3 2E 40 D7 6B 68 AC FD 0B B4 1A 70 C7
 CF E3 50 55 6C 4E 73 24 3E 6B 69 08 7E DE 57 82
 E9 7F 60 12 7F BF 19 39 62 CE 76 6B EF 19 57 47
 A2 11 F0 5F 6B 93 C5 12 D9 08 21 60 BF 69 52 C7
 E2 8B 04 4C CF 37 D5 14 0F 95 6F 00 56 AB BA 24
 95 F0 6B A1 BE F9 3F 42 5E ED 07 82 D8 D8 BA 6C
 7F EF 24 7A 6E 1C E9 44 F0 88 82 52 66 CE A2 CF
 A5 35 50 96 F4 A3 D0 17 E7 05 13 45 E7 F4 B4 65
 FE FF E7 94 2C 76 AC 6E DB B9 79 35 AA D1 1F 99
 0E A0 2B 3E 25 9C 53 05 A8 6F 09 56 25 E3 3E 56
 17 B5 F2 93 32 13 3B D4 D2 63 DA 88 DE A0 A5 E8
 01 45 3C 95 85 F5 B6 63 5C 25 E5 D0 32 73 61 EA
 6E DE 35 18 60 25 01 C5 03 E5 77 84 70 7E 51 96
 B9 F8 59 90 C6 2F 17 F5 E0 1B 82 3C 07 A7 6C 0A
 E5 98 70 99 6D 30 71 0D D2 B1 6A 53 32 22 84 41
 F3 62 B0 6D 9D 64 6D D8 6F 46 3D 87 1B 95 98 C3
 19 1A 0D 25 41 C1 B1 65 E4 35 1C 21 98 13 E4 9D
 1D F3 B1 7D 20 34 55 F1 F5 BC 9B 9A FB 7A 6B 8E
 A4 CB D1 9A 3F 3D 79 24 C9 05 7A FC 1D B4 D7 BA
 25 A3 D2 B2 CD 8D CF A4 07 AD C1 F6 C9 A2 36 0A
 56 5D 43 17 C4 4F 2A 01 D7 47 F7 B3 24 78 22 61
 4E 03 C3 62 9D E0 2D 8C A4 92 52 36 0D 3A C0 BF
 BF 40 E8 BE 8C 5C E4 9B 4D 89 A6 95 4B 44 36 7B
 0A 01 E3 40 1C 46 64 9D EF 8B 97 D0 B9 78 A0 F6
 95 9C 64 EB FA 38 01 2A E6 02 69 6F 19 99 F0 AB
 7E 1B 85 8D 01 0B 5D 84 35 6B 6C 4A E2 18 5B FA
 85 1A A8 4A D0 7A 99 C6 B7 21 BF C0 93 23 28 34
 83 65 7E F5 7A CE 78 2D DE 87 CE 72 78 A6 C2 57
 DA 9E 35 63 AA 1F 58 65 B8 28 F8 D7 A8 7F 3B 84
 E7 1A 00 CA 27 AA 7E F4 47 9E 8E CC 26 95 84 69
 07 8A 10 F9 FF B0 50 21 DA 94 51 23 30 5E 94 36
 76 78 7D 5C BC 86 2E EB 3A 1B 14 15 C7 63 B6 D3
 72 8D FD 62 00 89 0E 2A D1 15 41 C2 6D CB 63 4E
 19 43 52 4D D1 83 67 B4 33 0F 9D 36 52 32 AA 9E
 A4 DA F7 D0 58 82 D6 A3 B7 FF EF DF C9 2B 7C EE
 7B 2B DD 82 CB 52 56 68 B9 EF AA C0 FA 75 32 7D
 F5 28 7B 2F 0E F7 A2 AA 56 C3 FD 12 D1 B1 E2 73
 3B 58 55 7A 41 AE 1F C6 19 7B C3 CA 58 9F C8 85
 6C AF CD 84 0C 93 FD 9F E5 17 DF 09 AE A3 0D 47
 69 FF 7C E0 F0 02 5A 17 F2 34 7B 2B E1 8C 2A 42
 9E D0 C3 EE CD 90 63 73 3B ED D2 1C 04 2F 05 02
 79 60 0F 4A 39 D1 88 9B 83 0C 63 48 EA E3 4F 0F
 14 B3 72 EF C9 0D AB 77 45 2D 99 D9 AB 5D AD E4
 FD 15 6E 12 10 50 D2 B4 CE D1 8F 19 80 5C AE D1
 56 96 23 88 84 90 5A 13 47 A6 6E 53 15 BF A7 71
 ED 7C 97 FB CF 6F A6 91 33 D9 67 04 6D 56 D6 4A
 74 DA 99 29 80 31 19 4A 34 23 47 A5 91 6E 60 C0
 E6 F9 27 E3 76 72 C9 9D 3F 5D D5 91 B4 E2 77 CA
 7E D3 90 1E 48 AD 4E AB 72 6D 42 C5 17 E3 8A F2
 AE 68 1D 44 46 D2 49 E0 9C 5B 4B A0 B2 C1 70 D2
 A3 69 EC 37 4C D4 66 1A 48 66 16 9D 7F B3 FA 20
 79 9D 3C FF F2 51 32 3A AD CC 0A 45 BF 0B 33 AB
 46 AE EC 86 15 27 AA 86 91 0B 22 28 A8 A9 E2 A0
 F7 54 CD 56 93 2B C9 C6 AE 18 B0 A5 9A 30 33 74
 39 07 D9 BB 31 38 58 BA 5F AC 37 38 72 17 1D 80
 80 19 C8 3C 37 97 3B 5D 18 2E 40 0F 98 FB 2F 28
 0B 8D 42 63 15 6D 33 3D D7 8D B7 EE 6D 63 82 E7
 9E 0B C9 91 EA 37 59 FE 00 B6 A5 4A B8 60 9A 40
 FC 49 65 FD BB 7C 8F ED 30 94 C4 0F A5 39 C5 8B
 78 39 F9 E7 F6 10 1B 2D 35 5E 9B CE F3 BD 79 09
 BE 88 84 EE 5F 7F 93 51 66 EE C1 8C AC 5E 30 00
 39 37 F4 D0 8E CE 1B 41 16 AC 8E 17 27 2C F5 BE
 B3 EA C1 C9 4E CF DD 44 5D EE AD 00 65 C6 F7 62
 0A A2 D0 90 0B 65 CC 3E F0 13 37 92 25 35 8B F6
 DB D1 41 78 AD 96 BD 7E 8B D7 CB C7 7F F5 AB CC
 29 AF B0 5E F7 9F 2B C1 39 DC D7 1C DF D8 07 7B
 9E 72 A6 7F E8 05 E7 91 F5 34 39 96 0C 71 CB EB
 F0 6B AB FA 9E 21 DA D0 10 86 A9 6A 3E 54 DD 2D
 37 D2 42 1E C4 72 90 04 F5 9C DE 75 A8 A9 FF 0B
 F4 68 1F E0 F7 E1 2D 92 F9 36 DD E4 C4 D8 BC 67
 14 39 99 0F D5 49 9E 35 FC 18 87 FE 76 5A 88 66
 C8 71 6E E9 E3 42 DC 04 E4 9F 08 DC 2A 19 8C 2C
 02 02 85 4D 34 8E D4 7C 1B 31 5D 3C AC 63 0B 69
 49 A6 FB 06 D7 F3 C2 49 55 EC BC 7E 9B 36 E5 8A
 C2 42 2A AA DD C0 2A 2D E5 04 7E 26 FF FB F4 FC
 6F 2B 69 77 11 0F 97 BB F8 66 B5 9D FE 13 EC E8
 FC EA 0D BC F0 EA 4A 51 79 6D CA 06 36 7E 3D 11
 F6 F2 AE 9F DA E4 DF 31 BA 92 D7 FC 91 56 62 4B
 D3 6E 35 EF 28 B2 28 87 74 7F 4D FE FB DD 6E 01
 40 1B 55 13 E6 96 D7 0C F1 DE E9 29 A8 20 26 36
 FE AA F7 B5 D4 66 3F F9 EC 52 2D AF CE 6B 3A 72
 E8 12 DA F2 4D 7B 59 22 45 A8 0D B6 C0 E3 C7 C6
 00 4A B7 6B 51 46 41 FA E9 B2 C1 74 6E 62 33 33
 7D E2 75 D3 71 4B 20 A6 6B 23 C6 79 15 C0 53 C0
 9F 32 94 1A EA 70 BF 58 3A 99 A9 9B 0F 97 9E AD
 92 2C CA 61 4A 98 CB F1 11 F2 E9 F3 17 D4 BA 27
 62 B8 B9 90 20 93 E8 73 A2 86 4B A9 BE 95 66 3A
 FB DB 8E A6 BC A1 75 B2 94 4D E4 49 42 E5 CD 10
 26 7B C1 FC D0 A0 23 B1 6F E6 41 04 64 05 51 4E
 82 51 20 2E 00 FB 72 8F 49 F6 75 99 62 C4 01 9E
 8D 07 59 31 A2 62 D0 96 5A 9C B7 61 FD FB B9 EC
 F9 31 6D 5C 4E 4F 8C C0 67 F0 D7 97 89 D1 3B 72
 EF F6 3E 56 F0 17 0C C3 F1 CA 55 C4 F0 9E E6 A8
 81 94 4F 6C 5E BA D2 66 E2 84 B4 39 8A 42 BC D8
 A0 88 33 F8 DC A7 21 29 A0 23 E8 28 34 62 36 E6
 25 3E 6B 7D FC A9 A2 FC 1D 23 23 45 F8 EF 59 00
 79 3A D3 12 20 ED FF B2 E0 46 84 52 B8 44 76 65
 B3 7E 59 67 E6 AC 36 9B A7 15 BE 3C 80 10 02 00
 F5 26 76 3E B9 2D 05 C9 3C F8 A9 33 4F D2 78 C0
 F5 7E A1 20 F4 6A 40 22 83 EA C5 8E 68 CE 88 95
 88 FD 0D 81 F4 CD C5 D1 5F 1B E5 62 F2 56 7F 55
 53 0B 24 5D 3D 4E C0 9C 40 D9 7A C7 BF EA DF E8
 54 01 41 B7 4A 67 2E CE 11 AE DE 64 76 0F 0A F3
 AF 12 FE 03 24 FE DC 41 BB C2 5A 2D 29 AF 0B 7E
 2C 61 28 CB BB 29 02 74 01 8E 9D 97 03 C0 ED 16
 9D 7C 9D CE 23 F8 26 50 00 C7 78 97 C4 8F 09 38
 98 F4 2E 92 73 6A C0 06 7F 8C 5D 59 56 DE 10 EF
 89 80 C4 4F 73 B0 8B E7 61 26 C6 27 82 44 AF 15
 E7 25 BF AE 3F 2A E8 1A D5 9A 09 4A 36 87 A2 B6
 8D C7 28 44 AA 13 9B 6C FC 06 1D BD 95 7D CF 56
 CA 48 A0 32 6F C0 6D F7 8A 35 3D B6 85 0C 1A FE
 38 E8 48 A3 A8 72 88 30 DB B4 43 00 AE F9 B1 65
 26 50 8A 09 20 CE 37 BD AA 48 C1 8F 9C 5E F8 AB
 CE DF 27 13 09 B9 AF F7 16 CC 72 3C EB EA 2E 6A
 63 CC C5 FF E1 C1 C4 BE 9E 1F FF 5A 72 7E 41 A8
 BD D3 2E 29 72 ED 31 3C CC 1D 3F 3E 1A 70 91 4A
 17 CA D9 45 36 B5 92 7A 5F 1E E9 4C C4 8E CE 5D
 B3 2D C9 65 9B 2A B8 E4 5F 5D 80 3B 23 45 28 14
 C4 3B 77 FB 0C 2F 93 CA 67 52 67 28 42 66 0A 59
 1E F9 21 AA C1 72 30 6F C1 E3 61 4D E0 8E CF 5B
 72 AF 64 2E 58 B4 1D 57 0E 8B 21 D2 B2 B1 C0 80
 D3 3D C8 AF 19 DF 35 EC 98 36 43 4E C6 68 67 4C
 24 86 9F B2 0D 21 39 6A 7F 81 72 FC 40 A6 5F 17
 E0 B8 A9 B6 1B 58 2C BB CE 7E AB 5A 7B DB E1 45
 4E 86 1D A6 92 7C FE 01 DB 1E E4 2A 48 22 18 5E
 96 C6 2E 43 7A 92 BA 3C 74 23 49 E8 3E E6 D9 D1
 67 5B 4B F5 23 D1 DC 3C 14 15 5B 93 FE C6 7E E3
 1D 18 B5 90 2E 79 40 10 28 35 E6 F4 A1 62 34 2C
 0B EE 18 55 E0 E3 1D 2C FF C1 39 31 95 61 E6 DA
 E2 80 E4 22 31 C6 35 1E 80 D5 6D 89 FC C6 D9 CC
 C2 AB AE 4A 91 02 80 EE A1 81 D9 05 CC FF 9B D6
 BC FC 57 B6 99 30 0B 8B 2A 83 00 11 27 9C B2 78
 62 81 72 7C FB 15 5D 55 5C 2B B7 D5 D8 CE 8B 22
 58 AB 60 DB 3C BB 03 F5 65 7D 91 D8 52 84 BF B3
 2D 0F DB 49 D9 17 4A 28 69 D6 AD A8 D5 DF ED 70
 F9 31 E6 BA C2 BB 8E 47 48 0E 86 A4 57 BF 42 CF
 04 18 75 CD C1 27 4A B3 D5 51 CF B4 14 DF 10 F9
 EB 10 58 EB 34 A7 80 F7 E7 BC 2A F9 00 77 CA 17
 A1 AD 51 AB AB 8B 87 9B 60 DD 2A 2A C7 3F CB 2F
 9F 2F 76 F1 5B 0D DA AB EA 34 FC B2 3F BD AC 59
 F9 86 AA 51 80 15 7E 7C 33 6A C7 45 9F 38 EA B7
 63 D1 CF 4D 4D 01 5E CE 76 07 A2 E3 F8 C9 F8 04
 B6 76 07 05 15 19 1F 06 70 AA 11 7D D5 2C 56 23
 D4 79 BE AB CA EB 83 F7 E1 FE 05 16 BB EC 45 42
 F0 57 E6 EC 17 C2 64 96 AE CC E3 63 CE 4D 7C B6
 20 07 46 1C 27 1F 4B B4 39 46 AA C8 E7 BA 78 F1
 DF 84 97 AC FD DD 0C 9D E7 A8 48 12 F5 0D 51 B8
 42 E4 70 98 98 CE 30 2F ED 47 9A 3F EA FE 88 7C
 FC C2 32 95 00 BD 69 F0 38 B9 75 6D 05 C7 EE 24
 8A D7 71 8B 17 37 03 BD 1D 3A 7D 15 72 46 F5 91
 75 E3 62 CD F8 B2 10 F2 70 41 90 4C 58 E0 AB DF
 80 37 A8 C1 DA 4E 44 47 0D F1 B1 A9 5C 3A 40 B4
 0F 4C 1A 2B 02 7F B6 B7 A5 01 C4 4E 05 8C BA 1E
 56 DC 0C 16 8E 7D 78 85 60 20 D9 BE 26 A0 5A C3
 D3 B6 C9 6F CB 2F 6E 23 C1 32 A0 F5 6E BB AC 52
 94 D6 FD 94 18 48 2E FB 26 A4 1B 36 7A 9F CB AD
 4E E1 85 E5 56 1E 11 05 60 E0 BF 34 E1 5F 79 00
 26 5B 14 3B 63 85 EE 30 C3 07 FB 53 0C 9D 1A 61
 3B BE C8 E3 E9 34 24 58 63 FC D8 12 DA B8 DA 29
 4C 4D 76 BE BA 55 6A 51 00 89 CF 0E 3C 35 AD 4F
 EC 5D A5 EB C4 B9 A8 90 5E 59 C4 B1 98 7A 5D C2
 CB BB ED ED 6F 32 88 B5 C4 0F DD 3D 4C 47 6A 88
 90 AB 75 AC 1D 6B E2 24 E4 41 90 F3 D4 B5 B3 ED
 6E A7 E6 CE 9A 3F 10 CA FC 22 68 CF 4C B9 55 53
 73 B3 28 86 66 D8 C6 6E CB F6 41 1F 14 13 BE 77
 82 D8 04 F9 53 7E E5 13 D9 36 AC 7E A7 1B 0E E4
 26 9E 91 B7 F3 6D CA F0 EF 85 93 19 85 A2 8A 32
 23 1F CD 39 87 BD F0 B2 9C 84 AF 0C C3 50 F2 EC
 FD 83 3D 61 62 29 AE 56 8F 2D CE 34 B9 D7 A4 58
 5B 23 16 1E 30 1A 98 06 7E D1 27 7A 48 BB 41 D3
 71 E5 A2 FB 6E 45 0C 2E 2D D5 94 5F B4 65 7B C5
 94 EC 24 60 DF 61 9C 55 72 84 70 37 20 83 2A 5F
 5F 01 06 70 FB 69 9E B9 BF 41 92 25 7B 4C 4A 3D
 57 F6 CB 87 2D 59 1A 85 B2 29 65 E2 BE 87 FC 42
 7B 68 4E AA 6A 49 C8 7A F8 09 A6 7E 17 72 C3 99
 0B 36 D2 3B 94 30 E7 61 47 AA ED BA BD 9F 2C 31
 B6 69 DB D4 CB 6E 4A 33 C2 4D 64 0E 3E DB BA C8
 B8 3B 15 45 ED 2B 48 2F 49 2E 6A 75 17 5D C5 20
 26 31 68 E1 92 96 9B 97 E5 DD 47 55 33 17 92 F9
 D4 57 18 99 4D 68 F3 54 9B 21 B3 73 C3 81 B0 BE
 42 8D F6 E2 F9 0C 59 1B B4 87 D1 5A 3D 3E 4D FB
 8C 05 1B 97 BD A4 70 68 9B 51 1B F1 92 93 AD 3E
 7F 5E A3 DE 85 9C 35 05 A2 71 54 88 92 41 66 9F
 41 B6 4E A4 54 72 92 07 51 1B 50 F5 65 EE 3A 10
 C4 F2 0E 1D 07 04 77 40 2C F4 D7 CB EF FC FD 28
 2B F6 4D 93 17 0E 64 35 F2 F0 D5 C0 43 E2 14 AF
 A8 4D D1 C5 99 C2 DF CC C3 3C A2 97 04 62 75 1F
 E8 8E AE 3F CA C0 19 48 85 F3 F1 61 D8 8C 16 41
 6E DA 33 64 AD E0 3C BB 22 A2 7A D3 10 AB 14 E9
 8C B9 50 A4 E4 CC 08 56 5F 44 FC FE 45 63 5D 26
 71 89 FA 4D 69 50 35 D8 15 DD 9A E1 B2 78 B2 66
 59 CC 96 60 AC 52 2A 3D 31 A8 93 2B D2 34 19 83
 7D 39 63 55 36 88 C4 A9 26 57 6E 2F B8 9B E3 C6
 70 BE 6B 53 58 1E 41 60 24 32 2D BA DF 85 89 F4
 92 9F 7F A5 89 47 7D 0D 1D 2D 4D 63 CF F2 9E B3
 71 9F 44 CA 42 1E AE 9C 5B 44 BC 1E 9B 76 55 46
 43 42 45 27 59 6A FD 73 ED 00 F8 8C DB 35 76 A8
 5F 98 E4 2B DB DE 67 40 5C 99 EC 1E 58 27 57 FC
 D4 DE BD 44 26 4D F1 A0 E7 8F 6F 65 82 60 FA 79
 7A C0 8D DC 37 44 06 D2 A4 C4 BE EA 5E AD AA FD
 92 24 D1 2F 44 F4 B3 52 F7 C8 E5 A6 79 7F 0C 20
 7A 71 70 5E E5 58 D8 41 1B 3D 7C 4E D9 31 83 A0
 4E 4F 7F B9 BD 34 41 4D C8 B6 E9 C1 56 CC A4 23
 E4 1A 5F A4 B9 DA 66 56 43 DB 21 BD 1F 3C C9 12
 6A A1 E8 8A 4F CA 2B EC 46 28 EB 62 5C 3A F6 2C
 10 A7 F3 B8 28 2D 62 34 CF 60 7F D5 2D 51 40 F0
 8D 2C 6E 48 D9 F6 2B 85 10 5C F4 4D BD BE 7E BF
 DE 5D C8 0D 41 93 E2 54 26 EF 91 6B 28 B5 DA 35
 68 63 D1 37 27 1B 57 8B 4F 44 05 0A 5C 12 63 6B
 38 DF 67 7B 7D 37 FA DA DC FA C5 ED D7 68 0E 41
 F0 EF B1 6E E7 E6 4A 44 09 7B A2 35 E2 CB 09 B3
 A3 3A 33 ED 3E 82 08 C9 CB EB 09 45 B7 85 7F 4B
 67 1E 03 FC BD 23 C6 3E 40 86 60 85 23 DF F2 7A
 82 A9 1A F0 EC 78 6C CC 66 4E 90 92 AD DD E7 AE
 A2 FD BF B2 7A 6D 20 2E B4 26 02 DF 47 AA 4F 05
 2F 34 79 1D 47 A3 75 35 23 85 2E B3 C8 5C 8D DD
 9F A4 C6 0A D0 79 A3 E1 F3 A0 34 39 41 B0 1E EC
 E3 95 B8 39 A6 E4 39 B9 40 EB BA 10 3E 96 06 93
 05 34 33 36 87 BC 79 0A E4 49 5F C8 4A 14 19 66
 46 EB D6 57 67 B6 40 8B 71 E4 24 4C A8 22 E1 A0
 9D F7 8B BA 48 5E 37 74 42 87 31 AE A9 4B AC 4B
 5B 4F 9F 44 02 5A C3 BE EA 3D FB F8 48 5A 67 74
 E5 FD 50 FF 17 3C 2B A4 FC C7 F0 BF 89 B5 78 F3
 3D 50 E4 E6 BE 6D A2 36 CC C3 DE 5F 7C 90 81 F4
 C0 7D 0F A2 AC 29 7C 85 8C 21 6C 82 5A 54 88 49
 4D A8 84 4E 83 A8 99 3F 0B D3 B6 89 4F B4 00 C9
 44 9E D4 A0 B4 71 EE 62 43 02 93 34 A6 C2 76 4B
 79 F4 40 E0 EA 1C E3 E1 0C F4 62 26 E9 9E 9F BB
 B1 17 02 FA 74 CD FB C7 9E 41 42 06 DD B1 87 74
 67 04 0E CD DE 26 05 50 B4 3F B6 1C 4C 94 1A C4
 01 99 FD ED 46 8D C5 F1 93 70 3C 56 D1 26 70 5A
 DF F1 C7 EE 46 F4 A2 E1 AB 52 40 61 09 84 5A E7
 DE B9 98 BC 11 C3 0D 06 E3 CD 27 C7 70 78 89 F1
 9A BC AA 06 79 6F F6 7E 18 58 09 D6 A8 2C A2 B8
 CB F9 8E D8 D5 AC 3B CB F7 B1 12 F5 47 48 82 E1
 D9 44 76 04 31 81 FE 57 42 BD 81 4B 85 7D FD 36
 6B 07 ED FE F0 43 57 45 5B E5 DD 50 DF B8 8B 54
 8B 35 4F CA F3 CB 32 4B 13 FA 87 24 13 B2 06 92
 12 87 04 2B 49 3A DF 8B BB 52 37 42 DF 89 83 8D
 56 C2 C7 9B EC D8 7A 20 8B F8 A7 50 E9 98 EA 67
 71 C5 6C BD B0 7B 55 A7 1B 14 AC 73 05 9C DA 5A
 F5 4E 29 EB 66 18 93 23 CF C6 C0 34 09 91 C7 2D
 35 FC C5 3C 76 8F 71 CD 9C 4C D7 20 2A EE F4 42
 65 82 FF 73 7A 24 92 55 AB E2 5B C3 37 2D 24 27
 26 FF 1E ED 9C 28 78 E9 3F A4 CB 65 44 A5 B2 6D
 92 D3 F8 AE A4 1A C2 63 39 7E AB 95 72 0D 54 A4
 86 FB 40 68 54 B8 A5 C2 3E B5 68 D1 07 26 43 87
 79 B2 53 5B 79 AC 5E 8B 37 07 D7 17 6F 58 AC 99
 BB C9 B1 68 F4 F6 57 31 90 DE 34 CB CD 9A FE 30
 20 46 F3 24 60 4F 87 5A 54 61 92 D1 3B 54 41 62
 41 38 25 CF 5B D4 64 8F 83 29 D0 74 DE A2 26 57
 0D AA 29 4C 14 87 19 A5 1B A6 3B F4 5B 07 F6 7E
 84 72 BF 9D DD AC 37 3A 20 4B D2 FB 52 DF DA 01
 BC 7B 4F 27 8D CC 24 51 3A E0 05 04 DA BF 9C 0A
 6A 24 90 A5 8D 28 16 F1 78 77 FB B3 95 5D 51 43
 1B AC B1 F0 45 28 37 07 5E D4 9D 7C C1 B1 3D C0
 BA 73 2E CF E8 D3 E6 D0 9D 45 6E 51 B8 C1 5E A7
 D5 E1 E2 95 B2 CE 79 9C 00 17 2B 5D 07 B7 A5 22
 5A 78 8D 39 14 3C 94 02 35 7E A9 55 F8 BF 6F C4
 3B B7 23 08 B1 9E C3 CA 5D 15 91 A9 C9 A1 45 20
 55 49 12 01 62 0E D2 85 02 20 78 54 6C 21 AF 5D
 FF 04 61 4D 54 E7 27 90 1E 79 04 20 A6 1F 37 5A
 AA 42 93 D9 DB A8 01 C3 28 6D 30 31 E6 24 D8 7D
 88 C4 3A EF D4 54 02 65 06 1B 40 02 41 48 FA 71
 8B BF 00 94 A5 F9 EB 17 99 CA 46 00 3C 53 F4 0E
 42 AA F3 E1 2C C4 49 7A C1 54 7E 8D 42 E4 81 02
 A0 8D BD F7 C1 A1 B0 19 3A 3A 7D DE FB 2E 11 61
 18 D9 F6 C7 6E 9B 7D 21 AC B9 09 01 EB 6F DA E4
 A6 C0 B3 C7 C0 08 A1 4E 6B B3 D6 9B AB A2 65 86
 19 3B E3 8E 56 8C 2D 51 FC 08 80 90 91 54 56 73
 E6 3A DB CB 55 13 F3 79 A1 5B 4D 1C B0 09 66 94
 6C 60 B6 F8 9F C6 46 48 E1 AA 8B B4 2D F3 22 75
 CC 79 3C FC 7E 12 E5 10 9B 23 D7 B8 8D 34 85 07
 CF AC 77 CF 02 B3 2E E1 A3 46 E0 34 33 55 B8 07
 4D 61 17 70 DF 54 09 B5 99 10 59 31 9B 3A 88 81
 B7 21 4D CA 8F 87 48 94 E0 EA C7 64 31 3D 92 92
 2A AB F0 CD 0F 8F 73 98 CD 05 8D A3 47 E4 9F 20
 F6 7C E3 B3 65 28 A0 2B 42 BC 01 8D 0F 8C F6 0E
 AD 4F 66 E0 B3 19 4A FE B8 30 F8 24 08 5D CC EB
 47 7C 80 DF FB D8 97 B9 63 6B 35 DA C3 F6 64 C8
 7D D4 97 36 10 33 2C 47 D3 FF 56 7B 9D A3 D3 4F
 14 03 EC 2E CE 44 80 3F 3F 66 DB FB 50 4F FF F7
 E5 8B 16 C4 1B 1B 93 87 D2 2D C1 28 62 3A E6 9B
 60 34 B9 0C 46 A9 92 CB BC 9A BD 22 14 DC 1B 8E
 51 FB 3D EE D4 1B C5 72 54 5D C3 F1 0E 6A 18 38
 AF 6D BC C5 F2 9A DC 8F D5 03 A2 4C 35 B1 6C 58
 A7 BB 20 5C 11 12 A0 D5 EE 4A 7D 98 58 B1 3A 17
 15 FD 94 06 45 D9 52 6E 06 53 8E 43 26 8A 44 30
 E2 80 D7 96 C0 62 BE B5 3F 8C 19 8F EA B8 C6 A2
 45 67 70 8A 68 10 4A 58 0E ED B9 5F 72 2B 6A 48
 C6 6F 45 E0 48 2D 40 FA 9A 6C 95 AA 14 70 C5 E2
 B5 D8 EF 83 99 AD B5 D5 D5 73 60 6F 46 3B 70 0E
 B5 C3 70 6B A8 37 26 18 E5 90 52 1D D7 7F F2 C3
 16 87 92 EE AE 0C 4A 88 F2 3A DA 38 90 5A 46 E1
 D6 2F 77 7A 44 4E CE EC 84 73 35 BB 79 34 3E 3F
 98 23 86 29 A6 57 21 4B 10 66 B0 59 D6 F3 7F 79
 6B 1B FD 72 A3 56 99 7D EB 36 19 5E 2A C9 DD FB
 A6 07 2D 79 C8 CE 2A D8 2B A0 C8 C9 3E B6 8E 8B
 8A 41 20 0E 37 0C A2 57 CB D1 90 36 A3 9F 9C A5
 BD FB B0 AB 78 F9 E1 69 8C E3 1A 36 DB 1B 44 05
 BD 3A 29 95 E5 D6 EE 72 5A 9E EA 9B C7 D3 D9 81
 6E 90 EF 2C 4C 01 33 34 15 BC 6C D2 13 7E 4E D3
 F9 F4 F3 A1 E7 C8 30 3C 63 1F 34 C8 F3 ED 51 64
 1B EE B1 F1 0A 99 5F 66 6A 80 06 FF 51 91 70 38
 35 39 6D EB 35 89 3E AB B8 A2 CE 79 78 C0 C0 17
 F7 88 5D DF EB 50 3E D1 35 FA 63 22 2F FB 1A 42
 2D 68 E5 A0 D8 74 81 87 06 03 E6 E1 4C 7F AA 32
 AD B9 A6 AA BA 4F 32 95 70 8A 0F 1D 62 90 FC 8F
 09 66 BB 85 BC EF 34 11 F3 72 27 AB 65 7F 09 A1
 0D 5A 92 FC F0 1F 0C E8 AB 87 BB B6 68 5D 18 FF
 57 48 86 7B AC 89 D4 1A 7C 9D AC A2 B3 7C 7D 54
 8A AF 7D 34 BB EB A6 60 DF AC 8A 38 B5 76 90 BB
 7B 6B F2 F1 7C 50 76 30 C2 F4 2A B8 9D FB D6 3A
 DF 1C 00 A6 DB 57 C2 9B 81 7D 66 D7 9D 22 C2 34
 98 71 F2 FB D8 A2 27 3A 1A 94 4B 38 CD 47 E1 CB
 C8 8E DA AC E9 59 F8 0D D0 69 DC DC 57 F7 1E DD
 20 20 E8 80 45 B6 AE A7 56 7A 50 DC BB 0A B6 11
 34 74 34 61 02 22 90 76 EF 14 07 9B 3B CD 08 D0
 BB E7 23 44 88 36 AD 12 70 E7 18 98 0B F7 9C F6
 15 93 57 BF A1 F9 EE 80 B7 7C 0D C2 88 0B 7D 81
 43 EC 39 5D 9A 78 B1 FF 8E E9 95 D3 99 2C 40 2E
 73 F4 70 DB 2B D9 67 E0 C1 AC 27 F3 13 3A F0 BA
 B5 F0 BD 0C DC B4 43 09 61 E9 2F 55 DD B7 E6 67
 C2 60 B0 36 75 A5 57 88 BC 2F 43 84 4D A1 AB D6
 80 77 19 23 56 13 57 C6 7A 0D 51 5D 54 33 96 70
 D6 50 BA 0A BA 62 20 18 46 59 71 F9 67 9C D0 00
 25 23 CF D2 D3 71 65 47 F4 FB FB 5A A9 DD EB 1C
 81 74 2F 93 0F 5E 9A 65 CF EB 79 46 42 75 28 08
 44 BD FD 80 49 FA 1B 41 77 39 AA 0B 7D 5D 8E AD
 01 AE 42 FE 1B E4 F7 61 99 BE 79 EB 72 B3 EF A5
 84 B3 A8 FE D7 3C 5A 13 ED 58 78 AB 39 5E 23 53
 DC D4 EA 73 06 A8 87 36 03 EC 96 69 7E E0 38 16
 0D EA 12 64 BB 0E 9F C7 9E 2D E9 57 C0 FF 33 3E
 E0 CC 3B 58 5A 33 9F 8B 85 D7 C2 82 84 09 2B 7B
 FE 8C 22 69 49 22 E6 8A 56 83 43 07 9D 5C 5F AA
 CA 26 B6 E9 E4 FA 50 96 2D 0C 82 4D 03 AC F2 90
 82 BE 20 8A 8B 29 C2 22 1D 06 09 52 2C CC C6 E2
 F0 26 E8 5E 83 A3 BB 75 A3 28 39 97 C7 89 71 39
 0A F4 44 5C 28 CF 3B 53 42 7B 2F 6A 24 A4 76 8F
 F3 90 0C 1F B2 F0 B8 6E F0 B8 AC B1 B0 E3 85 FB
 2A F3 B3 55 E5 2C D7 2C 17 3D 2A 83 27 3A 96 0B
 9A 67 58 FB FC E8 68 65 D2 A2 B7 44 A6 03 BA 8B
 44 58 9C 94 58 79 17 B7 91 05 C8 6C A8 34 6A 2D
 2A C5 DD CC C4 85 A6 37 76 2B E9 4E 66 4B 19 72
 80 AD FE C3 80 70 5F D6 E6 C4 91 C9 5C AA 29 97
 ED CE 3D 57 26 76 12 BE EF 4D 71 52 59 1F 5B A1
 41 70 A0 4B CD A6 66 73 F5 30 48 09 5D F4 3F 96
 53 E9 08 D9 6B FC 57 48 C8 DB BE 34 9F 01 B8 23
 26 6A F0 20 6E 63 52 56 EB 64 44 F5 FA 91 4E 75
 35 56 B4 A9 82 44 C4 B4 FA 9A 22 BD B9 95 AD 96
 E2 C3 52 B7 79 3E 86 09 09 C9 BB A9 4E 53 55 CB
 C3 5B 3B EA 4F B8 50 6D D4 B5 94 1E 3B 58 13 C8
 02 C9 A1 A6 1E D3 E8 FD 29 6C 40 5C 10 49 46 E1
 A9 20 CC 9B BD 15 6A C2 2A 97 FE 67 55 31 B4 6C
 4C DC 92 16 C2 79 74 43 4E 46 A0 C8 90 AD 3C BB
 A2 0C B7 A6 E9 67 52 BD 2E 43 EB 34 B8 7E D7 8A
 75 D5 BE 64 80 07 97 6F 8F 1E 52 C8 81 D2 86 E4
 75 97 D8 3D 75 B0 CB 3A 57 29 AF 45 6C 08 3D BE
 88 8B 7C 1B A6 AC 48 6E 00 18 85 0B 53 16 9C ED
 FE 9F 22 73 3E 8B D8 AB 53 4A 17 72 C2 C5 2E 7B
 3F F1 33 C2 BB 2F CC 8C 89 91 42 D1 9D 83 AF F5
 ED FC C9 E2 2C BD 2A 49 E8 A6 64 60 5B 1E C3 93
 92 7B 91 B6 EA 5C EA FB 43 E8 B7 D7 CA 2E C8 1B
 AC 36 96 1B C4 A4 9A 15 F2 4C 47 B7 D7 BE AD FA
 E8 19 38 62 1A F3 48 B2 72 23 2B DC 97 4C 1A 1B
 00 74 9E 12 5D 89 CD 5C 0F 1C 9D 94 F2 D1 FD 55
 FF 0D 7D 3D AD E0 AE 87 EF 7C 95 BC A2 0D A2 42
 63 00 71 5F F2 56 83 6C 10 C4 A2 60 0C 27 00 61
 DB A8 5D 7E 9A B0 6D A2 DD 96 EE C7 07 C7 67 DE
 19 C6 21 CC 3A F2 57 1E 91 1F 68 62 E2 09 32 2D
 70 F1 FB 3C CB 77 17 CF E4 16 D3 D6 5B B0 19 2B
 E3 68 80 22 A1 54 81 EC F9 C0 27 BD 95 A9 BE A9
 96 C7 60 27 DC E3 43 1C 92 51 55 47 1B 7B 92 F9
 1F 41 D4 C4 43 D1 BC 1A 04 91 22 0E D6 FD 76 39
 EA 66 FE CC 7E 2A 1C 01 67 B8 6B C6 5A 95 E0 CD
 29 75 CF B9 CE 68 F0 C0 34 56 56 B8 19 3C 27 08
 C4 A8 62 04 22 14 F9 75 2A 6D 08 A6 5D C3 EC 1E
 83 F7 50 50 05 41 8A 2E 68 64 5D 0C DC CC 03 BE
 E7 80 C2 58 0F 3E 82 D0 7F D5 DD AF 0A 6D 0B FB
 C0 55 70 A1 84 16 D1 C3 08 FC 1B 58 9B 1B 51 85
 EF E2 1A 16 B8 5F FE 12 CB 26 6B 4B 18 B3 6D E9
 55 A9 82 FB 87 FA C2 9B 2D 7A 22 73 4C 1F D7 50
 49 7B FC C9 F5 46 7C 7B 1F 96 E1 49 04 26 5F 71
 8D EB CC A7 56 1D EA AF 85 7F E3 41 D4 2A 98 BB
 7B A9 A2 82 E2 9D CD AA 30 D9 60 6A E7 0A EB C2
 27 4C 17 DA BB 9D 7C 73 B9 54 19 35 38 C2 6E 20
 19 68 24 C6 59 7E FC 8E 0C BB 6E 6F 59 3F 36 7F
 3D 49 67 6A 55 22 77 7E C5 87 74 71 17 1B 3C 28
 69 12 D3 EB B2 DA 76 2D E3 43 FA FD D1 72 B2 42
 E7 6E 0E 1B F3 3D 25 5E 5B A8 76 A4 B1 A2 4D 9A
 BD EE 7E AE F6 CA 44 89 DD 14 EA DB 72 39 89 A7
 98 B1 62 FB 9E E3 D2 27 23 DC AE 47 D5 B8 B3 21
 00 91 27 A2 55 26 A1 89 CB C5 FD 52 60 DD 6D 83
 A1 BF 80 99 5F E6 ED 09 78 8C 2A 2B B4 AC 2B 83
 CE 17 C4 AE 71 D5 79 04 E1 7A 28 A5 3F 43 38 A5
 08 80 06 D1 51 A1 05 11 6B 42 F5 00 13 A6 B1 CB
 50 8C 8A 2C 92 01 7D C7 6C 78 70 E5 44 9E 91 6E
 58 FE 9F E1 FD 5C 9C 83 0D 82 B7 DB 9B 21 CB A6
 BE 61 E9 3A 3C A9 62 28 CB 39 DC D3 9B 7E 62 C8
 AB BC 83 25 15 C5 EE 81 ED E2 0F 27 4E 16 82 22
 F0 1F FA 7A EC 26 6B 1C B5 94 00 A7 20 83 69 67
 28 43 DA 21 68 40 FB EA C1 EA 83 A2 AF EE 32 36
 79 91 FB 20 B4 09 06 AE 02 43 86 C7 BB 2A 1D 27
 A9 F8 6D 95 BB B1 35 E0 FA 8E AE 8E CC 4E E2 23
 25 B0 83 B3 C0 17 17 C1 C5 3F 9B FB 61 A5 37 E9
 E0 EC BC 75 2A 9B 2B E8 AD DD 4D 13 F7 4A 28 F4
 84 50 27 2F 60 FE 60 BC 82 3F C2 4E 45 87 B8 B1
 65 93 65 D8 0F 8B 24 1C 18 DB 84 37 2E 03 1A 8C
 F6 15 14 2E E5 F9 96 48 F6 69 E4 DC F2 1E 63 4F
 A9 55 1A 99 A7 03 C4 F6 5E D9 A0 66 CE 66 B8 93
 86 C2 CD 8B 80 E1 31 A5 8F 41 38 83 34 E9 2B 97
 BF 07 0A 5B 27 A9 13 06 2F 01 EB AF AD E7 4F 39
 C5 3E 65 30 C5 DC EC D1 78 97 FB 41 B0 F6 B3 9A
 54 5B A1 41 8A 2F F8 0B 2D FF C2 45 4E 42 CC 61
 57 95 1A 8F E7 EE 58 23 BE 5F B1 2E FC 4F 3F AA
 46 B7 7B 16 01 68 BC 7F 40 AD 70 85 ED 8A D4 4C
 69 E7 85 AD 87 1C BF 8E B2 5A F4 43 64 B7 50 8C
 B6 59 CC F1 40 96 F9 55 59 92 07 49 5D 40 B6 42
 82 2E AC 3A 1B 7F 0B B7 48 4E F5 9D 8D 34 FB 7C
 48 A4 3D 03 DD 2A 15 2B DF 01 EE C7 AE 86 90 99
 67 03 AE 95 5D 92 05 5B 76 C3 67 C1 90 3A 4B 19
 F4 AD 51 5D 35 DB 88 B2 2D 45 CE 03 A3 07 4B DD
 F5 CA B4 EB D4 DB 22 CA D2 45 FD 59 DB 31 7B BE
 A5 8F 9D F2 5D FE 24 97 D1 83 14 5F 29 78 70 ED
 9A E9 DC 64 0C 16 5D BE C9 13 1E D3 EB 21 3B 38
 A8 72 EB 9F EE 5C 4B E8 32 3D 5D 65 B2 58 10 C0
 81 3A 5B A1 2C BD 1D 86 A2 A4 3F C2 44 D0 BC E8
 E9 BD 57 DF 84 FF 8C 57 5D B0 C5 7B 41 C8 E0 A9
 F7 4C 3E E2 44 24 F4 A2 76 0A EA D2 F4 E9 E5 30
 F6 CF B0 93 BE 1D 77 71 7D 42 24 2E F3 6D 7F F0
 46 E4 08 73 DD 00 40 87 7C 8B A6 C4 B5 9A 40 5B
 1A E6 64 5C B8 D3 87 F2 5D 30 E6 6D AB 56 9B AC
 96 3E 78 2F B0 4D D8 7B 94 7A F4 24 E7 75 C9 7E
 47 6C 0A 72 F5 E9 B7 50 84 4F 69 48 71 C4 23 DE
 77 1D 45 D5 2D B0 1E 93 DB A4 10 EE F3 92 58 3B
 07 3A 49 06 62 78 F0 7E A8 D6 12 C9 9F 13 E5 70
 FD EA 12 A1 D4 29 80 B6 EA 2F E1 C2 BF CF 09 92
 4B 2E D6 21 75 18 32 B4 79 BC D5 C6 CF 12 7C 5C
 A6 37 DF 1E 4C A4 55 B7 D3 34 CD 00 1F BE 45 DC
 1F B8 B8 F1 C5 76 05 18 83 FA D3 0F 4B 89 B1 2E
 B5 ED 61 26 7B 8F 97 EE 1C A5 6D C7 19 91 5D 94
 CE 18 D6 A4 70 66 45 8C B5 49 86 4B BB 66 AA FF
 D2 DD 8B 43 DD 1F CB F6 BC B3 DC 7A 2B 3B E9 1B
 A4 DE 5D B1 58 7D 33 5D DD 28 D3 EA C7 BA 45 E9
 1B EA 4F FC A2 DD D3 0D DB C6 97 39 40 00 6F 2B
 B0 A9 29 5F 1E 1D 16 6C F4 64 A2 67 EF B3 6A 49
 CF AD 79 22 65 80 48 27 CF F7 F1 95 50 53 84 FA
 C1 89 8E FB 0E C9 80 71 A0 95 56 37 6A 6E 60 59
 17 A4 18 9D 6D D9 B0 20 8E 9E B5 70 87 62 1C B2
 31 4D 76 8D 08 F8 74 6A 2E D0 B3 CB 86 35 F9 67
 B9 11 DA 58 59 DB 65 CC BA E3 A3 4F 26 0A 9F 8A
 12 03 F4 84 7E 9F 90 1E 57 F1 DF F1 5D 33 EE 48
 E0 83 91 A2 52 F7 55 9A 58 71 53 95 DD BE 13 6A
 35 86 79 06 72 F8 31 70 12 55 41 BC 9E 36 D9 5A
 A5 80 53 45 B0 D1 B2 21 E0 B7 C3 A1 28 1A FA 34
 B0 E9 FC 89 C6 DF BB 89 C8 24 A3 91 BC 99 5E 73
 7E 49 88 A5 C5 CD 68 7A 44 EC 2D 34 88 0E 34 B6
 EF CE BF BB 52 1E 0A E5 3C 77 5F 62 38 04 49 37
 58 7F A9 7C 3C 62 5C 9A D5 36 CA 0B 54 1A CE C1
 EB 52 5F 0F 4A 50 75 BC F5 22 52 0E AE F5 81 A2
 52 31 31 20 51 3A 42 14 C4 B4 AF 00 74 8F 8E E3
 F6 71 22 EB FD D1 DD AD F2 71 34 B4 08 12 66 0C
 DA B3 9D 06 85 13 5C 3A AB EF 74 B7 38 10 A3 6B
 BE AA 4C 7F 30 EC 48 59 68 1C AB DC 3B 92 74 9E
 07 D9 5F 4E B8 FD 75 66 DC 22 1A A9 30 D9 97 CD
 E4 5C D5 4F 64 3F C4 85 21 A4 03 38 01 67 B4 86
 F0 9D 41 5B 78 EB 1B 60 11 26 20 70 16 B9 9B FA
 70 FE 91 10 0B 20 4F 1D 72 4A 1D 3E 0D 48 4C A8
 49 D8 05 A6 57 2C 40 DD B6 0C 60 AD 42 A7 A3 19
 65 56 CF 46 07 22 95 04 4D 18 19 12 73 0D 71 16
 0C 0F 67 63 35 3E C2 A5 83 C1 C5 00 04 F3 7A DB
 E0 2B 8D 51 A0 CE 01 14 68 37 6A 49 8A 2E 54 00
 4C 5F F9 CA DD 45 49 1F 65 B1 E1 CC F9 00 BB EB
 25 BD D1 C1 1F 62 2C C5 11 28 41 DB F3 83 01 02
 C8 89 0F F5 83 E8 84 BA 9F AF 3D 31 B3 01 32 94
 77 89 35 B8 C9 9B 1C 4D 0D 8C 50 1A 2F 02 BA F4
 E1 88 87 FB 3D 29 B6 10 4A 8F 20 24 A3 FC A0 42
 63 10 50 27 ED 26 44 A6 3E FD E4 FA E7 F7 D6 C3
 D1 A4 CD C5 EF 01 B0 FD F5 73 13 E7 75 16 C5 63
 AD 29 89 F7 50 B5 5D 49 9D 32 A2 63 2A 28 85 0B
 1E 47 28 1F 3B 40 3E 8D F7 1E 06 37 04 C4 D0 89
 8A 3A FF 36 5E 85 B9 0C 91 E8 79 55 50 C7 ED 6E
 3B D3 3F E7 4E 5A D9 D4 4A B0 7A 72 AE 38 FB 2C
 B5 AF 41 02 69 A2 61 A2 72 F4 06 2E B6 78 31 A8
 99 D7 9B 1B 12 FE 49 05 8D AE 00 B8 32 37 71 5B
 66 AA CC 22 3E FA AD C9 31 1B 8D EB 55 B5 FF AC
 6E 20 4F 85 6F F6 9E 63 18 BA 15 48 4B 36 54 1E
 9E EA 88 A1 99 78 A1 41 8C C2 85 A9 30 3B 49 C0
 07 F1 97 7A 90 2B 2F 38 8D 30 74 3E 7F 73 7C 17
 5C 1B 97 A8 5B 3F F6 90 4D 3B DF C0 31 68 E1 ED
 F5 F8 D3 C4 54 00 67 81 88 10 F7 E3 17 83 75 5F
 83 CE 30 B3 5A 7B 57 A5 DF 57 2F 42 55 65 95 2C
 C3 08 B2 D0 D8 84 A8 2C 74 C4 4B E8 35 CF 33 EF
 FF 4D FD 2B BC 04 6F 7A F0 E6 A8 EC 49 4F 85 62
 61 5D B3 C6 B1 E4 42 6C 05 96 2D D2 CE 31 78 8D
 87 30 41 AA 2F BC DF 4F AA 57 BB 7E 52 EB 30 FE
 B7 74 D5 6F 5C C6 5A 29 3C 3C 6C 01 18 97 F1 EB
 8C 17 70 4C 14 DF 7B 5A 32 67 70 42 D2 2B 2E EA
 06 66 A0 2E 80 99 58 98 E2 A8 91 C7 F9 BB 58 16
 00 1D 92 3C 6B AA DB F6 14 F2 C0 84 B0 BE 01 93
 60 25 1E 6A 52 FF BE 14 4D 95 77 09 01 B0 8F 44
 43 3D 29 D2 41 59 45 73 4A 34 1B 4F 6C B6 45 38
 70 26 34 BE 2F B2 63 F8 81 3F 66 A9 5B 1F 09 31
 B7 23 F2 3A 98 C1 8D 84 D1 BC F0 3D 22 39 9F 34
 83 94 53 47 AE 64 BF 0A 4A 22 32 F0 E4 42 F6 9F
 AB 45 FD C1 D6 25 70 65 F0 74 8E F0 58 E3 38 74
 B3 4B E0 10 D9 8E DA CA 1D 8C 59 16 ED 1C BF 91
 04 EE 59 1F 23 73 2E D9 DB 74 24 B2 5B 24 1B B7
 2B FA 0B 22 8D 3B F6 85 22 CC D9 C6 77 8D D7 5C
 D8 D3 A8 FF 7C 6C 76 AB 7B 88 4C FF B5 6F 01 FD
 2A CE 2F 5E 2C 32 14 62 AB 0C 1C 41 4A 91 8E 89
 7C A6 4B 6A 8D 66 4E E4 BC 14 8E F9 6A 19 27 BD
 6A 31 FF 43 8B 72 C3 98 0E BD AD EE 86 66 39 73
 76 F7 5D 12 79 C0 E5 F4 5F CD 8D ED 61 71 CF 1E
 5C 36 86 ED 0D 9D E1 67 DC 47 21 74 22 B9 E9 B9
 44 5D 44 6A C9 BD E1 83 FD DF 03 82 B0 8B E8 F5
 10 C8 EF 63 A9 68 40 48 DC D1 EC 79 77 B6 A6 09
 C0 48 42 DE EC 42 E4 11 A1 32 4C 64 89 15 AD 29
 EE 93 8C 07 4C 0D 96 52 4A 5A A0 8F BE FF 8A 4A
 82 22 35 07 0A 41 31 78 8B FC AE 98 F5 BB FF 65
 E4 3A 2E 7E D6 9A F4 0A 5A 8E DE 93 3B 79 8F 32
 17 9A 73 B3 40 D4 83 30 8A C0 94 5C F5 8A C1 2F
 22 1A CD C0 2C FD 4F C5 FD 97 17 2A 2F 2F 4F C6
 0C E0 FB 88 96 E5 4B DE 5B E9 9E 8B 83 8C BE 81
 73 68 9B 72 F5 0D B6 79 D6 F8 7C C8 7F 4C E3 08
 25 4D 9D D6 44 80 7C B0 92 E3 01 C5 B4 D4 32 EE
 D7 0A 32 13 C4 0C FA C6 A5 46 3F 5D D3 BD FA 11
 79 11 57 19 3C 46 10 34 F8 78 44 D5 D9 5F A7 CA
 C7 16 8B F2 6B 50 98 4B 4E 3F B7 53 AB 7A FD 3D
 6B 67 D1 AC DB AF 67 0F 51 5E F5 8C CA D8 92 4C
 10 89 4F 74 C4 5E A9 19 A4 9E ED 2A 87 5A CC 48
 5D 6B AB 40 15 14 9B F9 69 72 CB 44 CB 1C DD EF
 E4 51 E8 EE 22 4E 29 18 FC 05 D5 99 40 2D 67 73
 F5 12 75 40 5F D4 C9 4A 0F 7D 1F AF EB 48 35 E3
 2E 53 DF E3 44 FB D0 4B 0E 80 74 74 94 CC 38 7F
 54 50 72 AE F2 C6 D3 F6 CA DB 98 28 26 A6 34 5C
 0B A7 BC 80 43 E1 8E AE E2 11 53 91 DD B1 39 2A
 B6 1C 99 BD 41 67 80 8E 7E ED F3 39 2F 11 FF 5D
 6C DE C3 19 2B 5A 27 1D C1 7D FF CD 69 50 6C 2E
 B6 A3 CF F3 6B C2 E6 AD 59 23 97 B8 CC 16 63 17
 FC B1 FB BD 39 59 55 54 C2 6C 91 47 18 4D 04 DA
 A7 76 A6 E7 1D 29 46 70 3F 3F 65 61 0F 3F CE 2F
 AE 91 0A 6E 05 33 B8 68 FF 02 41 CD 23 DC 15 E5
 A9 AF 98 3E 54 8E FB C2 96 E9 58 DE C0 08 EF ED
 7F CB 06 A5 E7 F9 17 6E 2A E1 EA 7F 99 CB E2 18
 B1 F4 A2 76 9B 9C 7F 0C 1A 00 78 81 23 81 24 76
 55 A1 91 55 DA 45 7E 79 62 9B 24 74 5F 72 09 E5
 9E 14 22 38 5E B5 D9 45 6E F3 B0 12 1E 11 CF 1B
 CC A0 B3 1E 63 78 9D 4B D5 74 EA B5 2D 71 B1 DE
 AD C1 1B 86 68 D8 FF 22 A8 1D 0E 40 22 30 DC E4
 A0 5E 7A D8 FB BA 0D BF 6F 10 D5 D8 52 01 FE E6
 4C D7 D1 FF C3 40 DA BC AF F6 E6 B3 3E B9 78 6C
 33 BD D4 A2 9B 10 2D AE 28 58 87 0C 2A 22 93 DF
 FD 12 D8 83 E8 0F C7 F2 F0 27 A9 C4 9D 0C 5B 81
 DE 25 C1 B0 D9 5F 36 2B 7F 41 3D 35 EA 7B 3F F0
 16 25 05 C2 3B F8 89 E7 92 A2 FC F6 63 57 31 9E
 BC 1B 3B 00 6F 4F 99 FB D2 51 FE 7F DA DE 93 82
 94 75 BE BD 07 24 19 8C C5 1B 59 CC C6 94 53 74
 F4 EF 15 B5 8A FD 95 B6 6E 4A 3A 09 B3 A9 0E 14
 01 36 D1 5E A5 C8 4E E5 4C F5 6F 9F 27 CA 3B E5
 41 24 CA C8 AE C7 BD 35 28 3A 73 21 53 7F 2E FA
 88 21 C1 FE A5 81 95 1D F6 77 13 19 77 62 0F 56
 E4 A6 94 5E 04 BC 5D 13 86 3F F7 A4 9D AB 62 9F
 B3 D2 46 62 C9 75 5C 36 CD 30 47 44 67 40 32 01
 71 37 54 09 EA CE 13 CF DA C5 82 58 F3 86 2D B0
 4C CB B7 BB 0E 46 3B DC 7C 80 F6 CE F4 48 C1 41
 85 95 55 42 B2 BE EE 15 3C FB 4F 5D 58 76 C8 C3
 3D CA 27 83 C1 50 19 92 04 F5 62 68 ED 36 AF 9E
 B2 D6 44 49 DC F3 68 69 E3 B6 88 1D 8D 6A 0C 8F
 6A 33 20 FE 49 8B E1 B2 CF 06 23 39 EE 2F 04 46
 B9 DF B4 E3 11 D6 24 27 7A 40 FD 42 A1 AE 97 36
 0B 74 85 A0 C5 9B 97 6A E6 30 A0 C3 1F C2 6D 55
 3A 2A 66 3F 7B B9 CB 34 00 6B C2 3D 07 7D 8B F9
 1F 9E EF 01 93 D0 BB 66 8F FD 0F BC 73 A7 B4 84
 FD BE 1C A2 CF 14 A2 BD AA DF 6B FC 47 99 16 00
 65 02 B9 91 94 D0 9E 33 48 D1 DA 41 04 89 16 F5
 55 1D 51 3E 43 AC ED 0F C1 9C C8 48 58 DF BD 15
 F5 68 74 88 95 39 7C B1 94 00 E3 8D 14 90 A0 63
 FF 17 67 C5 EA 39 24 E1 B0 4D 05 8B 9F 5B 45 4C
 91 BE 56 10 AE B6 58 FF 99 D9 7A 3E 62 A4 A0 27
 07 E5 20 FC DD 8B D6 AD EB 15 B4 6E 8A 46 A9 3F
 C9 B0 09 B6 B0 2F 45 79 0E 07 30 AA 60 00 AE A3
 50 32 88 56 AB AF 06 95 0D D2 AB 1A 99 29 30 C0
 AA E2 68 FC 34 AA 02 D3 8F 63 A6 7C 93 93 0B F4
 48 05 C6 61 A0 CF 78 9D CE 21 99 D9 16 E8 DC 37
 94 CE 52 21 30 30 7A D9 D6 94 41 D8 B6 EE 3C 60
 63 AF 29 F9 88 1F 8B 93 6F 53 3E 4A A9 0F 30 4C
 95 E4 CE 4E FD 71 A4 80 1E AC EA BC 34 22 5C 55
 09 86 37 0B EF DE 6A AC 86 62 8C 01 7A A1 F5 F1
 59 7D D4 13 B2 B1 51 2D DC FA 4F 56 DE BF 59 3B
 48 39 34 82 AB 5B 32 46 19 33 9A 97 62 DC 43 F9
 93 8D 20 45 57 FB D4 1E 9A 5A A9 5A 45 60 C3 D6
 DC DD 8E 63 D4 92 F3 6E 9F F9 FB 6A 97 A1 52 2B
 64 65 A1 87 2A 27 59 A7 8C 36 57 32 CD 20 E2 15
 6D 14 EB D7 50 4D CA BC 35 9C AF 87 2F 4A 9B 49
 49 3D CF 01 17 6D 0B D1 74 A4 68 4A 88 24 2C D7
 11 12 24 84 1D 44 13 0D 7B CF 3D F0 3C 44 6F 89
 C2 BC 0E 4E 68 3C 6F AC 98 25 D8 A4 23 C7 53 89
 62 C3 20 4B 7D 4F 62 DD F0 EC 80 D6 C5 60 9A 70
 02 EF 1F C3 0A AA 76 A5 06 60 C9 7F AD F0 64 84
 F3 FD 88 68 D7 BC 84 1A DA 65 0F 6B B0 73 D4 CE
 B7 E7 AC 87 EB 7D 25 42 8A 41 A6 20 9A DA 8D 7B
 AE 7D C7 DA AA 30 04 11 88 39 F2 31 79 42 AD 6C
 4E 22 4B AA 25 DE 6A 9C 91 BE 21 4D E5 CD 93 71
 82 05 43 78 05 9E 4B 69 8B C3 A9 F1 F4 AD 55 AC
 92 DF 25 19 FB A3 34 D9 C5 39 03 33 AF 42 39 AF
 09 C0 A8 04 7C C3 57 EE EC 2F 4B B6 27 7E AA BE
 5B 07 86 78 CE 0D 42 8E FB BB 95 20 35 EF E9 4E
 06 1F 63 24 33 88 3F 9F 3F 39 DB 68 BD 42 3B 21
 49 99 E8 E3 DB CF BB 6D 42 70 9E FF 13 95 B2 08
 BE 15 6B 9F 6A F8 67 C9 4C 91 29 38 29 75 85 39
 DA C4 CE 42 41 40 5E 4C B4 41 8B 5C 56 3C 77 FB
 2F C1 75 B0 C4 B5 F4 FA 79 14 1B 55 BF 39 49 06
 61 AA E5 32 30 0E E4 A7 52 01 BD 8E C7 87 83 35
 5E E2 12 34 01 14 D3 D2 76 BD 14 B0 0B 1A 32 B2
 DF 3D 1F A8 10 DB 0C 95 EF A5 A4 32 99 B1 0A EA
 CA C8 F4 6F 06 48 39 BC D6 C0 B9 F2 3C 43 5C 8E
 87 97 B0 29 55 C0 08 A4 BA C2 79 B8 67 AA D0 2E
 9E 77 32 F6 A2 49 4B 6C 9D C0 18 06 C9 A1 4B 74
 4A F6 D5 6D 7A A3 E8 7F 13 FD 55 82 0D 27 2B 04
 13 D2 B5 0F BC 9D 3F E4 28 CF C3 5C B9 78 4A D0
 6C 4F 25 39 5B 57 16 DB 4D 46 23 39 E1 9D 72 EC
 22 F0 C8 63 B1 7C 63 BF 38 51 BF 1F 7C 78 E8 AB
 62 1C 76 7B 2D 46 9B D0 97 47 17 FD 14 64 85 AA
 DE C0 82 BC 11 E5 6C F1 FC F4 BF 3F 6D 54 BD B5
 48 22 B1 96 AA 34 78 07 B3 58 F2 99 0F 6C 81 76
 3F DC 3C E9 62 32 3F 21 E6 1D F4 B7 75 7D 7B 57
 5A E7 57 D3 42 12 B5 8C 27 FD 1B C0 1D 69 7D 57
 CF 51 EF 33 89 23 EF 0C 21 7F A2 90 B0 B1 7B 23
 A6 B9 03 97 41 A0 E5 13 25 0D 45 D9 95 1D 52 06
 BC A5 EA C6 D6 CA 67 66 90 77 6C E8 B4 13 27 50
 54 6B 29 7B 59 3E EE 38 7C BC 1F ED B8 06 1F 54
 3A 44 67 58 6E 73 1F 63 0A 28 08 E2 C8 9A 05 D4
 4B BD 5B 70 EB 46 68 42 5D 43 39 CC 1B EC 5E A4
 0F 05 FB 66 DC F2 65 52 B8 2C 6E 99 43 C0 71 03
 FC 10 E4 F8 31 CC 2B FD B7 0D A0 4F 8B 78 23 5E
 D9 66 60 97 2B 14 C7 07 AB 48 33 79 35 31 60 6D
 38 66 D0 C8 92 44 54 E8 F0 DB B4 37 D0 2D 30 78
 F1 B1 C1 6B 24 33 25 FE AE C9 B8 D6 34 9D 16 1D
 CA 98 E3 02 8D 3A 97 5C 72 E0 8B CF F3 4A F1 59
 DB F7 5C 8F CE 3D 15 22 0A FF 5B 53 68 04 24 12
 C9 39 24 C2 E1 37 03 09 66 EF 8D 4F BC 9E 20 D7
 5D F3 52 D3 C8 F6 87 85 94 26 6F 66 91 F2 2D 5A
 E7 77 7F 13 CA 05 71 B4 7C 13 88 20 6C 32 95 D2
 AB E2 93 CE 6C E2 9A 4A 56 A9 C7 E4 6D 09 DC 17
 B5 AB 47 10 2A 36 05 90 BC 1A 51 43 75 DC 48 D7
 EE F2 AE 7B 80 52 A3 D3 3A 66 A8 86 0A 0E 1A 19
 81 5A 9D 5D 93 0C 8D 58 C4 E7 32 11 5B 87 21 C2
 01 7D 6B 36 02 79 A8 7A 47 F7 98 3B 0B 51 96 98
 B3 23 2C EC F7 98 BF E6 FB 10 8C 91 DD 99 19 AB
 12 0D 99 F1 22 0E 8B 7E 81 B4 42 57 A6 44 B4 9A
 E8 3D 9D CD 75 B2 A1 23 FB B2 6F 43 7D D6 BB 0F
 CF 91 66 F1 7E BE B2 D7 CA 22 18 43 66 5F A3 48
 9A AC 99 D8 44 2B 99 8A 03 D6 85 BF FA BA 5B AF
 CB 98 1F A6 C9 3B F7 2C A3 E1 5F 5D 80 2E 40 02
 F2 1F E4 6E DA B1 DD 34 CB 9A 96 CF B5 31 76 98
 23 1A 4A B0 0F E4 D1 1F 71 14 51 6E 88 70 E0 F7
 D4 14 39 EF 7F 1F FB 83 1B 89 76 CF 39 3B E0 CE
 5C 95 AE D5 38 CC F8 AE A1 C4 DB FA 45 E6 0B 5A
 59 6F DF 88 CC B4 71 7E C8 75 FB 27 5A 5A F2 19
 E7 45 6B F8 41 ED D8 88 E3 FE 58 95 9E B5 84 7E
 20 A9 36 72 C6 5A B3 A2 49 87 90 D6 AC 72 21 87
 08 71 4A 34 EA 5D B7 F5 5A 42 82 EE C5 1A 5A A0
 06 02 12 27 6B 19 B4 4B D7 D1 A3 1B 42 0B ED 87
 4E 5C 85 E7 4F C1 DC A5 B7 AF ED 81 03 B6 48 AF
 1F 8F FC 29 ED 02 A2 7F 83 09 6B 8F 9B C9 1B 7F
 FD 62 52 88 2E C1 23 70 E2 84 4B 9D B0 E5 A7 33
 1F 9F 7C 11 1E 5B 5B 40 7D B3 4E E5 2C 1F 9E 44
 8B 87 71 A0 E9 F4 AF 06 F2 63 78 AD 3E BF 5F AF
 D3 87 C9 AB B7 01 EC E8 93 61 36 C2 57 D2 0D D1
 69 DC FE 67 D7 65 CA BA 8F B2 63 0E D5 7D D0 91
 3C 25 6A C7 9E 75 03 CD DF D2 CF 1C 77 47 8E D5
 B6 BD 9F 2F 6B 7A 7D 99 B8 F1 FF E8 FE 0E BC 10
 62 87 A9 44 27 4B 43 66 E6 4A F3 5E 1F 08 6E 6A
 03 0A 3C F3 B9 3C 1D 4A 03 D5 73 DA AF BC BA 0F
 3A 84 6B AE 69 0F 11 91 56 C6 56 36 A1 13 81 A7
 12 6E 78 FD 48 AD 19 2C A5 5D E2 6C 09 67 1B 49
 29 6D D8 16 0E 4A 1C 1E AC 6A 50 F4 E2 29 99 75
 8D AD B6 73 65 C5 7F 53 35 14 1E 7E C7 FB CB 23
 3E D0 40 BD FC 01 2E 99 55 A7 1E 9B 2D 1C A5 BE
 4E 2A 7C C5 7E AB 25 8C CB 7C FB 46 BE 02 45 1C
 7B D4 54 78 F5 FC E3 51 14 8B 5F 05 7E 76 B1 2C
 14 A5 4B 4E BC B0 E2 B2 54 C3 AB 44 17 96 C0 21
 6B 83 FD CD 3C 2D CF A2 BF B7 8E CD 46 37 F9 F5
 79 EF 5B BF 4A C0 FC 4A 4F 15 7A B3 3B AD DA A9
 51 AC 6C 7C C6 8C 6D 70 9F BB 73 C2 51 08 E5 AD
 87 3F B3 1B 7D 64 B6 BD 67 AB A2 02 F3 A4 3F 08
 DD A5 9A E5 D6 8E 9D C6 C4 67 22 A4 AF 7D 06 C2
 3F 95 A4 F7 79 33 DF EA A9 0D 30 AB 60 58 DA F3
 4C F7 83 F2 EB 53 64 9C 30 11 10 B2 25 5D C2 B0
 C0 89 19 C4 54 8E EC 06 56 1C AC 5F B8 FF B2 DD
 AD 30 22 98 0A D5 E4 9C 86 41 70 F8 84 1D F1 C0
 37 D5 55 B1 BF 86 55 36 E4 6F 4A 4B C5 10 CD 69
 19 9E 63 36 49 80 7A C8 52 3D A0 FB AB 8F 4A C0
 62 BF 5A 25 82 22 9C 6B BC B1 F7 C9 CC 0B 20 6E
 0B 17 6D 12 18 A7 02 2C 49 FC A5 B3 FD 55 B2 E6
 25 3C 6F 5F 21 67 9C 98 90 27 C6 2C 04 D2 93 F1
 5D 0E 00 76 0C EE 53 89 B4 AB C6 06 E4 46 B3 F3
 A1 37 BC 4C FF 03 E2 55 80 51 7F 2A CB 94 0C C1
 16 37 51 2F A6 F9 2C 3A 93 1F 97 AC F4 6B 15 01
 C4 22 B5 CA 2E AB 8C B1 A1 46 27 68 00 1C AF 38
 9A BA 7C DF E2 EA BA FA E9 A2 0C B0 C3 30 D2 22
 5E E4 8B CE 8F E3 A8 0D 7B A0 DB 42 50 CB DA 19
 89 D3 23 2E 12 D9 36 A4 56 81 25 7B 6A 6F D0 1F
 25 29 0E A9 18 3F EC A7 F6 1B EC 3A 05 6D 8A 46
 BC 9D 58 DD 83 41 E5 40 76 4A C3 65 61 AD AA BE
 F8 EB F7 4E E9 38 3E E8 53 12 BA D7 D6 A3 BA A9
 17 63 3E 74 DB BA A4 D5 74 18 05 AB 35 50 60 32
 99 8A D8 4E 87 AA 84 A7 22 74 28 C2 73 96 53 5E
 09 F9 BF 2D 6F B8 9B 75 F6 1C 6A 6E C3 E3 CD 7D
 6C 81 91 AD CA 14 D5 F4 DE 1F 19 F3 F2 D8 FA AE
 5C 3C DB 27 96 96 A0 AB 3F 62 12 AE C7 2F 90 7C
 BE 50 73 92 E7 2F D6 03 14 67 82 AE 5B FC 07 1C
 16 5C E8 A9 AD 1C 88 6C 20 94 1F AA 10 C9 9F 2E
 35 34 C4 9E 30 D4 B5 01 EF 2B 6A 00 36 EE F0 05
 27 64 86 CF E5 15 99 AD CB 5B EF 2C 81 78 B2 E3
 5A AC 74 DC 38 F9 2F 92 71 29 82 03 0B 2E 27 4A
 F3 38 82 3C 59 75 93 34 F6 98 4D 3B 41 68 FF 24
 DD F3 5D 07 72 FB 30 BE 21 33 BD 1D AC 3C 13 F3
 2C 09 A4 4F 33 43 13 1B A0 A7 FC A9 5D 6C DC B7
 D5 0D B9 32 5A 9A 74 95 D5 0E 41 4E 5B 00 3A FB
 30 C7 60 87 BE 90 28 22 65 52 6A AA 82 6E 50 4C
 6A 3F EF 47 6C 18 96 E0 2D F9 A9 31 20 2B 7F A3
 DD C1 D0 B9 62 B7 F0 2A FB F8 A3 CB 31 10 CC D3
 D8 DB 7E F1 1C EE 85 88 33 F9 BF 13 E8 BA DC A8
 76 40 14 53 A4 E5 6F 2A 63 45 5F B6 2A 91 8D 9C
 E2 66 3A 56 0F E5 3B CA 2B 2A D5 11 CE 69 FF 9F
 FD 63 49 16 9E 89 BA 46 21 E2 19 96 23 3F 8C 56
 1F 50 57 03 DF EE 25 0D 48 80 78 EC 90 3A 2F 3E
 E5 7D 47 EA 5A 59 BE 5E DC C5 C1 22 42 CA 4A A2
 54 43 A4 D8 4E A4 7D 3C D6 81 01 6A EA 45 B6 D7
 3C 4D CE C8 0D B5 9E 3E 4D 23 81 83 8B 35 4C 01
 92 DD 6F 7D BD 58 BE 96 84 6F CB 1B 4E ED 25 C7
 A9 4F 8F C7 75 AB E6 A3 5B CB E2 AE 3A 0E 1D C8
 A9 57 97 A6 48 F2 C1 CE 9C 41 E7 F5 B5 30 7D 47
 1A B0 CD A8 26 6C 93 C4 EA 29 DF EB CC D8 FD F8
 9B FA 93 5F 00 13 40 A0 02 4C 7B 00 03 39 A2 CF
 E6 5A 11 2D 39 F0 62 96 18 5B EE 72 D0 B0 FB 19
 F9 4E 85 27 DC EE 44 A3 53 27 EE A8 A7 04 4A D9
 61 C1 7B ED 75 90 04 F8 28 66 3C 0F 50 72 3F 85
 CF 33 33 D3 66 36 BC D5 F1 50 30 F2 CE C5 22 BC
 18 A5 4B FC D4 54 FD 0D 5E 1C C7 7A 8C 68 78 E2
 3C 53 7A A1 37 BC F4 3D CB E3 8C 74 F3 5C 2C 73
 F3 57 E2 3B CF 78 BD E4 3E 47 D4 0D DF 8A FA 26
 0C B9 98 88 AF 6E A3 51 75 55 EC AF C4 25 3D CE
 CE 31 35 BD 8C CA CA 99 D2 0F 21 02 B1 BF DE BE
 71 8A 15 59 BE 36 63 87 5D FE AF CE 46 2A B8 AC
 4F FC A4 6F D6 28 75 4B 89 9B 2E CA 94 91 5F C7
 F2 08 76 E1 D6 64 C4 55 7F DE B5 8F 0F A7 F0 3B
 EB 06 8C DE 57 68 99 A8 50 0D 82 08 B5 6E B3 97
 66 C9 8E 54 A1 79 67 FE 73 2A FD 4A 79 8F 60 B2
 F6 BE B8 80 DC 13 C8 38 6C F9 48 FC 49 80 62 25
 AE FB 33 80 31 AC 58 C5 58 E2 BB 9B 6C F0 55 BE
 A9 CE 25 BA C5 DE 4F 77 B9 5A 2E 9A C3 C8 03 65
 81 DF 2F 05 B7 5D 6D 77 D6 D2 5F 45 55 B3 39 FC
 B4 62 45 78 A7 CE C3 51 96 50 DC 34 F7 EE AC 3A
 8A 0A C7 8B 0F 7F 9A 7D 60 92 4E 95 77 BC C5 36
 74 71 DF F9 E4 C6 16 A0 7A EB 77 4D A3 8C 54 FF
 3E 4B 2E F3 11 07 A3 3A C5 25 3E 5A DF 5B 86 05
 25 58 56 A9 F1 0D 2B AC D7 22 17 33 22 E7 8B 02
 3E CD 40 BA 32 4F 73 E2 A6 97 6E 26 D7 67 7E 0E
 25 C4 8D A8 01 39 0C 99 7A FC D4 33 C2 E6 94 1D
 32 BB 4D 46 CE 17 3B 82 74 6D 46 14 BA 1B 6F E4
 B5 46 6D 9F FF A5 77 D3 D6 E0 19 43 96 97 BB 8B
 5D 30 3F 4D 70 7D E6 C9 1D B8 E4 E9 05 1B 93 69
 AB A7 28 41 62 95 AE F7 79 12 17 9B 7F 93 C3 FC
 77 58 9C CF F2 38 76 D6 73 CB 2B BF BB EB B8 6F
 77 AF 0A 50 4F 89 C1 5D D7 5E F1 96 7E CF D0 6A
 B7 9A B9 C6 05 4B E2 83 DB 7B 76 2F F3 1C 65 5C
 EE 76 A8 85 E6 27 93 32 6D 8A D1 AC 0A 89 B9 9A
 61 CA 46 E1 9D 43 0C 9B 74 34 D8 59 59 CF 5C 80
 92 51 E7 DD C1 98 15 91 80 67 C1 13 3C D7 0E 14
 07 BC F5 5E 68 16 82 C6 3E E5 C6 D4 1A 08 28 B6
 58 7D 9D DB 8E 11 73 39 5E 14 40 7F 1A 81 51 7F
 81 68 4F 77 B8 C4 CE 4B 48 64 B8 E3 B4 65 3D 44
 D7 AB 80 21 F1 3C 93 D9 9A E8 78 87 71 DA 85 D1
 72 CD 51 DA C3 7B 71 D2 D3 73 BE 22 19 FC 3B 81
 A8 88 A5 D3 25 D9 0F C5 7A 16 AF F1 D7 DE A0 6B
 B3 83 FF 46 E9 C4 CD D1 5E 0A 26 8C E3 7E FB 0F
 0F B8 43 C4 D2 E9 8E 53 07 7F 4E 62 C8 EC 5C 5A
 1D 0C 8F 19 AC 26 0B DE 04 8E 4E 97 00 9F 7C 3E
 EB A5 98 7E 00 29 75 2A E9 6A 7A 69 3F 51 64 ED
 25 B8 FA 53 4B B5 12 97 4A 04 9C CC 24 3F 3D C0
 55 4D 18 D6 3D D9 B8 4F A1 CB B6 9A 49 6C 67 5A
 9F 35 14 6E BD 9D 84 B7 9B 8D 9B 51 E0 FA 33 E8
 52 40 FE 3D 34 EB 4E B8 E4 73 5D 9E D7 8E 43 56
 42 F8 4D 0B 33 17 FC 98 41 36 42 76 DA 89 BA 63
 3C 1E 9B 2F 42 0C CE EE C6 8E FA 12 30 5C 01 CD
 C9 03 1C 73 EF 24 07 7C 1D D9 DD A4 E2 95 00 63
 C9 64 24 82 26 16 25 D3 40 98 20 B1 BC 18 D3 30
 D5 5D 93 9F 35 B2 DC 17 83 4F D3 09 9B 2A 92 58
 FD 5B 93 43 2C 45 A8 50 02 80 07 D2 32 20 F8 B1
 EF 70 8E 0D 7E 97 75 1B 59 E4 CD 9D F9 74 FC 7A
 7E FC EB B3 C8 A0 E9 31 B5 94 6D FA 5E 9A 59 6D
 74 1B 9B 77 1B CA 9B 6F 1C 90 AF BE 7E 7B 38 FF
 49 B1 43 B5 16 B0 66 EE 10 3E 5F D9 D8 14 E5 F7
 80 DA 0C E7 DD 76 B7 AA BD 66 13 68 B6 0C 02 16
 08 3C B1 EE 35 08 1F 25 D9 67 51 68 3B CE 2F F5
 39 5E E7 18 52 D2 54 F4 E5 0E 2F C8 90 04 52 65
 0A 4E F8 A9 E5 ED 92 FB ED F7 61 A4 F0 6C 68 81
 D4 89 CA 32 3E 31 45 63 30 4E 2C CA D9 3E 86 03
 14 ED 0D DF E5 AF 60 91 7E 3B 14 3F 89 59 99 4E
 FB 88 AA BB 58 D1 AE 6A C7 52 C0 34 AC 08 13 19
 30 4D 84 A8 BA 9D 15 8B 69 AC FB B8 7C 3E 56 01
 F9 E8 9F 13 F0 6C DC F0 DA D5 3C AB 79 98 29 FA
 BA 33 85 7C 79 8A 5D 5D 7E A4 58 1E A0 3E 82 E1
 6D E0 5D 1B 67 2D 56 41 71 8E 99 04 E8 4A B9 B4
 6B FE 1F 6B 3D 20 BE 9C 72 A4 12 A2 0F E5 D6 9B
 AB E6 88 28 65 94 BF BF 6D D3 EC 54 FC 3D A3 EA
 B0 E0 F2 16 05 A6 24 26 FC 99 77 C4 65 92 34 00
 D3 38 69 4C 76 D4 4D 4D 01 19 8F CB 25 3C 50 EF
 64 9C 39 7E 54 24 9C 97 F8 95 94 9A 0C D3 C9 EE
 4B 64 81 A0 2E 69 34 39 A3 04 7D C4 1F D0 9B 4D
 2E E6 80 85 51 62 19 70 6D 10 EF 5D 72 5F 8A 5D
 45 41 CD CD 8E 99 FF E7 7B 6C 44 22 18 95 78 BD
 A2 06 CC C5 50 31 B6 57 F1 4B 71 CB 61 9D 15 6B
 B8 3A E0 18 CB 5F BA 51 99 32 B2 44 FF D7 5F 67
 B9 BA BC E5 98 CE DD E2 83 B0 AA 46 79 FA 08 A4
 7B F4 1F 19 0D B6 CB 4B BB 67 17 FB 4E 5B 6D 1D
 02 C2 F5 0D A2 60 F1 45 AB 0C D0 F8 30 2A 73 C0
 3E E6 7B 3E 5C A3 4B F0 7F 36 36 4B 79 76 D4 13
 89 5D AF 90 02 9D DD 16 0E C5 28 1A C4 AE 01 D7
 C1 EA 4A E7 A6 74 5A CA 36 85 07 CE 70 29 87 14
 0D 6B 88 72 C8 6C 21 60 AF 85 0B 4B CC 3E CF 3A
 32 0C C2 8E 3C E5 74 32 FA 4C D2 B8 44 37 79 63
 01 26 37 6D F3 DD BC A3 52 CB DF E9 A5 03 50 2F
 EB B4 77 8E 0C 09 07 38 87 2B 97 4F 86 71 C2 57
 D9 8C E8 C9 42 AC 60 56 67 5A E2 0E 68 89 CD 41
 51 2B 79 45 E2 45 0B 19 F4 A5 05 72 B5 AB 07 A4
 ED 5E 80 36 AD 42 C7 F6 BC 92 BF 65 4C FB B7 21
 7E 65 BD C5 70 2B 7D 6A E7 80 24 FF CD 89 38 F0
 06 F5 65 9F 29 57 D8 FC C8 DD 5A 26 FC 0C D8 4D
 BB D8 BC BB 09 B6 9E 08 6D 36 4D 8A 52 6A 1C A3
 F8 59 6F 0B 00 E6 A8 C2 2F 3A AE B3 97 17 8B 77
 8F AD 7F 01 C0 06 72 A6 C9 E2 35 65 4A 15 93 95
 B7 64 E2 03 FD 5F DD DE A7 EE 7C FA DA 3E 83 01
 FF 47 85 93 9F 8A B8 12 5A 33 6F 14 71 4F EF A8
 A5 3A 83 EE 33 B6 FA 16 49 CC B9 12 02 85 6D 63
 78 C8 74 70 48 E0 A7 14 B0 0C 8F 3F 94 D5 83 09
 19 CB 29 07 F6 F0 48 FA C7 D0 22 69 B5 AE 2E 1F
 A3 81 C4 43 29 D4 F4 2F 61 8E 6B 1E 85 89 C0 C7
 5B F6 92 F4 CD 2F 6C 8D 05 BB 52 B7 4B 46 46 7D
 26 AB 64 F8 49 A1 5A 19 A8 D3 E9 72 2E 07 F6 BA
 33 2C 73 56 0F 06 EA 56 FC 55 E5 A1 85 84 AD E2
 FE A4 BC 9B D9 0B 72 6F 09 44 42 EA A3 DC B9 40
 40 FD A2 D7 82 0E 86 77 FE 3F 8D E3 0A ED 85 09
 1D FE F7 3D 12 9F 45 20 B6 A5 FD D6 0E A8 92 53
 66 D1 03 69 0D 9B D9 CD 45 3F AF B7 C7 A6 67 B2
 1B 43 FE 3F 92 E6 CA B0 95 7C 05 3C B1 4D 81 24
 36 10 EA 50 43 EE 90 CE 5B 7E 04 7E B3 77 F8 90
 DC D9 47 2B 11 4F 88 1C 70 20 D5 F8 75 2C 5E 0D
 5A 5A E2 8A 56 CC 5D 56 B7 41 66 74 63 38 EF 34
 49 8E F5 F1 E2 D5 49 BF E3 1C B3 1B 95 90 F7 FD
 42 55 85 10 E2 2C B1 23 FB A1 D0 32 BB CB AC 4D
 E9 9F 46 A5 D9 23 A3 26 D9 34 B2 D1 BE E3 19 4D
 EE 7C EF CE 06 27 CB E4 67 49 DF 7A B4 0F 3C 50
 D3 26 BA 30 A0 1D DA 09 37 9D 81 86 0D 9D BF 3A
 EF 17 2B AD 2C B2 FB 76 BE 59 94 6F 65 D9 00 ED
 A7 4D 1A 90 2E DC EC D7 ED 50 FA 58 55 CC E1 3C
 C3 F4 5A B7 D1 A5 53 BA 0D 3B 0C F3 75 C8 C9 D4
 95 87 9A 6C 60 4B AD 19 98 54 FF 2D 9B AE 10 EC
 F6 1E 29 F8 0F 3D 8A 3D 72 72 80 1A 9F 2F 64 3D
 C7 42 E4 E1 BB 2A F5 56 C8 CF 23 68 5B DB 02 59
 FE 99 D5 CA 09 6C 6A 1E F2 F6 F8 15 8D 98 47 25
 C0 C1 E1 CE D8 BF 77 04 F9 D5 7B 58 E9 ED 7F CA
 01 79 B2 88 9F CC A2 4A E1 8F 43 76 C6 80 EC E2
 15 CB F8 B2 8C B0 15 5D EE D6 DD E4 B4 43 A2 4A
 A0 82 71 F8 FC 38 5C 22 44 B7 D6 98 BE 3A FC E9
 91 E2 AD 35 17 C8 AC 09 F3 20 D4 77 F7 C9 FF 68
 65 B5 21 E5 37 7A 9D 87 A3 24 14 F5 A9 22 67 56
 6F 61 76 FB F2 36 81 D6 6B 50 24 4A 30 42 08 1A
 5D 72 B4 7D 93 B9 09 6A DC 6D 9E AE E0 C9 A0 BE
 18 73 1B 5F 3A A5 90 0F 55 83 FB B1 33 68 C7 11
 34 3D CB 20 45 42 46 ED 6F 15 F2 C3 0A C7 A2 CD
 63 50 2A AF 7C 66 19 7F D3 71 37 F7 E2 BB 94 44
 C2 C3 0E C8 7B 2C A3 C3 40 A0 A3 E0 C8 CD 47 54
 D7 1F AE 44 6E 14 6F 9C F3 29 5D DF 6B 87 82 FF
 F5 76 6C 7B C3 B6 8C 2B 80 75 98 87 CF F1 91 49
 F1 2F C7 6B 52 DC 71 19 DE 6C 5E E2 16 DF C1 61
 B8 7D 63 B4 2D 6A BB 03 CE D0 52 1D FB 1A 2E 16
 B3 04 E4 BE 92 B0 6A 16 B0 64 6E B3 D3 41 36 3E
 DE 41 D1 1C B7 CF D5 E9 CE 68 80 9B 83 C1 51 CD
 70 E5 06 44 F1 C0 0A 8A 48 74 B8 8A 01 F4 64 38
 0E 25 7E 57 AB E3 B7 62 CB 20 44 AE FB 7F 17 46
 F0 CE 60 B5 B0 F6 97 C6 D3 F2 9A 0C 2D D0 D2 30
 14 14 1A D9 C9 E6 9F 8F 22 84 45 A8 8D D7 48 06
 DF FB 63 D7 F1 6B FD 55 56 93 A0 DB E0 4D AB E1
 71 EB FC E6 D5 AC 77 D6 8C C9 D9 B3 C5 54 16 1E
 87 29 7B 81 95 C4 AF DC CE 51 E2 28 19 CC E4 0C
 E4 EE D2 FB 26 1A 5A FD 9E FE DE 22 C5 4E D1 A4
 67 03 D0 4E 51 8B 61 1D 21 A0 8A 82 65 7E 2E 38
 88 9E 62 C3 7E E9 0B 90 64 A2 35 E1 AF AE 08 78
 C3 40 65 BA DC 7F 0E 93 D1 A2 1B 6F 75 5D 8A 41
 22 DF 46 FB D0 0A 1A 9B C9 1E 7B 4E 10 C5 92 D5
 40 A2 19 4D 63 8E 9C F0 60 D6 27 9B D7 06 15 21
 FC 3C 82 90 A3 04 32 3C 9F 06 8D D2 E1 5A 1C C6
 64 47 00 01 E0 EF 28 D5 5B 5A CE 71 CE 83 FD EE
 DD 15 D6 4A DA 15 B6 58 C3 FB 47 BF 70 5B 5C C2
 54 4D 2F 47 98 29 AE 2B 4C CD BD FA 5B 30 7E 60
 D9 32 C6 2A A2 45 7C 68 87 8A 40 05 3F 29 F5 B3
 FE 41 28 6A 43 35 06 62 29 3E FF 7D 0E D4 5E 94
 C2 77 F7 D6 C7 08 01 62 7F AC 04 F7 BE 9D FD 49
 09 D3 98 B2 B6 9A B9 E5 20 A0 D0 19 D1 3D E4 62
 BA 14 43 7A 2F 12 0F D6 2E B2 A2 D1 42 70 DE EA
 85 65 E9 1E 8A E3 25 EB 7D EC E1 B6 16 9E B0 BE
 F3 28 72 A3 72 58 E6 B1 AB 93 A2 05 CC FD DE 42
 7A 86 C7 B9 35 FE 75 B7 9E 94 79 7C B6 0A 60 4E
 34 BC 71 52 51 14 3A 6F 55 CA D9 06 4C 9B 15 1C
 E2 FF 90 30 FC 02 7E F5 1D 8F 7B 8F C5 CB DB 7E
 1B B3 75 2D 26 63 F1 B5 61 7F 92 E7 39 0D 45 C5
 C1 E6 62 FF EE 4C 85 0A B5 AE C6 7D BC 98 C2 8F
 A0 C0 2B F2 A3 D7 C8 76 8C 4B BC F1 E3 FE C3 7E
 84 B7 86 2A C5 A7 8C 01 36 99 00 D4 23 E1 96 5E
 79 B0 9A BF 8A 77 CE DB 32 8D EB C9 EE 43 BF C4
 7D CB DE B1 5A B6 BD 71 94 1B 80 B9 81 09 AD 81
 AE 83 F9 DC 05 D9 E6 E0 00 C9 4B C9 CF A4 C0 AB
 C9 91 1F FB 2C 63 26 C8 DC 82 FC 3B 71 BD F2 7D
 56 AB 45 DB 48 07 F8 8F CD 5F BE 08 DC E5 17 1D
 83 3F D4 58 AB E0 09 ED B8 DA 98 09 F7 D1 1A A4
 68 20 46 F7 81 F4 69 67 D3 D6 F6 8D 6F 41 6F 8D
 F2 3C 40 DE F1 BC 6D B9 9D 6A E3 EC 11 B6 95 5B
 E3 F8 A8 7B 02 4B 43 24 EF F0 B1 E0 98 42 19 4D
 F2 98 71 F7 47 3D 75 E7 0D CE F2 08 91 27 CE 5B
 33 9D D9 B6 D1 3C 15 4F 26 E3 B8 BC C3 B9 6C FF
 25 63 B0 F9 56 EC 37 D7 FE D9 DF 11 04 72 41 A9
 AD 68 80 76 00 A8 7B 9E 90 13 A9 F1 B1 B6 73 67
 8D 01 66 D2 A4 E2 06 D6 F2 8E 8F 92 92 D1 8F 06
 70 56 58 C9 AD B1 1D 81 EB DD 0D 18 64 28 B5 08
 F1 14 0B B7 FA 57 29 14 74 7D CB 68 CF EE 76 89
 F0 50 EA 34 E9 6A 4D 7D 56 4C 63 B6 F8 EA 01 48
 A7 C6 39 36 01 BA 5A FC B7 A2 C9 E0 02 A3 7B 22
 6A D2 96 5C 7C CD 41 60 E2 AD C7 23 33 36 B6 D6
 A2 9A BD 6B 3C 7D 8C 76 B7 85 0E 25 B0 B0 26 43
 EF 60 8D DB 6D 02 C7 3F 13 97 F3 4E F0 57 32 5A
 A8 FC 42 C2 14 BC BF 6E 67 AC B6 0E 59 57 A1 90
 E5 25 80 1F 3F 67 51 58 37 13 CB A2 D5 4C C9 56
 11 0E 34 38 32 AE DB 53 D3 71 4A 2D F9 C4 21 49
 B2 41 89 5A 71 5A C6 CF 00 41 BC F6 F6 6E A5 26
 30 96 35 CE F8 60 D7 B0 33 B5 A5 76 14 0D 85 2F
 30 33 EF 3F C0 C7 CC 06 7A DA B0 77 5E CB 87 BF
 97 FE CF 19 1C FB 34 64 72 67 7B 6B A1 D4 11 3A
 07 18 A1 6E 17 BD 98 9F 94 7B 1B C5 6A 8C C6 D8
 1A 23 0B 67 12 CB 7E 08 18 F1 DD B4 AC 08 6A AB
 02 D5 FF 48 53 A5 4B E6 D7 BB 5D 46 C2 62 4D BF
 9E C5 34 C7 0F 40 8E B9 B7 3E 57 A1 97 A8 99 95
 CD ED 53 4C B4 56 AB 6B 41 16 FA 9C 85 08 73 FE
 D6 28 29 C5 0E 5D 06 5A 08 A2 95 F3 80 BF 3C 3B
 90 BA 93 C8 10 73 AF 6A 7E 7E D6 EF 5B 16 AA B7
 70 97 5A 03 92 C4 96 FD B5 1D 43 CC A7 A9 1D 51
 B0 55 25 B3 EA 07 26 E8 6C D0 52 67 DD AD C6 D8
 9E E9 BD E3 5D E4 16 8E 41 C6 CC 07 4E 56 D8 E1
 AA CB 9D 6A B1 55 7D C4 5C 5F 06 F9 C1 63 8C 23
 92 34 2D 79 E0 32 9A 0E 7E 8A E2 B6 99 42 6F 24
 92 14 50 32 EA 17 01 50 FF 15 B5 FF 74 DE 8D AA
 04 7B EF A4 57 19 42 DF 22 AF AF 18 B4 89 8C D0
 86 A1 85 36 ED BA 85 07 F7 93 56 AD 79 16 CD C0
 E4 AF 83 F8 42 96 51 E3 37 EA 64 ED A6 3F 58 DE
 9C 63 54 87 47 70 3A 1A 5B 75 DF 30 E3 E1 84 A4
 05 BC 38 A5 33 45 96 04 35 87 71 7E 9D A9 E6 A1
 0D FE 0E C5 E2 67 19 77 EA B2 39 C0 2F FA 50 19
 B4 27 5A F0 D2 94 9B 70 0D 23 95 4E EE D1 9A A2
 FB 03 72 67 FF 85 90 11 19 DB DF 81 2A 9A 7D F6
 65 19 28 F4 CA 5A F5 88 E5 EB B2 C4 59 99 32 63
 16 5A C6 A3 71 08 48 35 40 2A 83 EC 9B DF 62 8A
 DA 12 9C C3 0F 83 1B 3A 3E 9D C9 55 49 79 AA D8
 AD E8 FC 5E B1 FF A8 D6 CE DD 65 43 85 6F DC 07
 38 74 E0 97 6C 11 CB D3 33 E8 18 B2 89 8D 2C 9E
 34 9A 86 B0 B4 DB 80 5B 0A 16 3A 1E E7 81 06 45
 11 D7 DC D6 E5 F7 3C A6 9E 64 57 A3 44 45 F3 3E
 55 FD F3 7C 1E 96 9C EE AA 59 5E 2C FB 22 16 C4
 75 12 B8 87 59 47 A6 74 0C CA AC B2 4D BE 1C 96
 D4 A7 0C 7A BD DC FF ED 9D 26 2D 73 AD 8C 59 E1
 14 45 86 10 33 C2 CA C5 88 7B DC C7 ED E1 51 91
 B7 B0 3D D1 78 12 2E A6 7E C3 EC 0E 9A 1D 8D 81
 05 CB BA 45 3F 17 1B C5 5D 35 52 2E A3 DF DB 14
 9D 4D C6 1D 36 73 6A EC 79 6D D1 6D 84 14 43 82
 7D 04 1A 2D 2B 87 04 40 D2 34 42 B6 FC 56 49 9D
 85 8E F7 8F F2 DA 15 C7 76 0D 4B 13 98 BA 8D B0
 BE 0C 40 C0 50 F4 BA 0A 25 CC B6 C4 3C DA 5A EC
 C9 34 CA D8 5A E8 3E CF 0E 65 25 47 4E D2 6B C7
 8C 39 71 F7 BA 65 54 B7 B8 F7 02 1E BA BC 81 09
 32 B5 D6 B3 11 0A 23 44 ED 0C CB 18 C8 3D BE 2E
 4B 7E 3C E0 22 9A F2 A1 57 AC F3 29 23 2C A5 66
 CF 87 28 A3 51 4D B5 F3 3B 8C 3B 8B CE E5 3B 49
 62 FF AD C0 80 0F CE E3 9F CB 38 65 B9 5D A0 2C
 35 16 4C 4B 0D FD B1 AD 77 AB 5E 8D FA 25 9C 42
 92 A4 94 8F 27 47 C9 9C E5 7C 15 4F 04 E6 16 8C
 2A EC 29 E2 A2 E2 25 2B F6 03 66 6C 2D 5E 9F A4
 A4 62 9A B9 B2 82 A9 A0 BB 9A 0C 46 BF 04 0B 4F
 24 38 2E B7 FA E5 92 19 3F 9F 0C 0E 88 16 46 52
 B6 97 68 FA FD BC 04 85 82 CB 38 82 BA C4 69 2F
 C8 A5 ED 54 E0 72 AE 39 04 F8 6C 1D C8 27 7E B4
 7C 31 F0 D0 50 AF 05 BC 60 CC 04 D5 4F 25 80 E1
 E9 D5 CD E1 54 FC FE 47 D7 4F A4 43 EA DE 53 58
 A8 4E 63 10 B7 E3 09 C2 BB CE AB 2F EA F0 76 FE
 BC 36 33 65 67 62 25 03 04 EF 8B F2 B0 E6 47 58
 51 33 1B BF 97 A0 D4 08 B0 5C C0 EE 2C E2 14 83
 E3 7E 00 74 BD C4 B1 96 79 BC 7C 2E 30 2E 2B 07
 36 80 48 47 AC 45 A1 27 23 0A 96 D0 D9 EB FF 8A
 23 B7 01 DC 05 3D 8D A7 83 29 A6 5E B4 D6 41 D2
 A2 AC B8 78 6D 84 0A 22 2F 3F 65 ED 1B AC 79 CB
 ED CA 18 6C 6A 19 69 40 84 7C 1C 2B 45 0B C1 89
 BE 8B 96 94 5B 9C 47 68 EE 30 F6 A8 BF CF B8 D1
 29 F0 99 14 6D 43 EC 37 32 F9 4B 48 C2 E7 0A 3B
 1D 86 E0 D5 AA B9 D1 6E 35 33 DA E6 BF EB 5E 59
 6C A9 64 39 5F 35 0C 5C AE 44 0B B7 3B E7 F0 51
 0B AE 09 49 AA 6B FA CA F0 1B 71 8D 49 BD C6 49
 36 7C C6 C2 14 D4 BE 99 57 7B 6F B0 6B F9 82 23
 DF A2 D4 4C D2 3E 57 57 E8 98 37 69 BF 14 57 32
 19 DB DA 3E 01 B5 AF B0 74 7B C1 86 26 B7 2B A5
 A8 CF 25 32 F1 FB EB B8 76 6E 1C 95 C2 D2 0F 1E
 C3 E6 02 43 79 AD 5C 25 E9 06 DA 5D 40 57 36 8F
 DB A5 C9 BE EF 4C 09 5E 91 B1 01 6D 0F 57 95 C9
 C8 30 B6 27 6E 16 4F 16 4C 52 92 8A 02 1C 36 13
 C0 E6 95 EA 7F 29 AB FE BB 12 F4 57 3D F2 EA 87
 CF C3 FE C3 65 A5 59 A0 27 39 94 EB 9F 89 B1 72
 09 D2 CC F0 46 A6 3C FA 79 0C 93 9F 6A 5C 72 72
 13 DE D3 A8 FE 26 A1 20 44 80 38 7E B9 CF DC 20
 B4 2C AB 8F 5D 31 03 81 82 AE 3D 5E 12 83 EC CF
 D5 40 2E 5B 50 BA 4A 63 76 14 9F C7 7F F8 84 0E
 93 59 DF CA 48 53 12 67 4F 0D 87 6F 2B 6F 95 40
 1C 47 F9 61 85 B8 A4 C5 CA CF 1D 65 CF 4B 93 6A
 39 FB A5 37 42 02 51 FF 7A 39 8A 30 7D 86 84 26
 55 63 88 6B 08 A0 54 86 B9 90 64 02 CB 67 7B D2
 D4 D7 61 D0 2D 7E CA 72 3D 8B 03 ED 16 92 83 B9
 2F 32 BF 51 23 85 03 1A 29 C7 E2 46 EF 9C 73 86
 EF 2A 6F C9 6F 7C 98 54 58 A6 BE CF 03 CC 5A 85
 72 1A A5 AF 64 FE 23 F1 F7 4A 28 B4 63 07 D1 5F
 BA 47 05 5E AC 40 81 D8 53 7E 33 69 FE C6 93 8F
 1C 17 F6 AE A5 FB 4F D9 20 77 32 83 7F B3 18 23
 6F A3 C8 87 BF A1 9D 0B 8B C2 B1 D2 80 73 BA A7
 32 11 9D 7D 42 0E CB A4 84 B4 DB 56 D5 44 E8 3B
 8F 20 81 1E A2 1D 79 41 35 BC A6 1A D2 95 92 67
 89 31 24 7B BA 6C A6 B9 09 6A E6 AB 91 98 A1 24
 63 6B 67 8A C8 0D 3D 7A 94 B4 85 27 AC EB 71 99
 9E 87 69 A5 96 8F 2F 09 AD 7E 9E CF 26 86 26 33
 68 21 1B 36 D2 A0 49 A8 74 2E AA 94 B7 AD C9 36
 0B 0B 33 76 AC 06 93 AA 63 08 F0 66 47 ED 00 C6
 FA EE 69 A5 01 86 88 AE 51 22 C4 C1 25 F2 9D BB
 14 D0 79 F6 E0 CD 2E 16 02 70 F5 AA F9 09 52 68
 89 2A D2 D1 2F 5D 90 AE B8 58 57 90 2E B9 B7 D8
 53 38 FB A3 96 CE F2 06 EB 07 06 AA BA 5F 29 42
 39 20 E0 E4 DC 53 47 63 27 99 1F 6F D0 65 7A D2
 43 CF D9 63 72 CE A9 E6 88 49 9A 82 50 58 36 7F
 02 5A 67 61 FD B1 CF AA 83 28 FE 3A 83 2E 5A 57
 2D 04 0C FA 17 83 C3 03 D1 15 56 EB 43 A3 3D 9A
 8E 30 24 92 56 94 0E 94 3D FD 57 6F 86 B4 9E CC
 BC FA 5F 7D 0A 8E 9D B7 88 25 5B E7 C8 AC 07 9E
 56 14 D7 F5 28 73 BE 1A AC BD 61 7E 86 BF EF 67
 C9 09 52 20 35 3A 02 D7 3D BA C3 BB 48 E9 96 A3
 57 39 11 10 2C A3 9F B0 7A FE 6A 36 AC 36 84 BF
 BA 86 BC 5D 02 AC EE 50 D8 CF 28 ED ED 3E F4 05
 57 09 60 3A DC BE 8E 80 97 47 67 25 8A F9 99 FC
 DF 39 6F 76 8E 23 FE 35 6E 62 17 AF 96 AD CA 30
 4E 9C DB 5C FC 97 60 B7 31 50 B8 C6 54 B9 D7 59
 83 8E 88 E3 FE 45 BF 99 A0 45 6C C9 EF D1 55 05
 83 7B EC 18 FD 18 38 CE 40 E1 83 51 12 49 16 F0
 EE 36 8D DC 21 F4 7D 1B 2E 05 E2 FF 57 70 3F 15
 25 B9 60 96 E9 D8 97 73 A3 6B 26 A9 5F D2 FB 3B
 0C B5 F8 E1 DB 6C 4D 61 4E 3E 9B D5 95 97 B4 4D
 2B F3 A4 BB DB A4 77 25 87 D9 78 FA 78 3E 87 D6
 4D 1D 7F 6F C0 18 F2 56 50 5C 94 25 F8 C7 7A D0
 51 BF DD DB 3C 09 28 13 88 E8 49 EA 05 EA 60 A2
 41 EF 52 CE 75 D9 3F 56 01 51 DD 29 C6 9A 53 8C
 58 6E 76 24 5D C2 7C EB 1B A7 30 95 8C E8 83 78
 AA CE BF 5F 2D BF 9F 57 E7 E4 7F BE 59 28 4B 8A
 F0 77 12 6D 24 CB 4A C1 21 80 F0 25 82 9A BF 45
 A7 86 6B AE 9A C9 AC B2 AA 53 7A 50 58 01 DC 96
 C3 72 FB BA D9 77 75 E6 6D 00 22 C6 5D 5C 57 73
 2B 16 47 64 CF 1B 95 A7 2F D5 00 C6 2F 65 EA A1
 0E 0A 85 EE EB 46 66 D7 0C AD 84 17 8B FE 06 2A
 1C FC C1 C6 AB 91 24 79 B8 A8 A1 4D AF A2 F5 E6
 BF 9F F7 83 BB 28 27 91 69 5B 7D D1 67 E8 79 61
 4F 06 D2 0D CB 0E 0E 43 DB 97 6E C6 8A 6A C7 B3
 94 1F 1B A7 54 EC 13 4C E5 59 40 5E 96 B9 37 9B
 D5 FC 0D FE 87 4F FA 92 36 AB 11 5F F0 B6 87 E2
 5F 1B 5A FB 71 7C 3B 00 5C 10 8D 27 D6 FF F8 CD
 FA 04 7A F2 FD C4 DA FA 27 FD 83 1A 05 FA A2 99
 75 1A 3E E1 39 43 31 B9 7C A6 55 58 28 65 1C 8A
 20 CF 5A 60 C6 92 85 12 36 14 A2 65 B6 09 82 53
 DE F7 C5 E3 5E 9A 4C 9B 3F A7 8C 9F F9 0E BF E2
 33 A3 E9 32 DC ED F2 88 4E 83 0A BB DE 1B 25 72
 9E EF 0E AE 74 E9 BB BC 24 53 6A F3 CF FC E2 90
 17 84 3A 60 E5 BF BA CE C1 C2 33 E4 56 A3 01 B8
 87 33 02 B9 E9 26 75 70 E6 9C 1A 95 7F 4D 94 F6
 38 84 07 DD BA C8 11 AF BD 3C 73 D0 9C 10 BB 95
 62 0E 58 B0 B8 1E C0 EA B4 57 4C 91 4F BE B4 DE
 13 7A B3 4D 28 72 C1 D2 BA 6D CF 3E EB 99 70 30
 1F 9B 6E 7C 42 AB 1F 0F 77 60 C6 0F E8 32 E9 10
 E6 2A 5B DA 83 CB C9 DB FF 03 95 A9 10 36 8B 08
 11 64 FB DC A5 AE A9 1C E9 CC CE BB F1 19 A5 DC
 6A 55 82 F5 EF 2F 87 6C 8C F8 43 41 C2 7A 8A D5
 F6 88 99 17 B2 A8 4D 6E 09 2D A4 CD C2 CC B5 95
 BC F5 54 5A BE 1B 1F C6 D7 0A 9D F8 D5 D4 BB 0C
 1C 2C 4F 30 B7 54 BA 20 0B F6 AE 5C 67 7D DF FF
 04 E4 68 65 60 71 AD 07 AD 0C 49 67 51 45 D7 B5
 79 74 8A 64 78 AE 85 4E 60 BF 3F 03 EA A1 77 2F
 DA 7A D3 6E AE F3 88 1A F0 CE 98 3F 48 54 56 9A
 97 16 87 D6 47 64 14 DB C7 71 27 EA 6F 3A 3B B7
 F4 A1 F9 25 17 8F 83 8E C3 6C 3C 20 99 FE 00 16
 76 8B 83 EC 35 AB 21 CC 98 CC DB 02 72 E0 3B 25
 22 DF 85 AB EC 8F BC 88 0C AE 06 17 D9 65 67 45
 94 AA E6 6A 7D AA EC 90 33 A4 9D 93 A9 CA CE 6E
 06 2C 0D 01 4A 3E 17 49 C2 22 7C 28 AA 1F A1 F6
 5A 71 B9 54 17 C7 B3 AA 43 EB 9E F8 E0 7C 10 F8
 48 CB 35 A8 75 77 E7 DF 18 DD 2C 0D DF E5 CD EB
 F8 B5 5A F6 26 8E 5D CD 20 4E 20 E4 29 B2 65 21
 A9 6F 11 7B 59 1F 1D 87 BD E8 F3 C9 87 38 BF 16
 6C 14 62 E3 D2 4F ED B8 9B 53 C6 EB DE 0F FE FE
 85 00 A7 E1 31 64 27 14 54 7C 45 94 94 60 67 A5
 8D 2B 9E FB 65 E6 AF 0B 16 D8 5F D9 6D 63 BE A0
 CD 57 39 15 FD 59 32 C5 D0 FD E6 63 F5 64 83 D6
 2B 51 7F 20 0E 43 9C AC 9A 04 0F 0E 41 55 93 7D
 79 99 6F 18 DF A9 39 A7 59 B5 94 71 1E D1 FA 9E
 20 9F 47 B5 6F 92 30 32 79 6C BD 86 7D 8F 2C A1
 D5 BE 62 6A D5 E6 4C 09 60 78 52 BB FE 70 EF A4
 4E 87 EB 53 7C 8C 8B CC CC 04 6C 5A 89 9E 9F F6
 85 CD BF E3 B9 C8 0E BF 65 EE 6D 24 02 84 A4 BC
 98 B8 83 A5 AC F7 C0 F6 79 32 AA B6 1B 0C 33 DD
 C4 85 5B D0 F9 17 9A A0 F2 DA 2D A3 C2 32 49 98
 67 26 D5 DE AB D7 82 49 82 5F 4B 54 7A CC 66 03
 9D 88 09 83 AF 98 CF 77 1B 1B 5E 43 FB 3F 6D B0
 8E 59 C7 B6 5F 19 4B 57 D8 C7 E7 E7 CE B5 5B 91
 5D E4 50 79 EC 86 8D 0C 61 63 C1 94 AB F3 E7 BE
 78 2A 7D B6 D3 83 CB 9B 6D 1D 55 9A 01 01 5F 7F
 AB 41 69 59 1B 53 DF 6E 81 AD 79 36 91 D5 09 B0
 92 30 E1 AF E4 75 8C 18 0A 6D 50 A7 3F 91 7E 6D
 AB 84 E8 AE 70 85 BE 0B 92 63 CC AF 8D 10 37 74
 BD 68 C9 96 41 0D 1D 4D 56 36 0B 4F 50 18 0B 95
 71 B2 C9 DC 91 82 B7 59 4E 97 60 B5 C5 09 7A 59
 F7 A4 2C FC 96 72 0C 69 46 F6 F8 9C 47 B4 35 92
 35 CE 7D 30 B3 56 53 BE 82 80 2E A0 FC 27 06 CE
 E3 76 BC 89 63 3B 4E 13 59 D1 57 CC F4 D0 60 40
 30 C6 D9 E9 E9 5C A0 37 CE 71 6B E6 FA D7 46 E1
 58 3D F4 8D 83 D6 E6 8A 35 96 A3 43 B5 83 AD 4D
 06 11 5D 64 EA 18 FE 58 89 D4 3D FB 44 F8 CA 85
 25 F7 62 B0 AF 03 78 2D D2 9D A8 FD CC 45 65 9D
 C3 75 15 93 EA 70 75 83 C8 14 A4 40 95 C7 D0 85
 D9 82 C8 5B EB 49 E9 F4 C0 AA CB CF 8F 0C BB 3A
 6A 44 04 F2 F0 50 E3 99 6E F7 3E 18 32 C1 5C 24
 44 27 F6 66 C9 C8 63 BB 1D 26 31 BB C0 50 C8 4A
 57 A8 11 D3 BC A0 FD 65 BD 72 F6 97 03 65 E2 EC
 4C 70 91 99 83 D4 3F 18 C9 B9 14 DE AB 64 EF 7D
 01 66 AF 97 23 EE 76 27 A2 9F 1B EB 7E 08 44 30
 60 46 EC 93 14 48 C1 82 D5 3E EA 5F E7 29 E5 E8
 39 FE 7A 36 E9 0F 0A 31 9C 1C EC 82 85 4C B2 15
 8F 25 57 10 44 74 CB 01 83 79 D4 FF 17 19 57 C3
 EA 9D C7 5E 98 52 87 83 B4 24 C5 D9 BC C7 07 16
 9A B2 14 A3 CB B6 C1 33 C1 9C EB BE B1 CA 74 24
 56 D7 D1 86 8F 72 88 05 1D F7 FE E0 76 19 19 38
 D4 B0 9E 3E D6 CF 79 90 02 41 FF 44 06 70 1F 0C
 EE 11 96 F6 E9 53 3F 1A 13 F3 7D CC FA 7D 6B 9B
 C6 9F C9 01 59 FA 28 E1 D1 4A 6D 1C 50 CA B8 02
 2B 84 AD 26 05 84 D0 63 0A DB 1D FC F2 46 67 8E
 F2 6D AB FB B6 22 30 D1 93 C4 97 9F BE 4D 8D B7
 2E 46 FA 6F F9 B2 9F 61 0E EF 7C 31 A1 3E 46 1D
 60 A9 FE 64 F1 18 56 C6 5F 27 56 53 F8 DF B2 28
 20 0E 6B B8 02 36 AD 33 77 6D 2B A6 15 B6 D4 04
 C0 06 CA 30 E5 B2 D1 C4 9B B4 11 17 03 30 94 63
 0A EE 42 5B 9C 4C 4E 27 C5 63 01 84 A3 42 54 DB
 B0 79 1F 17 D8 74 79 50 6A DE E7 14 0C EE 4E FC
 25 5D CC BE 7F 99 76 E2 EB 44 B8 4E BB EE 17 D4
 5C AA E4 4D 76 F0 D7 86 50 9F 2B 31 6C 83 6A 8F
 EE E5 CB 44 F0 AB B0 B7 C8 F7 E3 43 B7 81 CF 98
 5B AA A4 F2 18 B3 48 CC C2 B7 84 8E 4C 28 E6 39
 95 EC 39 BB 63 43 E9 23 7E AC 16 20 57 D7 8B 13
 92 84 C1 F1 54 78 03 28 DD 7D 5A 31 C1 89 09 1C
 56 19 6C AF 90 9B D8 28 55 9A 81 6E F3 01 9F B2
 26 EF 9F 40 BE 5C 7A 80 68 6A BE D6 34 B8 0E 6B
 E6 46 AB 4A D2 6F 41 4F 97 96 CA 95 45 1D B0 DC
 83 B4 A2 D6 AB F1 75 03 1C EA 30 33 E1 51 A2 7C
 B7 61 4F 8A 19 49 47 D8 5A 41 E0 2B 27 F5 CA 94
 97 44 B2 BD 37 7D D5 10 45 84 B5 1A A6 B1 C9 60
 66 01 3A AE C4 B0 E6 E0 C9 F1 20 99 8F E0 EC 0C
 B1 F5 1E 7E 38 CF 3F B2 63 8F 86 E4 37 D5 14 CA
 BA 5D 88 43 EB F9 8B 95 75 D6 1C A5 60 7F 80 AC
 B6 21 AE 27 EF E0 C5 6A F6 86 35 A6 D6 D7 DB 53
 EC 84 D5 00 E4 48 9D 6E D9 C5 B9 B6 37 D7 A5 E9
 7D 8C CC FC 0C 04 FF 83 21 77 E6 3F D7 55 F1 D9
 FC D8 87 0E 3E DF 99 50 DA EA 77 AC CF AC 9F A1
 4D 14 3E B3 98 EF 19 10 8C BB 57 E5 B7 70 17 2B
 A4 74 4D 2F 60 F1 DD 0E FA 78 E3 E0 3C 0F EA 2E
 4E 35 D0 16 36 B2 84 51 0F 91 62 86 44 73 35 31
 D4 1B BB 0C 8E 8F 93 68 53 1E 02 2B C8 A1 B4 F0
 23 61 C1 9B 76 66 2E CE D0 81 C5 68 AD F1 5D 8D
 80 5B C0 D0 23 5E B3 99 98 FF 55 4A 7C 5F B1 10
 F2 4B 92 BD 6A 37 9D 88 1E 3A 57 63 42 92 93 D6
 A2 B2 DE 19 6B 52 CB F8 BA 90 4B 77 3B 54 B2 E4
 36 02 58 C0 C5 F8 90 3D 8C C2 7E 0C 1A 11 FD 99
 1E 93 0B 9A 53 C4 5C 3F 02 98 C0 4B 34 1B 6B 46
 41 F2 BC 9F 7B E9 23 56 A5 6E B7 6C 8C A9 0F 73
 B2 0F 94 9C 85 A5 F0 D0 F6 82 9F 01 D2 29 97 E0
 18 12 00 0E E0 80 23 E9 34 E0 24 2A 66 54 6E B6
 63 9C 89 4B 3A 7C 42 8B C8 E8 A6 58 EE 70 02 B4
 01 CF 6F ED 0E 65 AD 31 CD 9F 19 B2 95 A6 EF 94
 67 A7 4F 0E C7 F1 F8 6D 19 1D EE 16 BC 60 BA 77
 F7 2A FB 03 C6 A1 EC 21 A2 89 3E FC 27 1B 9B 7D
 6E 89 81 69 FF 7E DF F7 E5 2A 07 2F 6B FD 58 2D
 69 C6 B0 F0 80 CA F3 E9 EA C8 34 86 7F 21 2E 31
 41 29 88 E5 24 DE CA 2A 98 54 7D 58 E2 99 E3 AC
 A9 48 82 68 F7 93 5F 41 FB 0C E8 2F 84 27 AF E3
 77 B3 97 7F 1A 75 DD C8 B9 AB 9A A1 EA 8E 9D 0C
 4E 60 94 47 9A AF 46 B1 E8 5E CC 3D 33 CC 20 F6
 E8 B0 23 D1 1B 8C 9B 0C 9B DD A5 22 5E E2 AC 2E
 4B CE 84 A6 DD FA 4F 2A E2 54 C7 48 2E 7B B8 63
 0D C0 BF 88 B2 6C 64 A1 66 FF C1 F9 B3 E1 CE 21
 3A 03 43 A2 9D 5F 3F 1B A8 FA 6A 6F 9C 12 9F 84
 DB 70 D0 A2 92 5D 89 04 49 0F F8 F4 F3 07 D6 32
 22 48 E0 9B 9D 34 DD 68 D9 A3 FB 22 46 B0 D0 2A
 8F D5 DB 8F B5 A2 EC 6C 3C 74 81 E3 B1 FB 9E 64
 F8 C4 0B 2F 28 A4 04 6C 42 C9 AA 3B 19 F5 52 CA
 EF 8B ED 62 CB B9 B5 93 A7 58 2E 14 60 FE 71 CD
 2A F6 E6 D8 1A F3 B5 5F 98 61 68 65 6C 4B F7 85
 8E 8F FE B7 84 69 55 5D DA A0 79 F4 32 E9 89 0A
 CE 61 C6 D6 3C F4 81 B2 9B 4B 0C 2A 7D BB EE D3
 A3 80 5B DC 6A 67 67 EF 32 40 C1 CF 6A D6 DF 2C
 34 27 87 CE 66 7C 55 B4 3E 27 AE A8 5A 6F 71 9A
 4D AC 52 79 8B 1F DA 4C 0F 41 D2 FD E9 99 21 1F
 05 49 84 69 DD 55 AF E6 D5 53 F0 81 F6 1B 11 90
 B3 D6 DB 68 E5 1F 09 83 01 71 6A 07 5E FE 2A 30
 83 04 46 BC 6E 80 6C EF 6E 38 6C 20 A4 E6 C1 F8
 09 F2 7D 0F 73 25 9F A6 2F E6 D3 C9 A8 74 5F 36
 70 1F D7 04 6B 63 6E 76 18 2A 8A AD A3 57 76 82
 7E 13 E4 1E 7E 6C 03 0C 85 AE 8C D7 7F 95 1B B7
 0A 50 87 F9 91 9B E2 6B 16 1B B5 69 D2 78 1F DC
 FA 5A 05 4C DB EB 0F 2E B9 50 D2 0C D0 89 3E 6A
 D9 0D 8A D7 95 4F 78 1D E4 8F F9 44 3D CF 61 D2
 F5 74 A1 96 5B E2 6C 04 36 99 18 37 4C 3B 18 8F
 72 2C 96 74 98 2C D7 71 E1 6A A3 9B 2D 11 CE 15
 8B 32 60 4D AA B2 B8 CD 9C 90 A8 85 73 FE A8 98
 54 9E 93 DB 74 72 FB CD 0B 68 3E 93 AD 0E 5B 1B
 8E 8E 75 EA 71 CE 28 7C 21 C3 0F 07 84 0E C8 DB
 BD C0 DE 1F C3 C2 E8 C7 6E D7 19 C8 8D D7 DD C8
 71 A6 3C 47 B5 D4 49 6B 8C A2 90 77 DF 91 D5 46
 25 87 96 DF EB C5 49 A9 F5 4B 2F C8 04 BD 42 4C
 37 DE 39 92 C5 F1 35 F4 D3 4E AF 93 24 E0 11 73
 AD 46 01 14 C3 29 78 AE AA 28 BF EA 57 D5 76 0D
 3F 76 F7 6E 46 7B 7C FE AF DB 64 82 58 9A 3D 69
 1E 2E F6 12 B1 5D ED 1A 9C AA 0B 66 A0 CE CE 15
 63 18 BF 73 DB 91 35 F7 38 27 23 CE 35 37 6B C8
 39 8C 44 30 53 84 CC 4B C1 59 9D 5F EA 55 5C DC
 ED 5E 4A B2 50 14 9A 88 99 05 D5 23 51 26 13 FC
 B0 B9 B5 88 21 25 91 64 97 96 C8 64 52 10 28 77
 4C D2 C3 EE 53 4F 67 14 B3 C4 7F FF 82 8E A2 6B
 4F C6 6A 37 42 6F 02 08 E8 6F CB 36 17 E1 0D E3
 16 B7 56 B2 BE 25 50 1E 73 DE 96 C8 86 39 BF B0
 85 E6 55 AC 67 76 1D 49 14 32 ED FB 6B 9D 12 4A
 9F EE 3C 18 17 1D 1B 46 7D 18 BC 72 AF E6 1E D4
 DE AA 36 E9 4D C4 79 A0 67 A7 E1 B6 FD 75 F2 4B
 BD A4 1C DC 1A 7E 51 F6 84 37 8B EB 87 4F 7D D2
 63 A4 5B 0C 72 36 1D 97 35 31 6C 43 40 91 28 19
 E5 24 00 66 44 4A 5C FA F3 1A E3 F6 E6 CA 6A 3C
 DE 1D 66 BE 0A 93 F0 89 5C 15 07 F2 78 1B C5 C5
 C7 8C 4D BE C8 59 B3 EE 88 6D 71 63 1A 83 39 33
 5B 75 9A 36 AB D0 7C 59 4B 79 B5 BA FE 12 2A A3
 4A 08 69 E0 98 32 3E 1A C6 A6 1A 94 7B 4F A6 D6
 3B 5B E6 AC DE 76 AC 62 4F 10 09 A9 36 E3 58 3A
 6E BC 37 F9 69 DE 15 19 E4 C0 E6 46 C5 42 1A 5E
 CA 26 73 01 40 D2 C5 86 71 CB E3 AA 8A 44 AC 1C
 D6 FF 31 3C 96 91 2D 8F F3 A4 92 C5 1C FB 3F D4
 9F A0 8C C2 21 65 DE E4 AC 1E E3 AD 5F 34 02 41
 98 82 50 D1 40 64 79 41 85 C7 01 9E ED DA 36 26
 C7 B5 DE 73 30 DB 75 30 D6 1F D4 82 15 78 A7 D8
 9B 6C 45 DA 29 F3 B9 1F 29 DD A9 61 E8 B8 FD EC
 C6 38 9B 70 EE 3A 3C 74 B3 F2 A9 AE 56 8D 7B 4A
 E3 FD 8A 66 30 0E A6 33 E6 FF 92 8A C0 75 CF 45
 BE 53 79 74 93 EE 0B 8E 5B 67 18 ED F0 2F 46 D7
 E5 D4 2E 9D 02 2E B1 7E 27 67 AA EA 6B FC 97 64
 65 18 78 2D 96 83 B3 F8 E0 AA AA 04 12 62 80 B3
 94 31 00 7A 4F 48 BA E2 60 41 09 3A 9F 68 F0 D6
 03 8D 39 DF FF EE C6 54 6B F2 17 2B 3F D6 80 0E
 F4 A5 94 C2 7F 69 D9 33 AB 16 C8 10 CE BE EB 21
 E9 F3 6E 34 9D D0 9E 04 B5 A0 D9 D5 35 94 DB F9
 52 15 A3 D0 FC CD E9 DE F3 31 21 B7 5A A4 BB A3
 40 20 38 C1 10 2E 24 E7 70 17 44 15 16 E6 BE 65
 51 37 57 F4 AF 58 A9 2F BF 0F ED 24 E4 42 68 8D
 74 AE 16 58 B8 8D 83 B1 98 37 8F E6 82 13 5D 83
 55 1D 5F 03 8E BC 09 1C A0 F5 26 DF D7 33 14 6C
 14 23 B3 92 2B 52 9F F4 C6 B5 85 7F 43 8D 47 2F
 CD 06 C0 A8 C0 90 EC 0A 62 30 98 EA E2 80 3E DC
 63 D8 F0 A3 A3 DC 91 04 93 01 3E 0D 52 A5 F7 92
 71 15 B1 DF D3 8D 0D 9F 8B 4F 90 E3 90 61 1A 69
 8C F9 FB 4F A0 00 62 0A EF 2F C2 AA 92 75 47 73
 C1 99 93 C7 11 5D 4A A8 37 15 C1 CE E8 D2 6A 41
 FC 07 AC 27 8D 4C B5 AE F4 4A 2F B3 C3 10 7B 14
 7A 2C 2B BA C8 77 95 EA 2F 68 D2 BA C4 80 32 55
 A7 40 49 EF F4 D3 5E 91 6C 19 F0 82 CC D6 94 43
 1C C3 0F DC 55 B8 47 47 3A FE 7B 81 A9 1C C2 67
 A0 E1 E4 08 3E E3 A4 D1 DF 7E BF CB 92 C3 88 03
 03 3A 4F 44 93 F1 DB CB AC 00 27 06 3A 55 FE AD
 8E A3 95 34 F8 21 6C 30 5B 38 C8 F3 42 69 75 C2
 C2 64 1F 0A D2 5A 47 EB 48 EA F6 56 A4 5D B5 60
 74 94 5F 05 A7 CD 51 A3 B0 9B EA 7C 35 79 A4 9B
 6D 4B 13 7B 3D 39 5B A8 A7 18 36 34 00 D0 14 8D
 E0 6B E4 F5 02 5D BF C4 EC 70 28 40 CD DD 2A 04
 12 BE 00 83 54 14 44 DC B2 1C 05 15 1C E1 A6 23
 B4 24 23 FF B7 ED 0E FE A5 B1 83 0B A9 7E 73 E0
 12 70 17 C3 7E AA 6E 31 45 09 74 3C 42 00 47 29
 0E 79 18 05 07 42 10 FB D7 A7 60 BA 16 1A 40 53
 EB 5B DE D2 D8 80 3E 8B BE 27 9E 24 E5 E8 46 BB
 33 A9 C5 66 C8 7A E2 48 EE C3 24 56 69 69 C8 3C
 F3 F1 55 65 5C E2 F8 5B AB CA 7E CB 02 28 EF 0F
 43 12 81 32 AA 33 18 92 2C E1 81 0A 39 0C A5 45
 86 12 6E B1 35 71 2A C8 68 D2 6D D4 0D 97 0E CF
 B3 FA F2 18 92 BF AF DF 2C 6C 30 BD 19 61 A8 A2
 92 7A 2D 64 3B 81 13 A8 EE 87 91 7C 68 BF F1 D5
 CE 62 0C F9 F2 30 F9 2A 13 10 9E B2 FE FE A4 E7
 54 48 82 0B 30 EE 37 67 20 A2 32 01 2A A5 73 3B
 50 02 FF 86 73 69 D0 4B 38 93 FD A9 15 EE 1E 2C
 DA 5B AF A8 D4 6B FE 5D 0E 8D E4 35 88 34 69 E0
 D7 40 8B F4 EC 31 8F CB AB 27 57 47 E4 6B EC B0
 09 CF EB 92 B9 F3 66 E5 79 1D 9F DC 35 6F BF 17
 AC E1 27 C3 58 68 BB DA 61 14 E1 57 62 FC 99 80
 58 F6 26 79 95 D7 27 92 41 2D C9 CB D6 04 61 3E
 89 7C 29 B5 30 70 E1 42 94 30 B6 CB E9 2F E2 7B
 99 F5 A4 26 55 DC BD F8 1B A6 DE 68 3D FE F2 36
 0F 94 A9 18 56 42 6B 50 91 21 02 35 7C 8F CF 11
 B4 BD C8 85 54 35 2F 68 DF AD B5 D5 FF 8D 50 7A
 96 C1 C6 82 CC 1B 42 9C 99 64 BC 8C DE 1B 70 E0
 04 8D 93 8C E6 F8 86 F6 A1 4D 97 B2 43 76 22 9F
 7D 8C 85 E5 BA C9 EF 09 E8 4C 23 0C 46 F2 5A 0D
 70 47 A2 E0 18 69 10 E4 56 FC 57 81 46 96 5F F1
 C6 20 DA 32 B3 62 AF A9 10 2F E5 3D 93 5D F4 01
 34 A0 C0 E5 C2 C3 9F 20 EB 37 DA 62 CA A4 46 AE
 7B 7E 21 56 9F C6 38 F5 95 2F 12 7D 37 1E D8 EC
 42 92 E4 6D 46 B3 E3 65 C9 2E 82 3B 52 92 5F 2D
 57 2A 8B 27 8B B2 D4 32 CF 3F A0 B4 16 9A 90 54
 E2 4A 24 26 9C B7 20 CE 6E 9D 28 7C B0 6C 0B D5
 EF 2C 93 D2 FB D7 67 99 36 72 4E 20 92 E3 E7 96
 DE F9 3B 91 42 19 03 E4 42 FB 34 27 AB FC CB 3A
 B4 74 15 7E CA AA 1F CB DA D1 59 41 D8 DE CF F6
 07 20 0A 81 F6 8B ED E5 EE 1F 2B 8E 99 47 B6 0A
 1A 01 F5 45 59 35 92 9F E7 77 79 22 00 70 B5 D2
 CD DA 3D D5 2C 7F 56 DA 18 D4 48 76 AA A8 2A 2C
 4E D8 5E F5 42 36 29 E1 B1 6E F7 8E 3D 4F 3E D2
 7B 84 D5 8A DB 09 E9 19 9B 76 06 E9 CA B5 7D 9F
 4B F3 50 89 F3 37 1B D6 87 18 72 C6 92 96 30 E4
 E1 45 13 A7 E0 11 ED 84 78 C8 FE 02 8F D8 C4 15
 A4 17 F7 78 E4 58 97 A0 5B CD 65 64 D3 DE E7 63
 52 C7 83 1F F1 FC 1E E8 97 35 CC FB 37 E1 7E 9B
 27 D7 E0 74 F2 EC FC DD 1C 7B 7A 32 76 41 1B 07
 1E 0D 18 E5 75 80 D5 8D D8 34 A4 CA 65 74 B1 14
 D3 82 83 E0 F7 6C 6A 14 E3 DA 81 4B D7 00 63 21
 75 E9 10 CF BD FE 01 3C 23 90 0F 4B 9C 17 90 AC
 3E A1 A8 29 BD 09 DF AE A5 76 79 51 B9 04 AB 5B
 55 77 E5 35 42 E7 38 17 8F 0E 37 5D 6B 44 FA 41
 15 A6 0B 4F B8 BF 5A F0 53 6F D1 00 A0 63 C7 EB
 1A A3 5E EC 75 18 41 9B CB C5 41 8E C2 5E E4 7C
 3B AD 56 60 84 06 A2 28 B2 A6 DC 19 70 79 A1 B1
 D8 E0 47 3D 86 C7 BB 66 92 C4 DD B7 1D 03 83 03
 B2 04 ED 1C CA CD 79 6D EB 61 F0 94 02 5C FF D9
 43 CE 9A FC 7C 0E A7 72 76 C5 FC 54 B0 C9 E8 E9
 75 FD 12 14 C9 F5 A8 1A 6D 82 D4 EC D1 7E 5C CD
 19 B5 7B 16 5D 39 3E 40 44 36 86 39 CB 82 39 0D
 7C D1 36 DC 9E FC AC DD 65 D3 CB B6 44 87 74 DA
 9E 3C 78 60 38 19 45 8B F9 F6 DA 05 57 29 3A 95
 B9 1B 02 5A 3D 10 1F 6F 68 7A 46 8E 3C 20 40 AE
 8E 0F 3A 00 83 C8 6F 31 B0 D2 20 4E 4B BB 2F E8
 EF 97 19 A0 15 D4 A9 03 10 04 9D A6 B2 90 84 D5
 97 AC 20 E7 F6 83 16 4D 02 5A 49 D9 71 86 25 19
 A0 4D D3 5B 43 C8 93 FE BF 94 B9 73 C0 24 70 92
 24 DD 62 DA A1 A9 FF 07 47 94 89 2E 98 7D 8F B3
 2D 86 87 D0 F0 9D E9 57 69 92 4D A5 35 5E AE 30
 89 F6 88 6A 4E 77 B3 61 E9 A2 BD BA 9E AF 0C 74
 77 E0 56 B2 1C 26 53 1A 25 EC 85 65 3B FE EE 65
 A9 1A F3 8C 18 BD C4 F5 90 4F EE 75 04 F9 05 07
 3B C3 7A 9B BE B4 C9 15 7D 03 5B E4 75 74 B0 F9
 B4 04 79 28 49 38 7C AA 32 C6 34 07 CE 20 E7 F8
 6B 3C E3 C5 B1 FC CA B7 CC 73 80 71 18 F1 C7 12
 97 86 5E FE 23 62 A3 32 11 0B 74 85 19 13 15 0A
 D1 44 82 7D C2 FB B7 51 39 F7 13 93 AD BD 79 E8
 A8 BF 91 C2 29 9D F3 73 48 03 7C 59 7D 74 F0 6D
 DC A2 47 BA D6 65 E0 D5 50 05 C9 6F 5A 45 53 9F
 F1 90 40 0D CE A2 14 6A 27 C2 75 35 88 98 35 D8
 8E 0F 80 5E 6A E1 1C F4 69 82 D6 68 9C 5B 43 DB
 3C 28 EA D1 B9 C7 12 6B 54 41 CE 65 B7 56 1D 26
 51 D9 3C 99 3C BE B7 6B 2E 5D 5C FA 4D 2A 81 7F
 D5 F4 51 64 94 62 DD A4 EA 0B D4 48 77 0F 21 23
 8B 44 A1 E5 A9 FF 45 C7 47 65 4F 64 85 35 AB 67
 DA DF 7E 61 9E 2F 2D D7 A2 D9 73 B6 DB A1 84 D7
 D6 15 C5 0D D6 C3 A5 CA 2E 1C E5 26 C6 C8 7F AD
 E9 BB EF 7D 6C 0A 33 DC 5E EF 05 45 34 90 86 D6
 1F 2D 68 9C 9D E5 D8 F2 91 A0 9D 20 D1 41 A1 30
 D2 62 C8 BC D4 07 BE 14 52 5D 81 B4 07 A7 C7 91
 13 53 55 BF 11 B6 A6 DE 74 20 2E D1 A8 D7 66 D8
 7A D2 62 16 DB 41 9D 7C B9 D8 F6 8D E9 00 1A 1C
 FB 69 9B 99 3E 4A 04 B4 4F 62 7F 8A 32 12 06 DF
 4B 66 DE 5F 8F DE D9 24 5A 22 90 EF 43 88 11 03
 8A 63 CC BF 9B 30 C0 13 99 D5 B8 14 82 19 8B A6
 0A BC 60 70 A8 91 83 9F D1 F8 32 84 62 49 32 6E
 87 74 DA 2E 8F 94 14 0E 60 82 FC 63 2C 29 11 E5
 E4 67 60 44 CA F5 3D C2 E8 85 1A BF E2 73 6E 55
 60 66 AB 99 D2 07 C3 CB 3D 35 85 F2 75 59 A7 28
 EF 60 A9 4F 71 8D 7C 63 65 82 AF EC BB 2D 47 65
 BF 6B 40 E0 93 0D 99 E2 72 EC 0F CD 04 83 9A 61
 6A 48 6B 87 0D 91 C9 C5 A2 C6 5F 75 BA 97 8B 5C
 A0 D5 4B 46 E2 96 5E D3 F3 D1 9D B5 07 B6 BA A5
 0F C2 75 85 AB 96 83 09 51 11 90 46 B2 34 00 C0
 74 33 62 21 F7 6B 73 DE 8D 6B 68 D7 8C D7 AB 24
 6E 93 0E A4 E4 3D F6 83 24 BE 3F F5 9E D5 61 E8
 1C 33 85 B0 9C 3B 64 FC 58 B5 E5 0B A4 B4 28 B2
 C7 C3 C9 26 6B 5F 12 7D BB F7 77 8B 97 FB 1B 20
 18 2B 56 26 9A 55 3F 1C 91 7D C0 5B AB 59 E3 C4
 B7 50 F8 0E 2F 48 6D 1E FF 4C 9B 5D CD 27 43 82
 2E 02 8B C7 E7 35 82 3A EB A4 01 B4 2F 24 77 B5
 3E A2 EA FF E0 09 E1 C0 8C 1D E5 79 9F AC 6C 73
 8E 33 13 13 BA AF F4 35 E9 21 07 D2 58 E3 E5 11
 63 34 7E 4A 71 A0 57 F6 25 26 8D 4F 4A 99 24 E0
 A1 07 6B 9F 11 10 AE 41 2F A7 09 56 F4 07 8B D7
 F3 A3 0A 56 05 FB 66 5C BF 92 46 41 69 37 D7 E6
 9B E1 D9 50 AF BC 79 D5 E0 AE 5B 61 7A F9 78 7D
 0A D7 70 BB 16 9E 06 53 F6 56 EB 8C 7F 85 7E E4
 91 63 1C 64 E6 7D 2F 27 07 1C 92 F1 0E E6 9E AB
 C6 D4 58 85 E5 51 D5 3B AE C5 BC 5C 0B 00 78 B7
 D6 24 27 AE DC 56 85 05 9A F5 A3 AD FF A3 80 8B
 CE F9 CF 29 7F B9 BA 06 DB 55 AE 83 DC D7 8E 29
 D4 A5 54 D7 72 82 CE 2A ED DD F3 24 10 11 9C 9D
 D9 3D 5E BB C7 31 D9 9B 34 F1 BB 24 D4 20 C9 B4
 03 B7 8F 61 8B 1D 60 F9 F9 71 01 4C E1 0A 49 AB
 4B 89 05 D1 92 39 44 CB 29 38 1C B4 DE BF C6 B8
 63 05 28 9C 28 55 6A 39 B8 73 D5 12 9F 1A CB 81
 D7 8D 19 76 7F 7B E7 4C 63 5A 59 83 7E FE CB ED
 56 0E 88 E2 49 F2 0E FC D4 73 EF E9 8F F7 C4 0F
 CA D9 81 CA FA 6C 02 87 C2 5E 38 9B 88 CC CF DB
 17 B8 FC 6E EF AA E3 61 6D E2 42 7E 69 A3 70 0D
 F6 72 FC 72 46 08 F2 0B 09 81 95 DD 7E 23 47 D1
 1B 03 DD 43 51 77 15 CC 1D D0 0B BE 95 1D DA DE
 83 74 D1 0B D5 E6 F9 DC BC C3 7C 98 95 0B 3A 94
 CB 07 11 DA 30 C9 95 F5 25 FD 3E AF 47 43 2F 1E
 ED A4 96 C0 42 6E EA 2D C7 49 A3 EB 39 67 32 C4
 30 B9 E9 EA B0 22 3D 43 91 2C 73 4C 83 AF B1 60
 6B 96 B4 82 BA 7F 70 6E B9 3D C5 2A 05 A6 C3 B3
 3C 1B D5 4A 41 C0 92 23 8F C8 9F A2 34 15 30 71
 00 1A ED 9D 51 1B 6D 76 B6 2C 9F D9 08 DD 2E DC
 19 C8 53 F0 23 7C A2 71 17 E2 BA 2E A9 64 07 6F
 33 06 4C FF E8 64 B4 22 1B A7 A9 41 5F D1 0F 59
 52 60 6A 43 3B FF 44 5C 97 32 FB 83 9D 00 48 F7
 7F 64 09 73 BF 4D BC 68 D9 B9 E8 75 82 8C 88 B7
 22 9B 67 87 1D 12 F6 AC 19 A7 0E E1 49 12 94 AC
 FD 44 FB 86 77 4C 3F 91 4D 31 23 BB AF 53 9C 8E
 D7 FF EC 30 92 A9 B9 94 C5 37 DE 99 14 E1 B4 D3
 48 75 26 4A 88 34 7E 49 75 2D DD A5 A3 B3 22 F4
 2A 55 F0 F6 2B 67 0F EF 0C 98 5E 95 4C FE 0A C5
 95 03 93 C7 9E 90 20 73 66 EB 4F F0 4C 66 88 73
 33 AC DA B3 D1 40 78 C7 6F EF D1 50 F7 D7 6C 4F
 53 60 3E 89 73 1F B5 D5 5F 3A E9 9A 17 21 D6 CF
 BD D9 66 B8 7D 4F 3C 55 89 FD E8 2F 77 15 6C E8
 13 17 55 E2 41 84 E3 75 C4 BF B5 AA A7 68 C6 C4
 D4 F7 3B 2E 97 22 15 13 E6 FE 8D E4 81 13 19 EE
 C0 2C B1 5F 48 F4 41 AC 4E B7 49 B4 D5 C5 3E 10
 E0 D9 7A 7C C3 2E 08 17 4B 52 ED 04 1E 96 3B 69
 7F A7 04 A4 48 C9 61 DA CA 3B B6 3F 71 C6 82 E6
 1F B7 5D 88 48 40 81 61 63 68 19 6C 9D 6E 01 D2
 AA 7A AE 6F 23 40 E3 9B 8A 23 EC 04 DE F0 B3 6E
 F7 09 D9 59 86 5D 62 6F 1D 42 3B 7E CC 15 86 1B
 F8 C7 3A 8A F7 A1 96 77 B9 75 31 9B D7 4A 4E BC
 74 9A 8E 32 35 7B 51 81 B6 4D 6F FE 16 63 49 48
 2D F7 AF 42 D2 98 7E 8C 1D 68 69 8C EC 53 DF 4D
 FA 4D C6 EB AB 42 C3 38 C7 89 CD 59 17 93 B5 41
 AF 29 23 D4 0A 34 00 60 C1 16 EE F4 4C 39 4B 3F
 30 00 B5 D9 54 B2 EB 69 7A 08 6A 7F 74 62 7F D1
 0B BD 81 87 B2 8B 38 89 34 47 81 59 BD 76 72 51
 01 1B 02 10 67 A7 5A 09 62 73 AB 2A E3 95 8F 58
 45 36 15 75 19 DB F7 A6 7A E1 07 B2 24 65 C8 C6
 CC 87 98 B5 21 F6 2D 30 10 6F 5D 56 D9 81 27 40
 B2 DE 54 6A C6 F5 A1 80 49 1F 11 12 D7 59 DA 4F
 AE B5 8E F8 9A E4 BF 00 BC A5 2C A0 BC 3C 0C 6F
 00 60 59 BA D2 0B 96 68 33 2C 49 E7 75 51 43 4A
 DB EA BD 94 2F ED 56 4D F7 53 3C B8 2E 64 19 EC
 FA 8D A9 81 78 78 0F FC 95 41 30 64 79 DD AF B6
 56 43 60 3F 2B 38 FE 0A 6F 23 8A 2E 36 91 71 90
 42 A6 63 55 07 8E DE A0 CF 40 81 FB 24 84 37 B0
 1F 8F F6 9C 95 1C 92 EB 80 2F D6 63 F2 33 0D FD
 BB D3 64 8E 2C 2E D2 B5 3A CE 15 5F 8E CF 33 5B
 50 7F 7A 20 00 66 20 80 F3 9F 4F 92 4F 14 78 01
 49 5F 47 3D 11 EE 30 EF 1D 3C C5 03 B6 78 5B 71
 6D 21 29 82 DF 02 3D 3A 0E 78 7A 1B 99 1B 56 30
 FA 4C 78 AD CC EE 3B 8B FF 28 64 E1 BA F8 31 75
 BF 2C F8 38 1B 05 71 D5 36 7F 87 10 60 5F 63 6A
 4D 51 DA 41 9A 50 D1 8D ED AA B4 B7 FD FD F4 BA
 48 44 CD 00 7C BE 36 B1 62 5F 24 EA 1C DE C5 78
 41 CB 2B 7B 7C E7 73 DB 15 75 03 EE 08 AA 1E A6
 1B 0B 5A 13 31 C4 DD 0A 13 39 63 15 C6 68 77 C4
 03 63 8E DC D5 4F 17 E4 C7 2D 41 0E 01 22 CE C8
 B6 38 1D BA 9A 83 A9 94 87 C4 4A 2A 9E 45 79 FF
 D4 18 19 28 40 7A B6 EA 25 7A 55 BF C1 43 57 9A
 DA AE B1 4F BC DB 49 4F 85 DD C7 78 57 BC FC F1
 D7 E8 D9 6D 61 EF 4B D6 60 E9 1E EE 43 27 65 42
 4B 2F E8 2D A2 BA EA 78 C8 D9 FE 5C FE 5C 06 77
 FE 1B B6 BC 47 8D 16 E7 5C F2 1C D3 B2 B7 29 4C
 49 23 36 DA 29 91 6C 29 74 7C 4E 43 2B DD 98 87
 B2 03 DA 31 CD CF 3C 66 70 82 71 9E 75 D5 82 28
 AC 63 B1 9D 62 A2 19 B8 D1 42 49 98 53 33 54 22
 02 7A 6A 2B 15 C4 29 2E 5D 72 05 EC D9 EB 55 3B
 DB EF 0A 7A 6B 88 08 E3 44 06 4A EC 03 37 EA 36
 61 5F D8 60 7C 55 FC 10 3F AA D9 C2 D7 44 7D B8
 48 F6 05 C8 68 CD 5C E8 49 D2 B4 22 23 FB 3C A6
 4F 87 F7 90 46 EE 10 A6 DF 5C B7 28 94 C6 75 1A
 5E 35 97 95 81 DF A8 A7 7A 1B 6C 26 2C 48 C8 E2
 7F 2B D1 31 59 ED 5A 07 5D EB DB 1F 34 87 B6 79
 2C 6F ED 5C 5D 4D E2 B5 49 9F 9E 75 1D BB 91 71
 28 33 78 48 FE 74 5B 59 2E E9 2A 70 46 53 3C 25
 BE 21 0D F8 DB CC B8 84 FA EF E1 D2 9A C8 B8 17
 72 27 54 0A EC EE E9 B0 DB 5B FD 58 B5 C5 58 9D
 C1 77 94 FC 2A F7 E9 DF 1B BC 9F 7D 3C 30 50 35
 8F 5A A2 AC 46 50 3D AE 43 34 20 74 83 86 44 17
 D9 04 22 49 86 7E 97 5F D6 AA 34 28 BA F1 B3 1F
 17 E1 EA DE 77 71 97 76 5A 5A 20 00 A7 99 FA 23
 14 F2 8E EB CB F9 88 F2 1F E6 1D 07 29 21 C5 72
 DE 1C 1E 0A 13 FD D0 89 69 C5 49 7F EA 54 DE FB
 ED 59 3B 6D 5F 20 25 DA 95 E6 78 9A 52 9E B8 FB
 18 57 50 78 31 97 6D E3 80 43 1B 42 5D D1 3B 5C
 AE DA 47 AC 05 35 8C 0E 35 AA 6F BD F3 7E F3 2D
 9B C3 D9 39 0F 5A 54 BE 46 60 95 C4 0A FC BE 97
 2A BF 78 91 80 A4 3D 30 E1 CA FC 28 13 61 D8 A2
 10 19 12 F2 3B A6 AD F0 29 54 49 56 19 B7 4F 36
 E4 E2 93 36 19 C0 FE 39 3F 3A 96 F7 F1 54 2F 06
 8F 36 CC 4A 3A D2 CE 69 3B 3D 4C E0 5C 87 DB AE
 E1 60 3F F1 BB 1E DB D4 76 C4 FD E0 B1 24 37 4A
 17 CE 96 D6 29 C4 60 89 6C CB 01 62 C3 46 B3 B3
 62 DD C0 4C 47 19 E0 3B 01 42 66 02 72 6E 7A 8E
 CB 05 15 C7 90 5D 2A 87 F8 3C F8 93 9C A7 79 CD
 61 CD AA 6B 1E 4F D5 84 B2 0D 33 44 C1 24 10 7D
 9B 77 3A E6 BA CF C5 CF 7E 96 32 A2 97 6B 7E DF
 ED DD 3C C5 18 11 C9 D1 0E 2C 0B 13 20 67 05 D3
 20 EA 55 E0 51 61 37 C5 5D 78 4B 97 7C E3 D6 48
 17 5A 47 9C D7 D5 35 A9 03 20 52 41 46 93 4B 5C
 98 54 61 F4 A1 32 C6 BC 8D E7 48 67 76 BB FC 5A
 E2 75 AD 5B 8F 9A C5 28 98 14 D2 5E 62 AC 44 10
 DD 09 68 2D EF 5A 5D 6C 26 1C 2E 1D 4F 63 3D 8F
 93 78 C2 66 25 EF FB 9F 62 DA 76 CE 10 02 F7 C4
 0F 31 84 AF 17 1B C2 86 88 76 BA 44 09 3D 35 43
 34 40 16 B5 CF 7E 1C A9 31 3C 76 84 13 77 70 57
 F9 51 5D DA 75 E7 6A 88 B8 3F 5F 21 F0 D6 04 06
 AF 78 29 B7 49 08 A3 60 31 96 EE 56 CB AF 8A D3
 9A A3 7B F7 D9 C2 C2 40 F8 77 C9 3D 0C 9A 65 28
 F4 CC 26 2F 02 00 89 3A 7C 99 F8 49 0E 35 97 1B
 58 A2 F2 A7 04 BA 01 21 2F CE 48 91 26 32 EA 85
 B2 47 EB 19 B9 93 67 55 58 C9 9E 15 33 70 21 DF
 2B 3E 4F B3 35 34 0E E8 64 7A 08 D0 75 33 61 F9
 35 B9 24 40 4E 0D 4E 12 A7 97 6B E3 D1 C5 2D 37
 54 FB 18 31 E8 42 F8 38 98 61 16 BB 3F BB BA 0F
 47 83 18 2A B7 DE 56 1C 12 02 E4 BA B6 E4 D4 0E
 0C 26 2B 85 95 0C A5 FB 66 E3 E1 5D 2F 80 BC 73
 7C CA AD 7E 32 BB DB 45 0E BE 75 82 16 63 15 5E
 70 D6 B4 30 65 73 99 36 6C BD CB 0D 15 3F B1 51
 20 F4 80 70 3C 64 31 A7 FE A8 D0 B2 DB 38 3B 20
 2E DB DD 89 F0 ED 94 51 CE 1B 10 01 C4 8C B6 4E
 01 9C C2 F7 FC 13 F4 B9 05 97 E0 63 95 62 76 BB
 4E F9 D1 98 76 A2 8B 01 1E FA 31 ED E7 6E 2E 56
 3B 35 67 9C 98 56 70 3A 71 A5 D1 BF 40 66 E7 C6
 75 9C 55 AA 42 64 C9 8B 35 D4 CA AB 73 9B 9F F6
 C0 4A 9F 21 1D 0B 93 EA 28 E9 70 DB 3A FE B8 F5
 7E 6A F8 16 DF E8 11 3A F9 8A 3E 70 E0 9E 67 3F
 B4 E7 77 4C 4B CB 90 73 08 10 D8 B0 3E 1B 12 D6
 06 31 72 6F 33 BD EB 5F 9C 07 B0 12 1E D4 65 8A
 A2 68 37 F6 F4 DC 0C BC CE 03 36 BF 87 EC D2 1D
 31 6E 17 25 06 2E C5 C2 9F B4 EB 34 AF E7 D1 70
 33 8D DC 1D 0C 0D 6E D5 70 97 D1 9A B7 BE 7F D9
 07 82 A4 AF ED C2 94 08 27 03 69 C4 E0 74 92 4C
 15 73 16 AA 29 EB 0E B7 E5 20 B1 69 98 55 5D CF
 AC 5B 91 27 F6 4D 32 FB 45 4A 91 5F FF 85 76 D3
 AB 34 AA 5D B0 6C 7B 6D 48 ED F8 C6 9B 26 69 D3
 D7 79 FC 1D AB E6 B7 78 12 F2 0C 12 49 7F 51 8B
 B4 49 4F 81 B5 2E EE 57 35 6E B5 A9 85 D2 88 D6
 5A 3E E0 49 6E 28 DD A5 5F B9 3C B8 16 B9 17 E7
 8D 75 50 F9 22 76 6C 1A F0 25 8F A8 2C 0F 69 42
 0D 53 EB 6C A7 68 80 BB 6E E6 0A 77 94 C4 AC 70
 9D 0E 6C 60 32 D8 C5 02 8E 32 ED 08 ED BD 57 8D
 F9 CF 42 16 97 1B 69 BE 78 20 FC A4 2C 98 5F B3
 18 51 4B 72 91 EE BE 72 18 39 9A 5D E3 34 60 D7
 6A 35 32 30 1E 87 3C 1C 2A 75 4D 66 4C 88 33 BF
 F2 0B 9F CC 5D 3A BA C3 29 1E 30 D5 22 6F C1 83
 31 67 FD 8F 7C 05 B8 BA AE 8F BE DB 07 C7 BE CD
 1B F5 E9 96 E9 4B 84 E5 68 9A A8 3C 31 52 0F 75
 22 F0 38 64 AC 7F 03 2D 6B 9F EC 0F 97 30 F9 0C
 C2 50 41 66 45 AC C2 03 63 BE BF 36 64 79 FC 69
 ED 48 5C D3 13 E9 53 86 70 DE 79 6E 49 80 AD 9C
 7D A2 5E F5 1C A1 AD 38 3F C5 4B E5 88 CA C8 B3
 95 5C 07 0A 8D 8C 5C EA 50 1E B4 D8 8C D9 72 BA
 1C D3 F3 E4 64 2D B5 77 AB 05 B2 1B 08 AF EB FD
 1A DE B4 40 98 FA E3 48 8F 54 88 D2 B9 CC 02 7D
 1E A3 E3 3C 22 0F CC C7 E8 92 FE F0 74 B3 5F 3E
 F3 58 4F 05 82 75 B4 35 48 B3 26 80 F2 9F 60 CF
 C2 CE 1B A4 ED 3C 30 C1 33 7A 97 65 9C 22 DF AD
 66 48 0E 62 82 A0 75 D5 1B 50 56 A6 7D 8F A1 FB
 39 70 11 A8 71 8E B7 55 04 49 E9 E4 CC 50 F8 E9
 79 AE 72 4E D0 5C 81 45 44 A4 58 24 1E 14 16 D1
 9B 6B C6 B5 44 73 62 CF A6 7E 26 EE 45 63 35 78
 33 87 EA 30 30 51 55 37 CA 67 34 29 0B 47 E0 B1
 2F AD 08 3C 4D 41 0C 8A 4C 8B 5F B5 7D 73 E9 22
 06 08 BB FD D7 5F 1A D2 02 5D 6A 4A B2 47 6B 84
 D7 1F AC 89 D1 DD 60 9A 1F B9 B6 E2 05 6A D0 B3
 16 85 25 75 74 5E 43 A9 51 BB F3 BF 80 D5 DB 22
 B6 DF 97 1D 84 EF 18 11 9C 8B 99 ED 2D 7A 4E 63
 A3 AC E3 DC 68 86 70 C1 5B 90 89 16 2B BF 17 46
 07 E4 62 09 36 09 60 27 94 A7 A8 C0 E3 49 28 1A
 43 88 A2 6F D8 7C 25 0B FE AE 03 BE 23 94 2C A2
 95 C8 11 DE 05 54 4F 3B 28 D4 0A 0F 23 77 C3 0D
 50 3D 1B 0D 91 54 60 5A 13 5D 56 A7 0C 90 6A 7F
 33 2B 38 CD 9E 49 B9 73 1A 61 37 5D 55 26 7B 2A
 7A F0 24 02 2C 7F 61 6C 9E D2 A9 37 AA FA 2A 84
 BD B9 8E 4E 96 CA 97 65 57 4E 17 78 13 50 59 60
 EE 32 65 6C CF 6A D0 49 21 A0 65 E7 79 7C 82 77
 2A 0B 92 9D 83 1E 00 40 99 D7 76 44 11 38 26 C4
 CE 53 93 38 48 61 B4 55 79 BF FB 45 1B 0B 3C 6C
 E2 3A 07 F5 A3 1D 36 B4 F8 F8 E6 ED B7 EC AA 1A
 2C FF 5A E6 16 AE 68 3E 53 B9 2D 06 4E DD 55 DD
 D1 12 E5 A2 A4 73 C7 5E D6 F5 5D BC 3C 25 A3 6C
 F3 2C 5C FE 8E E0 96 5B 81 83 A8 C4 AB 91 02 6A
 5B 01 84 36 0E 82 8D 92 F0 40 D2 25 F5 70 6E A4
 98 74 8D 60 71 2E C7 25 6F B2 51 00 9A 1C B8 DB
 B0 C5 98 FA 53 56 C8 96 02 1E E4 9A 86 DD E2 F5
 8F 3F 18 88 A4 8C A7 8D 6B A3 E3 58 F2 A6 30 3F
 63 5B FE C2 49 87 75 E4 31 EA FF 67 FE 9D B5 7C
 D4 54 D1 F4 89 76 91 A1 92 FE BA F9 2C 62 B1 D5
 24 BB 57 C6 DF 02 A1 50 B1 3B F0 BD 0F E3 E5 DA
 E9 E7 08 47 30 00 47 F3 79 DA C9 39 AE A9 A8 CC
 4C D2 FC 41 CA 01 EC A9 69 CE C6 1F 28 7E 93 20
 BB 94 24 AA 98 1B 45 9D 39 31 0E E4 A4 44 DF 8D
 F0 E4 26 D0 CE 2C 5D 9C DF F3 47 C7 43 10 D0 29
 74 8E 48 A6 56 CC EC 24 F0 42 F4 C2 90 F0 55 D1
 56 BB AB F9 77 09 0D 1E 5C 17 3C 5F EF 0E 96 19
 90 2B 9E 00 E6 1F 59 EC E4 97 CC 36 BF FB 86 CB
 1C 5D C9 8F 11 0F D6 B3 F1 50 15 DB 10 2F 9E EC
 41 C7 C3 67 2D C3 BD ED 79 71 1C CE 9B 4C 0C A1
 DA 1A 2E 93 9B 48 67 02 EA B4 DC D7 50 A3 18 3E
 30 FC 0B EC 05 C3 23 36 99 F5 3C 15 EA 84 FF D3
 1E A6 0D EC E5 12 F3 BF 4C 13 DA 21 7B 8C 54 3F
 CF AA AC 1B 93 45 17 98 DB D0 E4 36 12 D1 CB 89
 E4 3B 29 1D 23 B7 C5 55 33 68 6B 8F 0E 3C BE 05
 EE 01 D3 45 DA 4D 8E 94 6F 21 26 ED 9D 02 5C 28
 08 FA A0 77 D8 88 D8 CC C2 EB B1 EF 7E 7E 84 7D
 B4 3E 99 7D 09 0E 77 66 93 AD D9 37 7B 2C 81 4E
 AE 25 D7 CE 6E 39 8A C5 87 BB 45 1F CD 53 D9 64
 02 92 1E C8 59 48 BF 24 48 78 3F 90 59 DF BA 02
 AE 81 32 41 58 A6 E8 B6 D5 2D 5B 86 54 85 5B 2C
 F9 9E 98 4A BE 64 4E B6 4B 0B F0 34 D6 77 6E 5B
 48 BC BD 3D CC 35 C9 C3 F6 2A F6 37 00 EC 98 65
 B7 BC 70 20 D2 CB A0 9F 39 7A 13 6E 2B CE 75 19
 38 6C 29 EB D2 A0 E6 A1 C4 0F 41 F2 C5 C8 5E FB
 5F E2 98 D7 FB C5 F7 EF CE 72 90 AC 9B E1 EF F2
 92 08 58 9A 0B D4 83 55 22 D0 21 4A 23 ED 3F 8F
 30 E3 0D 5E 11 04 8C 6C C3 B0 43 97 D4 2C 3E CE
 8D 57 43 F1 6E E1 6C B0 58 25 1C 03 FA DC FE 6E
 A6 30 D6 CE BE A4 DB FC BE 8A 37 DA 98 91 2B F6
 4E 27 AC 4B 39 17 D8 B9 E9 D0 2B C1 23 46 4F AC
 FD 51 72 98 B1 C4 FF 79 6E 49 0C 19 C0 D9 40 F1
 34 85 E8 F7 6A 0E 91 D6 00 42 00 26 39 5D 95 48
 4D 1C 1D B2 7D E6 DC D6 00 E6 3F 0E C9 B4 44 77
 3B C7 3A 19 66 9E 4E FC 49 E5 A0 52 7E C8 5A 00
 75 17 7B 27 67 3D BF 16 15 74 00 A2 FD 25 8B 21
 6A 49 B4 28 9A BE CE 6F 31 5F C6 04 EC 4A DF 07
 3F 4A E6 A9 1E 03 73 55 1F 04 94 4E CE 0E B8 CE
 32 07 38 9F AA 36 A4 C0 EB 8B B4 5D 08 B7 D0 CF
 A2 B9 22 DF 8E 2A 04 EF EB 3B 0B 89 B2 B0 9D 6C
 E2 A6 1E AD 85 AB 09 8E 30 3D EC 6F DE 5C A8 39
 80 26 56 05 02 0A 32 8F 68 34 23 56 4B 42 BC 09
 4C 2E 94 52 BE B4 85 E3 3D 90 BD 90 13 D0 65 7C
 D4 23 70 36 00 AC 8D 5A D4 78 17 96 E1 F0 50 08
 31 46 E1 9D 6C 76 1B 75 3A F8 51 17 00 1A F0 37
 04 97 5E DA 8C 54 24 AB 8B 15 F3 6F 12 0B 16 D1
 2D 6B 0F DE F3 1E F8 5F C3 1F 30 2A 55 70 E5 96
 0C EB 5D D0 57 91 23 D3 53 B2 EB 5D C9 29 3E A2
 87 7D A0 64 00 79 B3 1F A6 CC FB E9 97 F0 26 78
 E3 02 28 E8 D2 05 F3 A1 EA C8 3E DD D2 A7 5E 01
 36 48 7D CD A3 E2 E3 48 66 3E C3 69 A2 BA 42 17
 C9 FC DF F7 74 39 23 9D 22 B4 D0 5B 77 B5 DC F5
 93 BA 63 FD E5 3A DE 5F 52 0B 49 93 6A 22 89 19
 8A 8F C7 5D F8 96 71 AD 1F 3C 72 C0 FA 83 FE DF
 6A C2 11 0C EB 09 92 00 7C 92 0C 28 08 3D 46 0D
 D0 EE 35 DA 44 CC 19 21 2F 1E 54 8F 74 36 0B 14
 22 54 88 C6 AF BE 1D 3D 6E 8D 7B 9B F5 29 7C FD
 44 2E 03 B1 16 9D 79 B5 4E 82 56 D0 DD FE 1C A9
 60 42 0A DE 20 26 FA A5 B8 D5 9F 25 5A 40 5D FE
 22 5D C4 D9 4C CF 0F D1 3A 78 34 A0 B7 FC AA 42
 39 DA A7 03 86 14 B9 D8 C6 11 22 17 57 87 5D 47
 A3 92 DD AE BF E1 6F A5 FA A4 B8 DF 7D 05 EC 71
 7C 1C 0B D1 2A 12 DB 48 3C 2D 07 DD 54 91 A1 4F
 BC 46 E1 18 9D 4E 0B 25 E3 D3 5A 9A 35 9D EC 10
 79 81 28 D7 78 8E BD 20 3D 72 90 45 98 22 63 8D
 C2 68 EC 30 ED 9F E4 24 25 4A DC 96 36 2E E6 2C
 5A 4E 54 39 ED BD 8B 6A 14 19 7E 4F 5E 32 A4 65
 3E B1 BE 38 A3 91 5A 71 E2 AD EE 0B 09 3B D3 1B
 E6 A2 69 F1 5F 73 36 73 02 67 09 20 55 64 03 25
 3D 45 5C 5E 6C DB E8 74 2C 81 D6 AA F1 F1 FC C9
 22 FE 7A 0E 61 61 7C AE 31 11 90 88 60 64 95 E3
 5F C7 5F 94 E4 EC D4 D4 D6 CC 27 B2 E8 2D 8C 86
 AF 0F F1 3A 64 C1 DC 70 CF B7 26 0C 7E 86 22 60
 11 F0 D4 7E 6B E6 83 97 8B D7 C9 53 70 5C 1C D1
 BF 82 E5 4C 69 E9 B4 51 62 45 97 E7 21 D9 CB 9A
 EF F6 A7 E3 E1 26 3B CA DB DA F0 40 B7 16 B9 EA
 AE 77 5B 86 CB DF A4 8D 84 4C 54 F2 24 62 8E 28
 DB B5 EC 4D B1 A4 9D 7B A8 94 E6 39 81 21 83 B4
 3E A2 94 E7 B8 D2 4D 11 ED 48 AE 2E 38 06 E7 DC
 D1 C3 EB A0 83 D1 A8 51 82 3E 81 C2 80 78 84 29
 9B FC 28 05 CE 43 E5 DD 4C 5F D5 38 D4 33 D1 BE
 F5 2E C9 F6 09 5C A1 14 5D 22 D0 6C CF 77 E2 BB
 64 11 26 80 85 7A 5B 0D 07 13 8E 09 2E 2A BF F0
 A1 30 39 2F 49 03 92 EA 15 D7 E7 19 AC A8 F3 C8
 FD 2D 6C 20 26 EF E5 24 57 BA 45 8E 1E 07 15 18
 DC 72 90 F5 BE 2C 24 56 F3 CA 8B BA 20 CB 7E F5
 42 73 80 A6 02 69 E9 AE 7E F8 4D E2 94 FD 19 3C
 96 D2 FF 5C 78 87 B0 A0 1B BE 30 7E FB 16 29 D5
 54 31 8B 2F A8 41 51 43 F2 74 40 81 79 31 C4 C6
 45 86 D4 A1 9F 46 26 7F E2 43 0E D2 3D 5A 40 F0
 07 4F B6 4B 7B 70 F8 07 B8 4C C4 18 DB D7 C1 AD
 E3 F9 73 D9 3B 4A 88 16 9E 51 00 BF 2F 15 0E C1
 D4 A2 55 FE F5 8C 88 B8 65 D3 24 6F 87 11 1D 4D
 DF 82 E2 82 2C A9 AC A5 F7 C9 8F 35 05 F1 69 93
 4A 38 25 EB EA 68 12 BD C9 73 C3 2A 17 1C E1 6F
 4A 52 86 EC 20 94 4D 1D 70 2F 8C BC EC 74 5F E6
 D3 40 EE 92 C6 46 5C 2A 83 E8 F1 09 8C 47 74 76
 86 63 08 9D BB 47 E2 F1 1A 88 30 BA 37 8F D3 52
 C7 0A 86 A9 3B 00 75 C3 1C 2E 9F 2A E8 AA 04 D0
 00 6F 93 B5 21 03 AE A2 9F 5E 7F E2 28 01 EE 61
 DE 4B E4 B5 58 A5 11 DC 3C F3 BB E8 94 F0 40 FB
 6E F3 62 09 F0 D8 27 EF 53 9D 8A 08 DE 78 7F D8
 CE 84 97 80 0F CF 39 20 43 6D F1 27 11 08 95 41
 99 B9 B7 3C AE 98 2D 4F D8 68 A7 E3 4E 25 65 C0
 4B A8 E4 D3 76 84 48 8A B8 36 AA BF 8B AC 3C 76
 73 48 9C 56 19 B9 6F 4D 7E A2 DC 64 79 EF 43 DD
 09 10 17 D1 5A 52 89 40 26 AD 95 7A 8D 0A 8E FB
 67 A5 A4 7E 7F 99 A5 27 DB 35 54 1B F1 95 88 3B
 2C 5A F0 7D 0B A0 69 86 BA B7 01 64 5D 0C 9C 96
 1E 7E 3B F9 F5 C0 52 7A ED DA CE C5 45 B4 7D F8
 E2 98 F4 25 06 D7 74 4B E9 9D 7F 51 83 15 EA 1C
 82 C2 8D 10 40 10 49 6F A3 5D F2 67 D5 BF 82 66
 7B 9B A6 AD 30 F7 76 0F 39 23 11 76 ED 87 FF DD
 A4 DF 44 06 BB DF 83 74 4C 5A 7C 7A F0 6F C8 8E
 20 AA 2A 14 E9 A3 00 EE 68 18 F1 85 9C 18 68 AB
 93 F6 62 BA 63 97 4D A3 C7 37 A4 C3 66 57 E0 51
 1D 12 0F D1 6F CF A2 C9 7E 57 87 54 BB 87 A2 A0
 6C 35 98 7A 9C 72 76 91 1F 18 9F 10 26 4C 1B 1F
 2D 26 66 68 C1 45 8E 0E AE C2 E5 F2 2B C0 C9 51
 AF CF 3D 17 43 AF F5 C2 E6 52 E4 D0 BE 59 26 E1
 B8 AF 59 79 CC A7 F7 EE 54 46 A0 57 80 69 B2 99
 5B A6 9C 7C F9 B8 65 C8 81 28 BC 58 82 3D 03 1D
 8F 23 13 F1 3F 98 31 9E 84 00 D9 01 C7 C4 7C 92
 C1 AF 73 B3 4B CF BD C4 28 38 29 CA 67 B6 83 42
 09 52 39 87 03 83 C2 60 B4 9C 6C E2 9B B9 AD 16
 DC FE A9 EA 76 28 D7 59 87 03 19 43 03 3B B4 7C
 7E 32 5F 6E BE 1E 6B F1 3F 05 AF 38 9F B4 6D 2C
 51 1F BC F2 10 3E E6 61 C6 C3 89 A5 FB F5 9E 35
 1B 31 E3 0C 3F 33 FD 1D A9 BB 3E F5 BD AF FB CA
 81 6F F4 57 8F 9A E2 F6 E0 40 20 1A 55 6E B0 2C
 85 FD 6A 78 D3 7D B3 43 8A 52 01 01 34 BD A0 1A
 75 F0 54 5D 4B DC 41 39 F5 F1 1D D9 D0 42 41 43
 FE BD 16 48 3A 35 E2 30 71 A7 88 C1 9D 51 0D 93
 28 BE 85 CC 55 D5 A2 FE AE A4 0D 5B BB 41 1B 8C
 77 E9 74 18 1D 6D 50 3B FA BC C4 A2 02 77 27 41
 20 01 69 8D 22 A8 EE DD D5 82 CD 4E EC 34 49 63
 00 8B 86 0E A4 93 32 10 19 16 10 C0 A2 5F A0 C6
 A8 14 6D 28 53 78 77 DE 1E 7A 55 64 C5 D0 3C C8
 22 90 C0 84 51 46 41 CE 18 A7 0F 84 99 B0 FE 96
 C5 E4 DE 15 A6 88 F8 79 ED F7 8F 54 B0 84 4A 07
 06 AB 6D 2C 03 CD 6A 57 5C AB 2E B1 0D CC 62 DA
 77 76 20 EC 17 A8 F5 E1 04 BB DE D8 40 16 8F DA
 B5 2B BC A5 D8 35 F8 AF 5D 87 D8 EA 08 B6 A6 23
 61 3D 1E 9B C9 46 0D 58 31 17 3F B9 ED 02 89 64
 07 2F 83 C6 0A 9E F9 CC 17 6F 0F DB FD 77 30 ED
 BA 0B B2 83 15 43 26 0F FE 44 19 EF EF A6 E9 45
 A9 0A 80 5F 64 CE E8 00 88 45 CC CE E7 0C E3 90
 89 2B 7D 15 8A 45 90 16 1E 70 67 65 22 F9 17 78
 58 99 D9 61 28 AC 2D E1 1D 0D 8D 98 7E 30 A6 7D
 7B 84 C8 03 F7 BB 26 BD 4F E9 FE 79 47 27 65 CE
 99 F7 DB 9E E2 70 51 C2 8B F5 64 32 C3 86 D8 93
 6F DB 96 CB 33 7D F3 FE 8D 47 CE 66 AC D6 AD 0C
 52 A0 8F 26 9E 35 3C D0 7A 22 2A D4 1F 55 EF 88
 94 B9 8E 38 37 65 D7 F9 AA 43 9A B8 9C 2F 29 EB
 52 78 72 F1 11 29 A3 FA 93 A1 6D 00 12 FF 8D 0F
 7E 1B 2A 96 9C 2C 56 94 7D 86 AC 6C AE 98 90 27
 30 4C 45 A7 46 60 83 5A 6D C3 DE 29 F1 7F D5 3C
 EF 5C 26 88 57 71 23 73 10 9C 95 F6 BE 68 51 F1
 81 D3 21 6F 7F 8B 49 35 A5 58 F7 D3 84 14 AE 79
 8B 75 A5 32 78 14 09 17 B2 68 DC D1 3B D3 B9 F2
 A8 E1 63 AD D8 FF 8B 50 7E E6 57 BB A5 E8 61 DE
 09 ED 5B 29 9F AE E6 ED B9 F6 97 3C 7E 32 49 7D
 6B 68 7D 81 C2 0D 30 70 C7 BB 26 30 C6 50 AD AF
 87 D7 F5 7D 82 03 39 44 B5 46 8E DF E1 20 D6 7C
 CC 47 5C 40 3E 2A 38 8E 1E AD FB C8 A5 1D E3 35
 6F 4B E0 5A 24 B9 CC 62 0F 72 DE EB 76 4F 83 29
 45 30 35 33 49 BC 67 A2 9C 5F 16 38 59 78 40 E1
 DD 0B F4 B9 B9 7F 3F 51 CB 97 13 B4 0A 28 5D 99
 15 14 1E C5 0F 22 9F 03 AD 66 DF 0A 32 6C 9F 75
 FA 02 9B 53 28 EF 3B AB 2F 7E 31 4B 8D 37 82 BF
 C5 10 4B AB 82 81 69 3D 1B 37 23 6A 71 3C C7 51
 2B 6B 71 07 60 64 32 19 8E 0C 68 ED EE 28 B0 08
 D0 BC BA 38 18 76 38 DC 37 5F 35 03 EA 7B BB 1B
 18 2A A3 0F E6 04 F7 41 15 E7 EC 0F AE D1 37 89
 8E 5D 05 68 46 41 2E F1 4F 0F 16 D4 ED 95 AF B7
 37 F0 48 30 A0 28 B9 E5 0E 62 5E 15 98 18 A4 BE
 EC 35 A8 63 A0 00 73 87 AE EC F4 41 66 2C 40 D0
 D6 40 4B 4E 09 8D 36 3C 54 43 42 40 83 5B 31 41
 A3 62 0E E3 06 04 58 AF 28 66 06 9A 7C 24 73 22
 CC D8 1F 1C B0 80 27 39 1C CA B5 21 4C 30 85 53
 34 56 29 26 37 32 13 E0 A2 2C 49 D1 93 F0 03 9D
 C0 99 A9 98 EB 69 25 F4 09 8D 6F 23 E5 DC 82 1A
 FD 03 E3 46 F8 C3 D1 C5 69 CF 76 94 76 C8 E9 BD
 78 CD 97 4A D4 B9 DA CB D5 4A B3 C4 1E 73 67 78
 9D B5 A2 71 31 82 F6 B9 76 94 34 74 09 53 29 1F
 EC 3F 38 31 17 05 90 4F BF 53 75 CF A7 34 BD 07
 0B 5A 00 D7 96 56 0A 02 0F 5B 19 A4 13 DF D5 61
 CF 3D 5C BD CA 1C 31 C0 82 6A 9A 52 AC 13 87 23
 B8 BD 0E B3 E4 8C 9A F9 FE 3C DC 83 3A 55 58 69
 42 DC 20 9E 1F 58 76 B7 D8 4D A1 37 38 4D 94 57
 82 1B 4A F3 67 53 06 98 B3 24 6E 33 30 D9 C1 86
 44 CE A6 9F 07 67 C5 ED DA 53 83 30 A6 D1 CD 4C
 89 AD 07 A1 C8 0C 90 93 E9 E5 14 A7 21 F3 76 04
 6C 48 72 25 08 D3 88 91 3A DC 0A 74 EC 06 41 1E
 38 EA 2A 9C 9F F5 B6 C5 45 1D 1F 2B 56 BA 65 BB
 62 B5 5F 65 3C 7F 52 6C 47 AA 8D 72 8B 4C 65 21
 77 CA 52 0E D1 C6 5D 2C 8A A5 9E BC 79 2D 42 64
 0E A4 FD 42 07 9A 56 AF 74 72 BC 8E 2A 68 B6 38
 2A CD EF BE 19 15 95 2E 08 82 5F 9C AB CA B4 BD
 BC EF E5 74 F5 E6 CE C1 45 97 67 9D 79 72 FB CD
 5C 43 CD D2 5F 03 18 B2 EF 03 2E BF CB 68 96 D8
 2F 1D 25 CD 30 13 AA 5A 77 69 7D D7 24 E8 AE FC
 8B 83 58 A7 F0 32 26 3E 15 92 86 B4 1E 9C 2E BF
 5F D8 51 84 57 2D 34 66 49 92 C1 ED F0 85 EE C1
 33 F1 40 13 CF ED 2B F1 1E CE 15 22 47 88 E1 5B
 4B 4A 09 B1 36 B6 9D 3F B6 AE 57 AE F9 D3 78 22
 3B 6D 93 B9 F1 C1 A6 65 39 13 33 5C CC 86 85 4E
 42 52 2C 67 90 AE 62 D3 5C A0 3E B6 1E B1 2B FE
 BA E2 06 08 97 75 31 07 B6 D9 29 C1 31 A2 C7 3D
 6C FF C7 46 9B 90 3E 61 ED 1C 5A F6 B2 9E 49 F2
 22 75 4E 18 F2 68 12 EB 19 E3 60 35 B0 BC 76 73
 55 2D D7 99 31 3E 17 1D DA E5 85 4F ED 4D E8 E6
 EA FB 1A 4D C9 D0 28 94 A0 49 FC 58 C0 83 0F EE
 CD 4C B0 7C 93 58 E6 54 C6 B7 6B 31 E1 FB ED 90
 77 E4 35 42 11 8E BD B3 7C 27 AC 3F 1A 5F 85 0F
 A6 08 45 E2 3E 7F 01 FF 3B 5C E0 38 83 47 C4 B7
 F7 F5 27 59 55 2B 34 E3 C3 C8 42 55 1D C3 61 14
 AB 59 E9 A2 17 BD 90 B6 FD CD 8C C6 E0 4C B9 E5
 24 16 70 5A CA 76 2E AE CB F6 7F B2 A2 74 B1 51
 38 45 6B CF 36 65 A6 65 BD ED 1E E7 B1 72 98 8A
 5F 6B ED E9 96 C7 24 52 7E D9 E3 6F 06 D9 6E 2B
 42 9A 72 45 84 07 0D CE 28 51 01 B2 78 23 D4 40
 49 F7 D4 5F DA B4 7F 18 FD 74 5C 56 BB BC 07 29
 C2 80 FD F7 E0 9D 78 C6 F2 41 11 B5 25 26 28 19
 61 5F D3 A6 3A 9B 70 85 B8 B9 0D 98 5B 56 CC 0C
 F5 08 8A 2B 51 F3 01 75 69 57 1B 47 1D 2F C4 AC
 67 D7 FF FB 53 CE 36 47 96 CD A1 25 35 AA 65 A3
 D4 6D 36 C2 2F 98 1C A7 11 CB EF 70 98 BA 2F 01
 F5 69 AC 72 98 FE BC 59 AC D5 6A 9E 29 F9 03 5B
 2A 8C C6 06 08 D2 86 AB B3 B7 2C 12 88 01 85 50
 8D A6 8D 73 24 D5 DC 19 27 CB 00 9F 39 1B 4A CE
 E9 25 AD 98 EB E9 98 26 7C 29 51 F1 E3 41 03 AB
 E1 25 19 18 01 A7 CD AC A6 1B F1 91 BB 1C CE 15
 56 B1 04 7D 40 51 DE CE F2 64 69 43 E4 EB AD 78
 1D 5D 2E 2B A5 23 3D F6 63 FB C4 50 0F 46 CA 52
 7E 9F 46 E5 30 C6 1A BC 4A 14 EC 35 9C 99 81 93
 0B 59 91 24 21 11 AB F9 63 D5 8C 78 BE FB 98 7A
 0D 5C 7C 7A C2 9C F6 CE E3 38 25 FF CB 40 41 19
 8B FE 32 30 B2 9D CA 1E 9E ED D3 74 44 F7 32 69
 1C 58 7B A0 54 2E 93 4A F3 4F C1 E2 44 2F 2E FD
 E5 9D A4 42 2C 36 42 84 13 2F 05 9E 21 05 ED 15
 66 B8 C5 49 3D 9F 17 62 ED B4 C6 12 B6 E1 66 2C
 67 51 07 23 C1 43 88 2C 92 10 4E D2 4E 9A 4A D6
 E9 F8 9D 3C D3 44 57 CF 13 92 58 E7 31 A3 7F 7E
 21 13 34 72 E9 B4 C4 49 2A 68 87 D2 80 57 2B A1
 D4 09 53 F1 AA 3C 31 46 04 79 EE 78 C5 DB EB 82
 A0 5C 07 3F 6F 7F 70 73 DC 99 0E 7D 1D E1 0E 20
 16 01 40 A7 03 08 49 54 E7 68 23 47 DF 3D 5B 64
 B0 BF 6F 3D 8F 3E 2A 19 D5 FE E0 DD 46 69 97 6A
 D3 00 DD 0C 1F E6 6D 2C 64 01 ED 56 98 0B FA 7F
 24 4F 80 8C 9D 44 05 16 41 12 90 74 E9 77 F4 78
 8E DC BD 35 3E 78 EA C3 FB 1E 75 D7 00 D4 A7 99
 FE 32 6D 96 93 2D 49 39 78 EB 46 51 50 35 8D 3A
 6F FD 4F 54 58 EF 0A 5E 21 E7 B8 86 BE 47 DB FE
 0C 65 4B 4B A7 99 EE 0D AE 8A 2B D8 DE CA B9 42
 91 70 31 81 43 C1 A1 07 E5 50 95 C7 4F EA D4 AC
 1D 73 30 1C A1 61 F4 EF 86 B8 41 71 AE 96 5E DC
 8F 3B A4 AE 4C F7 72 DA 2A 04 07 AD 66 D6 28 9F
 3F 09 8E 93 5B 1F 3C 86 20 48 C5 B7 76 6A D5 DB
 C3 CC 4A 27 1E CF B6 D0 3A 79 E0 AF 32 68 68 27
 A7 A2 2B F2 CF 4B F7 DA 76 B4 FD DA 3C 00 43 AA
 AD 4B 42 3A F4 67 66 97 7B 01 9C 78 3F D3 45 14
 B0 22 1C 43 EA 32 C3 58 81 02 F7 DC 16 97 4D 88
 F5 CB 73 50 5C 0D 7A 4A F6 1E B3 D5 8E AA C6 D0
 88 A8 68 55 3E 40 73 B0 24 03 95 31 46 CE 37 CA
 67 AD D1 CD CE 75 E6 91 01 97 15 35 49 50 7F CC
 8F 29 4A AE A9 1E 73 31 7C B6 DE DC 44 46 C4 28
 C9 FA 0E 15 EE 4E 9A A5 04 09 BB 9C AF 30 3A A7
 42 81 20 9A 6A 76 CF E5 9A 6F B8 CD 36 FE 9B 1E
 64 AF 6D 50 0E 82 BF FB DF 13 33 85 2C 8F 6A 0E
 E6 DB F9 31 2C F1 5A 75 98 01 0A C0 00 11 4C 89
 57 09 AA E4 03 FB BD 78 1A 42 6F DC C7 F2 8C C8
 68 E0 B2 04 5C 7B 1D 4A A6 81 09 FA AD 73 9A 9A
 FF F3 3B 18 E6 B2 C2 F7 74 9A 14 33 3F 94 39 59
 21 81 DF A2 82 CB AD D5 74 AF 97 B9 D4 D3 13 36
 8A 61 D4 98 63 26 60 F8 D1 71 05 04 DF 0C C4 99
 C0 3B 2E C4 9E 4F E0 BF DB 5E D9 53 FF ED F0 65
 E0 38 26 BE 47 FD 5D F4 C3 9A B3 71 68 7D 63 7E
 70 2A D3 0F 10 FE 33 2F D4 E7 34 17 77 E2 93 22
 8C E5 23 1C 0D 31 34 E4 18 DA D5 F8 4D 92 EE 8D
 8E F2 94 06 5F EA EB B3 C0 A7 2C E9 B0 00 4D 65
 82 A9 43 54 07 F8 D4 36 15 69 61 E6 2C 96 F7 E2
 F1 7C CB 40 41 CD 61 DC 35 16 BF 90 C4 37 30 B9
 A6 37 84 2E 90 4B 89 41 A7 4C 70 5A 74 B8 DF D0
 31 27 D7 B5 FF 7F CF D4 9D EB C6 3E 10 83 F8 D2
 BF C6 35 86 DB 9D 15 38 50 81 79 1C 53 7B 6B 48
 11 E8 E0 C1 7A 9F 6E 71 B0 13 43 57 16 11 5D 73
 AE D5 23 2A 2E 3D F6 9B 7F 64 F7 B5 69 5F D6 12
 2E 06 B9 BA 72 F4 59 C7 75 9B D0 2C 0B 92 B1 C3
 46 48 15 D3 6B BB 81 F8 AA AC 9A 56 98 DB E0 2A
 0E B9 0C 28 D8 5D 5C AB 20 B3 E9 9A 1A CC 23 EB
 AD A6 B9 AF 8E BA 8F DD 1F 41 97 3F 93 E2 32 7E
 0E D3 6B 46 D6 16 5C 54 E0 35 05 F2 26 D5 B9 90
 E8 68 BF CA 59 A0 E0 58 24 B2 95 C6 0C 1C 59 58
 CD B3 47 3F ED 89 B5 23 D1 01 64 1A 97 F7 4B 36
 09 D6 68 1B B9 CF 09 FD C7 4B F6 D5 EA 5B 30 B8
 9A 2A 46 88 CC 0C 63 56 AF 72 78 13 32 FE F4 C9
 E9 BD 35 FF 31 24 A6 FA E2 14 5F 7C 2D 7D 64 6A
 B4 43 8D 10 8A 3B E3 C6 35 85 67 C0 E6 93 5F 35
 04 4F CF 51 2D 9A 46 83 54 10 5C 7D 8D 93 CB 82
 F2 07 BC 16 10 29 58 97 6B 1A 12 E2 28 24 A7 CE
 D6 E7 E0 8E 34 38 63 17 CC 97 A7 43 9D 02 CE 3E
 52 EA 43 34 64 E0 27 85 37 6D FD 58 7B 31 D5 03
 6D 9F 23 77 6F 34 48 AD 70 A3 D4 6E A0 23 22 70
 42 6F 46 88 5F 45 1B 4F 7E DF EE B6 04 3A DB 6E
 D1 58 2B DC B2 F4 19 F9 5E A4 BA B0 7A 90 E9 D7
 FB B8 14 D4 96 92 5B 6E AC 1A FA 30 4C BC 4F 7C
 55 B8 11 51 27 AC 21 5B 1E CA BA 36 2A 3A 22 F7
 84 57 DF 7D CA E8 91 A3 D7 72 1A 3A 9A 34 84 66
 FC 77 9D 18 77 90 26 B9 54 80 C0 B1 6D 44 61 F5
 CE 26 63 A6 3F 2A 13 E7 88 71 3E 50 9B 71 12 EB
 4F 3B 20 F6 2F D3 75 FD 54 B2 EA 84 04 9C FE 48
 A3 15 12 E4 FE A6 CD 5D 40 F2 53 03 F2 9B A7 93
 28 87 49 4C A1 D4 B3 EC 9A DB D6 64 05 FC E7 0B
 C2 4E 4B DA B0 4F 57 CE 14 9E F6 25 16 46 90 E9
 8A 13 C7 AE E4 32 27 1B DB D7 B9 38 F5 D0 5B 36
 FA 7B 29 D2 79 C5 6F 0B EF FE 9B 67 61 42 47 79
 BD 47 30 7C E5 6A 11 DA FD 18 B0 F4 7A 00 5F 37
 DF 01 16 9B AF 51 42 78 DB 8B 39 AC 4C 86 9C 57
 FD 77 72 74 3E 7B B6 01 2A 4C 6C C5 08 E3 4E 80
 A4 9A 42 9F 66 23 6B 6A E9 60 A2 1E 76 D3 8A 6D
 DE 62 8E DA 93 A4 A4 6D 1A 16 7A 9F 84 BB B7 04
 7E 86 A6 AD 84 AF 22 F2 65 4E 77 2B EC 6F 37 EC
 3A E3 9E 8B 41 AD 84 0A D2 7E B7 A2 FF 51 1D D6
 FE C7 FC CD DA 91 FA BC EA 16 F3 9F A9 50 50 10
 16 CB 19 A5 21 C0 D8 93 CC 27 AE 93 8D 8A EF A5
 BF 3B AE B6 FD 99 A5 55 C8 37 F8 0D 96 3F 8B 94
 78 72 07 59 27 07 21 C5 C4 FA BF 84 93 07 BA F9
 84 20 01 5F DF 8A 45 C2 DF 95 C9 63 67 90 4A F9
 F1 54 2F F7 A7 91 56 5D C7 5E 1A 6C FA 9F 05 C7
 34 22 73 59 8A D9 8F A6 16 83 17 0E C9 EB B9 62
 91 71 DF 77 5E 66 11 01 13 AD 66 C2 8A B4 33 38
 43 B0 48 7B A8 99 A0 4E 95 55 13 C4 1A 03 5E BB
 50 ED 85 3B A7 73 85 FC 0C 28 83 0F 7D 5D 00 8C
 38 18 F0 6E D6 FD D6 E3 C6 35 00 CC C9 B3 FA 92
 72 9D BA 6B 5E 21 8B 0C E6 58 C8 26 CF 51 6C 20
 66 80 DD 39 5F 06 3D 1D EA 52 C0 AB 91 80 B0 A8
 16 D2 5E A6 74 BA 9C A4 09 9C 08 75 F3 75 37 5E
 AA DB C4 2E 6C 13 A4 C2 6A 07 E8 10 8E BA 82 23
 E0 72 DC 8E AC 80 D2 E1 ED 49 B8 23 BA 17 29 FE
 A3 6F 82 C7 95 B3 E7 39 D4 27 88 A5 AA 80 5D FF
 CB 15 42 27 46 12 95 C5 2E 35 F9 24 61 0B 0B FC
 78 1D E5 2C 32 EA 9C D0 DE F3 8C DF F7 34 A4 13
 BF 96 DC A0 44 45 80 10 26 54 5F F2 C4 BC DC 4C
 72 DD 9B D6 F5 52 3A 6C 53 BD F8 F0 BD F4 C9 B4
 A8 35 BB 69 72 CF A0 49 1C 61 4D FE 0D E4 2F E3
 E0 75 88 FD 51 1F F4 11 1A FF FA 74 A8 CC 3D 8A
 A9 26 E7 EF A7 8C EB 15 6B FA 3B 5B FB CC 6A 44
 BE 1E 76 F1 1E A2 6C 4C 43 3F 62 DA 11 9A 97 93
 E8 50 58 48 88 97 02 1A 06 CA 03 B1 88 A8 93 AD
 D3 BC 07 17 85 4C 11 1E CC 52 B2 66 E6 93 C7 FF
 9B AF D8 07 40 0A 65 FD 06 1B 8C 03 2C BD 79 22
 7C 7A CC CF 7B 17 A8 DA BC 02 0D C9 4B C3 19 9E
 F3 D0 79 06 11 75 0A A9 6A 1A A0 33 BA A7 BC 83
 2B FD AF 5C 67 D8 E1 8E FB 83 19 87 E9 D4 B9 56
 6F 84 8D 5E 60 3E 16 65 BC 18 AB F4 BB B6 5B A2
 4E B2 9D 26 9C FB BA D2 20 A5 9A 9D 75 E3 47 80
 D3 CC 36 9D 00 21 1F 03 19 DE D0 DE 92 A7 25 21
 1C 7D 35 29 92 15 CD 2D C0 50 1C 86 D3 0F AA 67
 1E 58 11 AA 83 AA BF F1 AB 9A 5D 34 4F 50 D4 15
 8D 36 2E B2 72 48 96 37 3A 1B 04 A9 68 03 46 89
 E6 D3 C3 16 29 1B 7C 8E 1A 35 C4 CC B3 7C F0 B4
 38 6A 3D 79 F4 A7 D3 EF 9B 94 DB 4D B4 1A 43 3B
 48 F5 89 FA C0 84 B6 D0 A3 3A 63 F6 D5 55 80 75
 A7 72 FE 29 12 A6 0A 16 05 CC 3F 85 9E DA 4B 85
 2F A5 52 E1 07 21 BE 46 FC 88 5D 49 05 BC EB FF
 93 60 FC EF D0 55 91 DD 92 86 59 E2 DE D2 E5 F3
 EA 33 64 37 3E 7B 30 5F 4C B8 30 60 4A 0F 36 0C
 7F 5B 0D F2 B7 DE 33 F0 98 2A 14 9F 7D ED D1 8B
 31 8A 60 C7 94 FF 8A 89 33 47 01 63 5C DB 41 47
 E6 E9 5D 95 36 04 20 89 D9 07 C0 F8 85 18 9E CD
 52 A3 04 E1 83 A1 07 5E C0 C7 EF 43 AD 0D A0 5C
 19 66 E3 CE A9 0F 4C 01 CB 45 A2 73 27 ED 7C BD
 05 DF 33 40 1E F3 0A 37 86 32 7B 36 BC B3 4D FB
 5C 53 EC BF 70 54 AD D4 63 AF F1 6E 88 A8 71 4C
 80 8A DA 11 BD AD 87 7D 80 9A EC A2 DB A7 48 34
 98 BE 82 AF 50 48 26 E3 C1 F6 89 EF D9 18 59 C7
 50 3F 3E A3 4C 54 50 81 CC CF 22 FD 28 26 38 83
 36 B0 B2 60 AF 5C 51 D4 1F 4E 8E 90 20 FC 05 72
 85 3A 22 CF FB DD D5 78 98 59 BD EB 44 31 66 78
 38 69 AE D4 22 C4 A1 51 BE F9 46 CD 19 A4 12 D5
 6D B9 C9 CE C6 71 11 C1 08 63 60 08 86 A3 1F 69
 6A 4C 3B 05 CE E6 46 77 1B 16 34 85 64 CA 0F 81
 69 D6 0E 49 06 FA 27 4D C6 55 7D FF 12 F6 4A 8B
 EF 8D 39 5A EE 45 69 B6 A6 1F B0 FC FC 37 1A 98
 91 52 DF 24 EA 02 36 33 91 6F 96 06 6D 3E 23 ED
 2B 94 D1 5B D2 C2 F2 92 6F 95 4B B2 FF BB C1 4A
 E7 AD 7A EB B3 37 F2 C5 D1 DD 54 C3 B9 67 78 C3
 FC 72 4F 79 8A C5 10 2F 9A A0 FD EE 88 47 39 79
 30 6D 00 59 04 72 F1 B9 3A C3 C0 0E 61 22 FE 28
 85 70 B6 2B D9 D1 BF 19 70 F9 96 15 DA 16 11 60
 9D 21 93 D3 95 7A AD E2 18 EA D1 9E A7 DC 24 65
 08 BA C8 34 E1 57 EB 90 69 02 41 8B C8 C2 04 0E
 36 61 C2 14 CD 1A B1 3C D3 8C 68 B3 DC C0 33 76
 30 75 E3 D9 43 CD D2 30 F7 A3 F6 EE 21 27 4E AA
 2D E0 1E B6 4C 2C CB 3B 66 F7 6C E0 D2 5E 19 90
 66 2B 91 72 F5 9D F6 9D 7D 87 F2 29 4A D8 8E F3
 86 CB 42 2A 00 BB A2 DD 2C EB E5 67 EE DC 0A 21
 AF A6 C1 6E A8 43 42 27 F8 FE 29 3E E1 86 74 3E
 B7 A2 EA F6 37 E6 71 12 71 88 04 F2 01 BD 88 82
 71 4A A7 56 3D 22 67 AC 93 8A CF 2C A7 EF 42 08
 15 0C 9B 39 12 44 E5 DF 2A 50 11 25 C1 11 5A DD
 F6 75 1C 0F A6 68 F8 BC 65 71 78 AE 94 38 78 D1
 E5 E8 BF 6D 34 8E 12 3E 82 1B 2B 15 A8 44 CA 78
 6F 04 49 A3 4D 66 BC B2 0D 7D 47 77 B7 A0 BC B0
 9C 9B 82 76 07 87 F6 34 B1 04 E6 7A 95 E2 BD 95
 7B 7C 57 C3 16 00 53 07 2C 25 79 FB 41 0F 81 F2
 B4 5D 7B 39 5D 34 97 E1 D3 19 62 8E 55 D0 AF 17
 E7 47 4D ED B2 94 2E 5B 32 5E 94 F1 E4 EC BA F7
 68 F4 A5 86 32 CF 40 F4 7A 38 9C 31 98 54 1F 6C
 3C FB 39 CE 1C D8 CD EF 38 C2 A2 6A 3F 4A C6 EE
 D5 41 4B 0E CA DC DC 88 A8 E0 4F 04 0C 39 FD E4
 94 2A 59 16 1D 5C 34 B7 71 20 80 59 94 0F BF 43
 BF C8 3C A1 2E 7D 4A 05 53 04 70 E3 8C 7B EF 7B
 1A 99 E4 89 F7 28 CE AD F4 F5 4B F4 0B 79 13 5F
 E3 1E B2 B1 51 AD B6 25 C3 31 91 48 63 65 95 CF
 45 76 50 01 4F 4F D8 8B DB 42 7E E6 6A 73 38 C8
 FA BC 2B 01 A3 1A 06 83 45 09 98 0C 9E 42 69 9A
 6A E6 1F BF 4A 40 B9 94 25 3F 1A CD 55 0B 2F 90
 FA 8F FC 0F 44 1E 46 0F 09 37 EB 21 9C 7A 45 D2
 99 76 D8 1C 2B 7C 97 5C A1 F2 EE D3 8E 40 EC 62
 44 F8 23 CF 0B 62 A0 48 DE FC CE 16 DC 3A 37 C2
 BF F7 A2 A5 FF 24 60 9E B7 ED BB DF 64 75 EB EE
 6D 51 0C 13 14 7D E3 CD EF 96 92 0A BD 09 3A 32
 55 1C 4C C1 E6 DD 01 FF 89 4E BC CD 7D FF 4A 57
 90 4A B8 AD 00 41 46 B5 7F 4C 94 36 69 54 C6 16
 3A 6B 4A 55 5A 2F B5 9A 69 3F 81 1B CA 0E 23 AE
 FA AA 97 BA E7 5A AE D3 FC F0 BB B6 B4 50 89 4E
 63 80 F8 F7 8C B3 9B 98 0F 2E 4E 4C 1A 5B 36 07
 C8 05 4F 72 3C 28 58 EC A8 82 8F D2 3B 0C 40 49
 E5 4E 9F 7B 05 91 58 B7 EC 83 29 D5 F8 E8 DA 65
 F1 CC 8A F7 37 06 14 F1 C8 AA DE EB 71 8D 63 A8
 EF 7E FE 42 4F 06 CE D2 59 FD 91 04 C9 79 55 33
 F3 A1 EC B1 A1 15 E8 45 4C 01 93 A0 B7 47 DF 1D
 F6 4C 40 ED D9 91 6A 51 AE 57 DA 56 B3 88 63 83
 B1 B9 CD 6C EC D5 D8 45 C3 4E 9B 01 3B 63 0C 91
 5D D0 DD 2B F3 54 D3 14 6A 72 AE 25 0B B2 50 87
 46 6A 81 08 1E 28 12 BA B0 F1 30 25 A7 7D 33 91
 C9 1A A6 FE 6B 17 0F CD D3 B5 ED B1 5E 44 4E 61
 2B 89 27 0B EC F7 E6 A5 B7 2E CB 50 14 92 4A 3A
 1A 7E 54 8C 32 75 0E DB DB F6 5A 39 FA 74 F2 30
 A3 A7 ED 23 1A 4C B7 F0 5A CF B6 52 CC 9C 1D EC
 4A 91 57 8A 5E 7A 6A 0C 23 07 E9 D2 AD A9 12 C3
 1D A1 D5 81 1B 0B D1 58 B7 03 C3 C7 31 62 FC 08
 E6 56 72 3B 40 36 69 53 01 C3 04 C2 37 43 6F CE
 DC EA EB 93 4A F2 7E D8 7B BE 84 6C BB 88 11 B3
 24 2D 68 D6 53 31 09 F8 26 0A 1F 83 43 65 4A 95
 1B 6E 7A 1A 40 4A 18 F0 A5 BD 22 AE F7 5B 8C 9F
 10 31 52 67 8F 06 54 E5 5C 27 43 4E 5F 68 5C 75
 D1 0E 52 05 FF 9F E9 B7 11 4D 2D 83 A8 50 9E F9
 19 F2 CF 53 D3 BE 6F 74 BC 17 5B A9 E9 E3 BB 2D
 1B 29 B3 11 B7 70 61 F0 B6 F8 3D E9 19 80 1E B4
 B4 3D BE B9 D1 3B 8B A2 DB D5 EC AF CD E4 10 BE
 30 79 52 99 F8 C0 07 FE A1 4B 4B 6D 41 DF 5B F6
 E9 E4 64 53 BD B1 7A 13 0C 7A E0 95 AC 0C 03 9F
 EA 80 05 66 2F 8B F0 06 48 E5 50 19 B1 27 64 82
 48 D8 B1 AC E7 49 B6 BE EF 89 09 23 7A C4 AA 38
 39 75 0A 7A 64 B8 39 26 8E 2B 17 8F BE C7 D4 09
 43 0C D6 F2 DD 3A 1D 51 EA 57 D5 39 AF CC 0C 1D
 F7 E7 AF 82 0C FB 29 2B 72 8D D8 19 B5 B9 95 FE
 E5 2B A4 6B C4 4A 62 C4 96 57 82 FE 5F F9 B3 73
 BB 35 9E 6E 25 61 4E F8 AF A3 4F 96 45 8E 41 21
 A3 F7 47 C3 AB 0D E9 FA C6 00 13 3B 9D 0A 1D 4E
 EF 83 75 B0 41 34 FD 3D 56 E2 1A 9B 63 BA 6A 8B
 84 A7 97 22 58 69 33 64 5A 89 73 31 FB D4 8B 89
 9F 89 2C BB C3 92 CD AF 4D 44 4E 07 66 21 A5 32
 10 60 01 F4 EA 13 4D 9E 77 44 08 6C 88 17 EE B5
 3C 13 45 C2 C5 88 F9 E5 AF A6 EC 1B 57 A1 63 5D
 52 5A 11 6C 7C B4 5E CF 21 38 F7 7C CA 76 B9 FB
 6D 6F BD 6D 73 C9 7B 7B CF 40 AC 57 E0 DC 38 47
 15 A9 0F BD 50 BD 6B 6E A6 61 9E 79 B6 AE BD 84
 57 E4 8D 42 B8 CF 4D BF 80 B4 3C 9F CA 99 0A B4
 FD C3 C2 35 82 BF EC F5 29 83 22 37 AF D4 75 CA
 C6 D9 6B AE A9 C2 81 14 A0 8A 68 68 68 1C F7 D3
 1E 5F 25 08 20 99 4D 65 55 7F CB 6B AE 5B CC 0E
 48 4A 19 D1 35 44 62 F3 DE A8 12 6A 24 EC E0 0A
 A0 A9 A5 08 15 04 79 4F 20 DF EE 38 69 D8 EA 9F
 70 E2 60 2B 2E D0 32 3B 17 4D E5 51 16 68 F1 A2
 94 DC E1 9A 08 D5 B3 22 0D E3 BE 2F 1A 4A 62 64
 6F 10 08 FA 46 AC 0A 90 27 7A 6E 57 DB 14 95 A9
 63 F3 C4 44 8A 03 5F 27 82 33 F1 2C F7 34 4F 2E
 06 F2 3D 6E B0 E1 40 5D 0F 94 8C 88 88 35 36 03
 A7 8F 97 0E F5 6A 46 DE 5B EC 31 A1 26 E8 10 80
 8D 3A FA D0 3E 4C F3 95 3B C1 63 12 C6 67 5F 1F
 EB 18 C6 B5 8C E2 C4 B5 42 06 8A 21 CC B2 A9 75
 54 85 11 C1 AD B5 1F 12 18 4E 5B AA 47 85 BE CD
 C0 E4 01 15 8C BD 4F CE FA 35 C7 A8 00 27 43 65
 38 F3 6F 47 A9 B1 EC BA 79 A9 D0 EC 1D A1 E0 CA
 09 E5 5D CA 84 C4 34 3E 38 F5 2E A0 2C E3 AA BB
 7B 97 B3 0C BB 2B 6F 6D 06 DA B7 BC BF 08 43 31
 01 67 A6 25 88 49 03 C6 CC A3 DD 32 AD 9E F5 83
 6E 41 FD F4 F4 A2 FE E7 8E 4C 93 D1 19 2E CA E1
 53 9B DB ED A4 CA AB C9 35 F1 FC ED 54 27 AE BB
 56 EC 3A FC 7F 27 ED 8A D3 6A 7F 98 B7 A6 33 A8
 E7 BD E4 6B 77 87 BD E2 25 66 16 3B 14 51 25 53
 0C B2 42 C8 D1 7F 9D DF 25 97 1E 5D 4B 18 15 E0
 DE DC EA 84 0F 89 D5 42 28 C9 7F 31 F5 D4 DA 14
 4A 5E 16 31 50 27 5E 15 BB E9 54 C8 EB 50 DD 6F
 AB C9 49 7E 73 AF 11 D9 F4 EE E3 ED 88 EE C9 FB
 76 8F 2B F3 21 E9 D0 4A 50 F3 DD 30 AE 08 01 D1
 F0 E2 75 E1 6E 38 CA 78 58 48 A6 B4 AF C5 21 DE
 D2 BC 53 2D 18 8E C0 09 F4 20 B5 AC A1 F5 7F 32
 CA 83 11 9F 81 70 18 CD AB 40 29 3F 92 BC 94 31
 29 ED 28 49 93 7C 49 E0 9F 48 D9 DF 30 36 E9 16
 AE 4A EF F8 1B A6 84 98 9C AD D0 74 54 5C 69 6A
 8E FC A9 F9 3E AD 80 DB DD 72 0F 25 A7 58 C5 56
 AB A2 9E 11 E9 49 FF A6 A4 A3 1B 48 97 CB 41 26
 72 3B 70 54 BA EB 1F 0B E5 21 AC 4B C6 01 CD 15
 F9 9C 96 1F E3 5D 15 AB 93 29 89 06 CE BA 39 72
 D4 1C A8 80 DC 6A 97 F6 56 31 96 27 D0 AA 31 EA
 D2 95 25 48 29 BC 6A 88 85 29 40 2C 14 6C D7 F7
 3D 5C D3 48 E8 47 74 B4 B3 55 90 C3 D4 6C D9 E7
 E1 29 9D CD 8A 4D CF 9E 99 75 3C 00 A1 6D 12 0F
 B5 5D F4 73 94 71 6A BE BE F5 A9 37 BC 1A 1C D5
 51 5C B7 12 48 AE 17 98 83 A0 62 6E EB BF C2 CF
 C1 B6 6A 73 19 AE 8E 19 F1 66 DC E1 89 E1 4C DC
 40 31 46 88 63 EF F0 B9 66 DD CF 04 42 14 36 18
 C7 B5 5C 44 6A CF 07 19 D6 3B 63 1D 4D DC 44 0E
 F9 3E 9A BD 60 E5 AC 0F 83 3E 7D 21 01 6E DB 57
 4C 90 0D 6C 78 FA 35 F6 82 09 68 EE 73 DB 86 FB
 43 34 F8 FF DD 49 45 61 56 91 EF 53 A4 6B C1 20
 27 36 67 50 0F 41 1C B9 A3 9B 3F 50 F8 74 3E AE
 78 7C D5 37 45 45 73 1E B2 F4 ED 13 E2 47 86 87
 CA CF 93 3E D3 08 EF 62 23 EB 00 56 0D 1B 52 AF
 3F 36 C2 2B 78 DE 13 C9 92 90 6C 64 FC A7 50 2B
 18 79 E2 80 2E 97 EB E7 05 43 58 9F 55 6F 98 FB
 86 9F 84 04 D9 EB C1 0B 89 F3 00 20 D4 C9 8C AB
 87 21 CC 04 8A 06 BE 8C 5B 50 F8 B2 B9 BD F4 DA
 71 54 3E 1B 83 37 61 A1 E4 F7 65 E1 77 6C 7B 88
 2A 97 49 3E 73 FD 61 60 BC 0C 8B 0C 5A B8 C0 D7
 70 A8 E1 D0 EC A7 5D 7A 89 0E 51 AB 24 E8 6C E2
 73 F8 FA 65 19 EC 14 16 CE 0F 5D B7 53 D1 60 F6
 E7 96 43 5F 99 18 BD 5E 45 D2 9A 4E 3F DC 77 B8
 D5 49 E2 9A 71 0C 89 0A 31 24 2A 6A F3 5A B3 4A
 C9 B9 30 97 B5 62 42 F4 3F 97 C7 73 EB FA DE C5
 13 AD 02 2B D3 8A 0C 2A B5 74 82 C2 9B 05 C2 5E
 11 3C A4 59 39 44 7C 19 AB 18 74 CB EE 38 DD F0
 B6 D2 5B C3 CF 78 9A 0F BB AD B3 68 AF FA 9E CD
 1D 99 6A FD 42 8A 9F CB 70 E4 E9 0F DA 97 7C F9
 76 EE A4 B8 38 EC E4 98 45 45 FE 2C C4 1E AA 50
 9F 8C F2 04 B8 AD 5A BD 23 2F 42 A2 89 6C AC 30
 F4 4B 9D 25 32 27 F1 29 72 C9 ED 46 3F 13 22 16
 53 BA D4 EC FD A7 3A A5 73 FA 99 FF A2 5B D5 99
 B2 78 99 B6 92 47 7A 28 9E 07 E4 4B DA 0A A1 55
 82 CE 36 A1 E5 81 11 B2 A1 4E E4 EB 27 92 BA A1
 08 21 C9 56 86 00 20 54 AD 21 09 39 C2 0F 04 F4
 F5 15 99 A7 9C E4 F7 05 BB B0 CA 05 27 75 0A 59
 20 35 A1 18 11 20 A3 3C D0 C3 CC C8 15 12 C3 A1
 92 F5 DB D1 D3 CF 08 96 4C 2B 95 66 A2 C5 2A 1E
 FA 03 B5 A7 A8 6E 35 64 76 85 E7 6E BA 9B 68 AB
 E2 7D 60 4F 36 FF A3 4F F9 35 40 0E 0A 4A 81 F5
 DA 1E 6F 8C 59 8E CC 13 D8 78 6E 28 31 3E D5 35
 87 05 DB 3E 95 D7 F9 FB F3 3D 2E ED 05 17 61 1B
 6B B2 47 1C 45 FB C4 58 ED 1E BF FB D3 42 7A 5F
 5A 6F 21 6C A3 6B 03 FF 80 29 05 2F CC BD C4 0D
 D1 63 7C DD AE F4 50 B0 B6 CD ED D7 EA FA 99 70
 0E 9C 53 5A 20 6F B7 33 24 58 3A 5E 27 84 CC AC
 C9 B0 A8 4C D8 04 48 B6 09 17 2F 53 13 E2 3F 0E
 85 2D 02 97 62 B2 1D 30 14 E6 18 5F 1F 38 D7 59
 2C 00 42 45 D1 69 32 AA 24 E3 FB 56 FD 5C CE CA
 03 0D 76 1E 98 11 50 CE 4D CB 04 53 38 A3 85 36
 50 24 2A C7 0D 05 79 F0 E5 A7 0B 5C 03 F2 14 97
 D3 3E BB 56 26 2C 26 BD AD 28 1A 49 DF 12 1B 6B
 14 B8 CA 33 CB A0 B9 10 71 44 69 7E 7C D6 FF EF
 A5 7A 58 3A 65 09 8D 13 88 A0 9C BE 51 3C 55 97
 1E E2 24 AE 1E E4 B9 6F 88 57 A4 54 2D 65 75 2A
 45 05 22 24 AF 34 3C 51 0A 7A 27 9F 3E 7C 60 76
 C9 DE D2 E1 D1 1C EA 46 B6 D0 BA CC BA FF 33 71
 B9 0D 8B 7D 13 14 5B 39 70 21 FA 77 13 F9 52 2C
 89 DE CA 7B 59 EA 91 78 C8 2D B5 7E 96 A4 60 92
 E6 E8 A7 7E 2B 7C 16 8E B0 DF D5 93 82 78 76 AE
 B4 D3 FA 4C 70 3E D0 20 B2 29 A4 A0 CE 0B 7F 6E
 13 05 82 F0 DA 9F 12 C4 DC E4 0E 3E AC 5F 18 62
 F9 6E 5B 6F D6 90 A2 C0 38 3B 95 0F F7 B9 5D CC
 FE 16 D7 6C 24 39 F5 50 1A 77 95 75 63 8B 4C E7
 2C B1 E5 3B 6B 45 F0 CA 8F 63 75 11 C9 30 6A 1E
 44 3F 73 DF DF 30 67 96 5E F5 D4 5E 00 C4 1A 96
 C7 C0 F0 4C 2B 00 19 41 91 E7 BB 25 AD E2 51 8E
 0E 39 F3 37 3E E1 F5 2C 13 A8 A7 A4 F4 58 2B D8
 4C F0 48 E3 3F 30 0C 2D AD 60 BD 0C 3F 3D 74 94
 D0 EF B1 50 5C AE 49 EA C0 AE DF 26 0F AF DC C4
 C6 9D 08 E1 0A BE 39 82 FF 66 A9 9C CD 6B B6 6C
 76 DE 1E CD 59 11 04 29 8A A6 37 A9 1F 91 17 08
 1C 6D 47 0A A5 68 3A AD 63 05 A3 B1 AA F5 82 93
 2F 9F 8C CA DE B2 B9 33 78 0D D9 0D 43 82 98 CE
 01 38 21 61 E6 3B AD 61 3A F7 29 3B 2F BC F6 23
 D4 C8 A2 83 E0 06 63 DD CD 65 30 07 7C 28 94 29
 49 15 1B DC A7 81 7D 7E AB B6 77 70 D9 CD A3 06
 BD 8D 79 49 02 19 E8 BF D1 15 0B 23 E3 61 87 CA
 8B 54 F4 67 51 6B FE 0A 97 41 36 80 36 E0 0D 62
 82 88 03 6B 68 56 FA 0C EC AF 27 10 96 66 6A 81
 33 A8 FE 10 D7 01 72 C3 15 1B 3C B1 C2 C3 13 B5
 E3 8F C0 47 99 42 E2 4E 54 05 9E EC B1 DE 77 A7
 BC 52 40 E2 1A A3 7D 7B 82 B6 69 19 D1 8E 8B 30
 35 9D 11 2C 30 86 B2 1A 14 65 12 09 68 16 13 55
 71 F5 99 1F D5 95 5A 66 48 6B 27 56 F9 96 E1 B2
 DF 5E 33 F5 CF 4B 03 2E 2B 80 15 C4 30 48 2D C7
 B5 08 EE 48 46 05 B4 28 5E 5D B1 E0 F1 7B 8B C5
 E5 69 10 51 1D 81 33 AE D7 1B 12 B7 00 5F 41 7A
 77 53 00 E2 F7 EE 79 AA 86 2F 0B A4 3B AD 7D 24
 53 A8 67 A3 E3 1C 57 02 A2 2E BA EC 82 7F 04 D4
 53 D0 6C 72 33 94 F1 68 2C 70 77 2D 15 19 D7 23
 27 D2 38 FF C8 08 B9 3D 2F 46 6B 46 59 1E 0B A6
 A5 73 0A A0 9B EA 93 32 A3 A3 B3 62 E0 32 37 DB
 69 29 31 1B BB 93 68 1D DE 49 B4 8B 4F 34 CA 3B
 B6 24 42 6B 3B 2A 64 DA B3 53 FA 8D 66 C3 69 5B
 46 FD AB 0D DB 3C 1E 1F B8 01 D2 0A D5 46 37 EC
 84 D8 75 48 B8 21 9C 38 41 5A DC 50 E8 C3 82 21
 AC EE 34 CE 96 7E EA 33 1F 00 B9 85 CD B4 7E 9B
 9D 38 D3 F8 65 D4 1B 4B 80 68 A0 E2 42 E1 38 58
 7F 34 5F 85 3D 58 A1 67 75 43 BC 43 F8 FD 69 F7
 63 70 90 27 AD E2 8F BF 9B 22 1E 49 CB 11 69 53
 B4 D2 6D EA B5 15 00 F2 F9 9E 98 DB 84 7B 0E 3F
 54 53 05 A6 10 0B 97 5E 36 74 70 26 71 A2 30 F6
 26 04 B3 F4 4A 1F 19 4B C8 F9 A5 35 14 7D 45 56
 B1 37 39 E5 37 AA DB 79 F2 91 1B D2 8D AB 0C 54
 96 4A 7D 57 2B F6 05 4F 41 A1 02 1D 51 F5 2F A6
 57 40 0A D6 9A F7 9D 22 5C F8 3C 68 73 C3 29 C6
 7B AB 55 8C A6 01 7A 87 6A 18 49 FF F2 5B E1 3F
 0B B3 80 81 40 8A 42 11 36 14 97 78 AA C3 F5 1A
 1B 45 4B 7E 8D FE FB A6 F2 D9 9D 6C 15 00 93 F0
 55 B2 4B 31 CB 37 79 DC 46 A7 5F 33 65 95 5D 76
 5E 7C 65 C1 47 A2 CC 0F 0D A5 75 59 BE EC 27 4D
 D7 F8 D1 B5 DD E8 E3 67 C2 FA DB B4 A4 58 FA 72
 26 31 90 D2 C9 D2 AD C9 07 93 F1 9C C3 A1 18 CC
 89 4F 12 2F DE 52 3C 47 5F 9D A7 28 8A D8 80 95
 0E BB 9B DA EE D5 3C 52 7D A0 A1 44 CD 9D C2 30
 07 99 DD 86 E2 B7 32 DB 1F 74 CD BE AF 1D 33 9C
 E0 05 8D D7 55 35 02 44 FB E5 67 BC 20 14 E4 C9
 F4 1F 80 0C FA 70 AE AF 17 08 BF 1A 8A 42 30 0A
 E3 43 DB A9 AB 34 B1 89 10 A6 12 7A 8A 4A 56 77
 C4 15 E2 5C 6C 2F B7 EC 7E 42 DF 45 90 E9 AA 6A
 37 D2 56 7D 3B F7 70 0A 05 EE 17 0D 2F B8 FE D3
 16 AF 89 24 94 6E F5 D3 E4 BF 75 A6 76 4B FE 3E
 19 E3 85 4B E1 3E 5A DD 78 6D E6 F0 5D 1E 9D DC
 A9 5F CB FE 35 33 D1 51 84 8C B6 BB 95 5C E5 C7
 F3 BA A9 5E 67 DA 75 DB 7B D0 4E E9 FA 6E F8 CE
 92 1A FB 34 63 58 9A F7 2C 2B 28 20 11 0F 03 BA
 61 AF F7 5F 4D 60 6A B2 97 4D 23 02 63 4F 81 88
 5D 95 42 9D 5F 1F 9F 2C 89 2C 65 B0 75 8A EF 95
 EC 36 6A DB 6A E6 BE 83 2D 3D 99 8D 74 2A F3 DB
 D5 94 09 ED 87 D2 ED 25 5F EA 4E 7C E2 DF D1 CE
 7A 9D F5 8E 50 59 03 3A A6 A2 CD 1B 71 BA B4 71
 CE E0 3E 7B D5 6F E9 2F A8 DD C3 1D F2 7D DC DC
 3A FF C6 05 F0 A7 C3 D7 2A BA 87 84 B5 E8 12 D8
 D6 61 3E C7 D6 1A CD 0B 96 0A 0F 39 56 D3 86 1B
 09 D0 6A 50 CE 81 E5 41 24 59 C2 AB CC B8 C0 38
 F4 D0 39 AB A8 63 87 31 C9 FA F1 6A 73 0A 4A 88
 BE 3F 3C D6 79 78 C7 D1 AC 3E 88 82 D5 E1 6C 37
 61 6F 37 AE D8 A9 2E 39 1A 1C 7C 38 BF C0 CA 80
 E1 7B FA 56 97 F6 6B 04 2B 41 8B FF DE BE 16 74
 B4 91 8B 33 63 12 F5 20 1C D9 EE F8 E4 4F 7F AA
 5C 66 4B 4F 8B E2 AB 1D 6B D5 19 53 7D FD 17 C5
 42 7B 3D 81 02 29 86 09 F4 7B 22 63 CB 75 12 4F
 10 50 8F 77 D2 AC C7 0C 29 01 6F 56 11 11 9B 10
 5F F4 9F 0B 65 30 85 42 81 5A F9 B9 EC 26 CF 18
 EB B8 FA 3C 26 3B 65 02 36 75 9D 42 CC 6C BA 5E
 A3 5A 0A 7E 63 C6 47 04 0D 43 ED 46 5E BB AA FD
 DE 6B 43 38 C1 80 06 52 44 A5 7F 36 87 8B 2C A7
 79 FB 1A F0 68 AC D0 2F A0 84 9F 33 77 F3 FB 6A
 20 36 95 09 60 E8 B4 14 24 F6 80 EF 08 11 0E 97
 D6 EE F1 2F C4 2B 0A 07 EF 6F 75 4C 84 D4 4D 18
 3E 2E C3 CE 2E 7E F6 9D 43 08 B9 AE 11 C7 22 71
 36 CD 8F 01 96 33 D1 16 8A 68 39 1C 3A CF E1 C3
 9D F3 94 8B D1 F4 BF D9 F5 68 E6 BA 4D E0 95 CF
 9D 6E 81 CB 44 8E 72 F1 B1 1A F2 E6 11 D5 21 AD
 BD 8A DE 47 EC 3B 23 1D EF A2 BE C4 5F BC 6E 91
 02 25 8F 56 F0 2E F8 81 22 F4 3B 86 05 B7 FD 04
 1A 38 30 81 CF EA D4 03 55 05 26 75 EA A0 8B 2E
 AC 0F 20 73 2D 44 F7 5C 46 AF 38 71 5D B7 77 06
 A8 11 DC 4A F7 70 C5 50 19 6F C5 F1 E4 E3 6D F8
 27 D5 C9 AC 4B 0C 64 8E 75 88 A2 C0 B9 E0 10 70
 56 3D 88 E8 E3 C0 A0 78 BB 04 1D 75 F4 CF A4 CB
 E6 00 95 9A 93 CF 43 E7 87 55 71 82 BE 49 80 F6
 B3 D1 DC 3E 20 9E 32 2B 7C A3 F3 06 EE 52 36 F4
 C3 AC 90 D8 4A 2C 35 08 0B 30 DF 00 6E D5 6D DB
 EC DC 82 24 D1 44 DD 67 77 04 A5 73 00 AB 60 A8
 E0 34 0A 2C 10 43 F6 91 14 BA C2 51 6C 3F C8 B8
 D4 28 8E 34 11 85 B3 6B 47 FF D5 84 15 25 92 26
 69 57 A0 A7 78 D5 E1 4F F0 3B 6D 7E 4D 4E B0 AC
 AB 00 21 8E DB AE 9C 37 42 86 03 68 E9 FC 1C B9
 80 27 51 1C E4 C5 FC 64 0B 61 31 E1 4B 49 A2 E1
 3F 04 38 50 DA EA 35 65 69 EB 99 B7 1D B2 C3 D6
 9F 57 C0 80 D0 7F B8 0B 5D 19 E7 0A 96 81 A9 22
 19 EC B4 DB 5C 7B 33 86 A9 2E F4 9D 18 49 29 64
 74 B8 42 02 FE 5E DA AB DC 6A AA B0 5B 55 B8 FB
 B0 D9 C8 7C 6A C4 C0 AB 6F 5C 8E CB 38 91 13 BD
 AF 61 A6 D4 6D 2D 01 7F 9D D4 86 5B C9 7F 9E 82
 E3 62 32 3A 8D E9 BB 80 4A 28 24 C1 83 26 21 8B
 9F 70 D1 98 F5 9D 86 7A A6 C5 8B 75 8D 97 E2 5A
 6A 28 71 B2 94 E6 3B F2 0C B7 54 4C 38 55 5D F5
 18 1B 09 47 54 EE 07 80 E9 9D 34 ED 0D D7 4E B5
 93 06 FD 1C 88 EE 9E 21 06 B1 8A F7 66 FE 14 FA
 22 71 2E 30 F2 14 48 3A 2F 97 3E F7 9E 7E 2B F2
 18 FA 23 50 0E A1 EA 50 73 4C 0F D1 EA 7E 8F A1
 8F 16 8A 9A B6 3C 9C 74 90 F4 23 9D 56 1C CD 9B
 6F AD E1 58 81 28 0F 77 C9 D3 D3 CE 6B 7A 29 BC
 E1 1A 50 6F 92 49 57 7E D9 D2 23 67 C2 37 72 55
 9C DD 7A 04 DC D3 B2 18 A1 24 4D 43 E2 3F B1 67
 BF 28 B8 F8 A4 B2 8A 88 87 41 52 DD 20 32 9D 4F
 67 13 3A A1 BB C8 82 19 02 29 73 93 AB 09 8D C7
 E5 30 7D 72 92 37 36 11 AD 66 53 99 4B B8 64 C6
 55 05 C7 74 E7 4C D5 18 AE DE A3 21 F5 EE 1A 80
 15 19 00 9E 3F B3 BD 3E 09 15 18 9B 2F E0 26 23
 E7 33 1C 19 B5 A5 33 9F 82 B7 7A 26 4D 54 FE E9
 38 35 5C 1C 80 F0 D7 E6 C9 1E D8 58 5F 31 97 B4
 3C E6 C3 D5 CF 78 0A 0A 6F 5C 6C 77 A9 0D D6 48
 A8 A3 F4 C2 61 32 05 9A F6 12 14 B0 14 A9 5F 93
 0B 39 E1 EB 33 26 17 F9 0A 9E 85 00 27 13 E3 DB
 D1 90 A3 4F 06 D8 53 D4 21 35 1F C9 42 1C 16 2B
 32 6F 43 28 02 BF DE 73 B6 55 1F 1A 30 AD E0 2F
 0A FC 69 B9 F6 82 F5 58 D4 6D 21 39 E5 4D 75 EE
 7F 03 F1 33 3C 71 8A DA 5C E8 3A 22 EB 2C D8 A5
 58 DD BB BC C1 55 45 E1 6B D1 FD F4 E9 77 80 83
 B0 13 8F BB 75 0B 06 B6 98 7D BD 82 F5 1E A0 5A
 FC 11 FB A4 8B CC 54 BD BF 86 5B F1 FB DB F4 F3
 78 92 61 FA FC A6 36 45 A9 6B 45 EC 93 FC 8A C7
 FC BF 4E 56 8B D2 93 96 7B 7C 03 83 84 BB 21 14
 A2 2C 1D F2 F1 DA 26 6F 4F 94 7C AD BA 99 E0 EF
 E6 04 D5 03 E6 92 D8 4C 62 EB 73 DC 65 8A 83 53
 CC 03 AE 05 E3 ED 28 42 EC 8E 1B 3B A8 B8 6B 92
 FC 7B 62 CE 78 6C B9 EE 80 9D DF 69 09 46 06 35
 44 3F A9 FC 8B D0 37 02 26 74 27 BB 39 D0 A6 1D
 34 ED 93 84 26 90 02 27 E1 A1 35 ED 12 0A D7 66
 7F 44 6F 12 FD 02 C9 F4 83 06 3F 05 3A 5F 8D 6F
 6B F6 E7 C6 E8 E7 3A 70 58 6A 01 E1 98 4B B3 72
 E8 1C CC 8C 20 03 E5 98 56 6D 66 FF 04 B5 4D 74
 D6 65 3D 15 70 C2 CA 12 E4 85 CC 33 80 3C 78 68
 F0 D5 82 82 FA 7D A7 4C 87 E8 B8 05 76 BE E5 82
 A8 93 9D 01 4D 1B 8C 59 E6 AB 1F 68 19 D5 5D 75
 7E 6D B3 47 79 E1 DD 54 AC A2 89 27 D1 C5 5B C4
 95 D2 64 C5 F2 B9 A0 C9 5D F1 A5 8C 5B C6 39 5B
 D9 C5 D1 C3 5E DF 8F 3A 22 4A 5F 74 3B 5D 20 B5
 1B 41 03 FB 4C 1F C9 12 A9 ED 62 10 5C AB 7F D6
 6D 6D 73 B2 48 41 56 6B EA B1 3E 69 1D 6C 2A 68
 66 6C 91 84 BE C2 85 57 FD 48 2B 27 8E D9 DD 08
 1B 3F E4 9D 47 4F C0 03 34 0B EA 60 98 42 CE 35
 2E 56 3C FC 3F 63 57 92 17 3B FA AC 40 C9 99 D3
 AE 30 12 50 A7 77 98 57 1F 89 AC F3 1C 4C 19 5C
 BF 64 54 7F FD 6D F6 FA C5 81 1F FD 10 BF 73 2E
 D0 E3 01 9E 0B D6 31 74 89 52 19 6D 61 7B A3 48
 F5 A0 B5 3D B8 7D A2 9D 33 12 6D 32 97 89 D2 5C
 DE BC C6 F8 2C 83 7B 30 38 91 70 28 5A 96 71 90
 7C 1E 83 BA E6 A1 80 C3 C6 F4 40 D8 F7 9A 44 9F
 17 54 6B 03 F6 4D FF B2 CA 67 58 4F A5 A2 6B AE
 2C D6 4C 7F E1 BD 42 46 7E 30 CC 80 36 B0 D1 47
 DC 12 E3 E3 9C 3A 44 93 C3 9D EC 96 AF D1 EA D1
 D2 31 FF A0 42 E3 D5 30 D2 8C C4 EB F6 43 1A ED
 B9 2E D2 C8 3F 19 0E 54 A8 DD BB DD B1 6D 0C AF
 0A EC 4F 6D BD 13 35 71 4D 27 38 77 2A 3E 64 7F
 80 4A 84 74 9C 74 2B 88 E2 15 3D 14 34 63 2B 11
 6E 82 43 87 8A D3 39 7D E1 6F EA 0C 28 9D B2 23
 59 69 6C 87 10 9E 85 0A 27 84 40 49 5F 63 B3 E7
 60 4E 79 C3 5D AB 82 19 4F C1 16 EF 7C 80 D0 C9
 EC F7 22 B0 EC 15 64 64 2D 42 AF 98 5C 4F A8 5F
 C9 A8 86 7A F4 99 B2 15 FC 33 51 CF F6 51 E4 EA
 3F 58 2C DD 7A E1 AC 24 F6 52 75 B5 99 36 71 63
 87 2C 11 D0 89 CC D5 62 F3 AB C4 92 DE E9 3D 72
 29 D8 DB 7F 28 16 32 31 BE 0B 46 87 04 3E 78 7E
 33 C1 DC E2 8F 7C C5 CA C8 36 CB 55 D9 0C 7D 83
 06 36 4F 71 65 27 DC 1D 9E 1B B3 F9 D3 E4 04 23
 CA EA 10 37 28 12 2C CB B7 E5 76 A8 EE 99 9B 9A
 05 56 88 93 D8 1A D3 EF 05 91 28 BA 2B 2B DC 7B
 C2 A0 27 4B 67 D1 07 E9 FD DA 78 4A C4 D8 BA E1
 4B 03 ED F2 D7 F8 6A D0 F1 85 72 91 CB FB E0 04
 FD 0D 1A B4 00 A5 E0 87 AA 79 DA 26 55 E3 26 23
 42 FA 0C 88 71 15 E6 8A FF 51 5D 64 0A 4B 23 FA
 F8 2C C9 BF 9B B2 CD 0B 6F BA A2 6A 7D 75 A8 EE
 19 AB 72 D4 AF 5F E2 1F 50 8A BA 8B D5 EB 87 2C
 5D D8 39 A3 48 8E 40 83 A4 8B 5E 17 F6 B5 DB 65
 87 B7 6D 7F F6 AA 7A 67 6B 19 AC EC D7 F9 B5 89
 A6 B5 AD B6 21 E7 73 DE 6F 97 06 84 21 9D 74 5D
 97 F5 EA 92 24 6C AB 8A 3B D9 84 24 A8 15 82 E0
 38 66 4D BF 18 C9 1A F6 A3 06 9A E2 C6 2B 26 E5
 A2 9A 45 FB 0B 54 38 90 41 C0 16 F0 40 06 CC 4C
 60 EB 6F 44 4B F8 B9 92 EE 19 4F 07 E4 7C EB 72
 42 E2 0B 04 BA 44 0B 1E 41 60 BA 13 13 33 E2 D1
 51 E2 BF 4F 47 79 2D CD 57 CF 98 E6 4B 82 D8 82
 60 5C 58 B4 84 55 F6 09 12 9B BD FE 31 F7 89 36
 E2 04 E8 C7 62 A9 0C D1 35 B7 23 B9 41 8B AC B9
 72 90 E1 A9 27 94 9A 81 56 45 FC 79 E1 FF 72 AE
 0A 76 48 B4 D2 4F 9B 90 20 6B 97 4E 40 E2 41 D6
 63 BF 0B 0C AC 5E 58 DD 8D 71 43 4F 01 E1 E6 9A
 95 CB 2B 09 43 56 E2 D2 59 15 F9 35 3A D2 A7 2B
 02 BE 3E 1A 33 36 10 6B 94 B8 71 14 7B AB B7 6F
 20 73 3B E1 76 B4 55 DA 47 0D 88 BE 1E B6 79 F5
 B1 AE 33 EF 3B 3A 2F 8D 9B E4 AA FB 03 9F 2E AF
 46 C9 5D ED C1 BE 07 37 04 98 D6 69 5B F1 13 E5
 93 F5 81 BF D5 B9 79 18 49 12 4F 33 D9 06 11 CC
 4F F9 53 7C AD AD 27 A3 53 C0 29 22 B5 22 0E 1E
 B7 34 62 2A F1 99 1A 4B 96 25 17 91 31 CB E3 E0
 B7 95 4E F5 B5 EB 79 96 22 2D 97 22 FB 29 FE 71
 AB 7A 44 78 B6 1C 9B AE 49 08 EB 35 85 CD 8B 8E
 76 D4 14 82 4E 08 AC 1B FA 61 F7 73 28 D1 B0 A9
 BA B6 47 7F 62 19 F2 2B 5C A2 8E CB BC 07 5F 5E
 73 92 7C 48 AC 7A 85 A6 22 F0 4A 77 06 43 8D 4C
 8F EF 0A 06 39 07 BA 44 C2 DE 2F C1 77 AC 8F 6C
 DD B4 A7 FA D1 D8 D0 7D A4 7E 27 20 78 F8 F8 59
 D8 14 A2 FE A4 E0 3D C7 0F F0 DA 0F AB DC 5A 8B
 F4 BC 08 BC 12 C6 70 52 E8 0F 64 81 F3 EB 42 E8
 90 54 93 CD 03 63 D7 97 70 E6 DB 6F 27 3D 3D 3A
 ED 64 20 2F FA 35 18 16 00 CD B8 27 3D C4 1D 36
 07 35 EC 75 A1 B4 1D 25 6D 0C 98 28 D1 4D FC F7
 BC BE 51 AC F4 D7 06 90 E5 AF 33 C6 E9 50 FB 2F
 8C B0 5F A9 0F 5C E1 DC 26 E6 F8 37 E3 2D B9 10
 04 FF 89 78 C1 1D 9F 4E 12 AF E0 84 93 94 57 96
 70 0C 0D 0C A8 CA B0 2D CA EB 2F 6B 0C AA 60 BB
 FA 24 4C DF 74 A5 74 9D D7 7A C1 11 AF 70 6C E4
 12 D3 74 43 8B 9F 28 90 D9 B8 97 8A 7B C4 D2 33
 EE AD E5 AB 52 A8 F6 D9 E4 5A 98 17 C8 2F 4E DF
 90 07 A3 7E 36 1F 17 9A 53 DB 81 7B D8 4E 65 CE
 7F E9 23 A3 CC F7 1A FF 6D E0 14 0E 34 DA BA 91
 F3 BE 89 03 B8 E3 A0 35 A5 19 EB B4 82 B6 2E 65
 D9 16 55 79 33 5F FF BB AF C3 42 85 1A 86 34 C7
 3B 41 74 03 10 38 62 73 9F F1 8C 86 07 66 C2 2C
 94 FF 55 16 5E 87 87 02 C9 B9 73 5F E8 B4 DE 28
 B9 E5 14 F9 C3 DD B6 9B 66 5E 30 70 C4 8F 55 AE
 94 4D D2 B9 1B 1F DA C0 AA 28 5D B7 A8 D8 AA 4F
 85 6B D5 B4 D2 EF 2F D8 45 2E 7B ED A5 B2 E5 1F
 FF 37 A5 81 4B 94 C0 36 56 B2 3C A8 21 56 23 0C
 82 F5 89 45 1A C2 6A 9C A2 69 61 CA A5 50 DF 23
 7A 6A FB 13 C0 38 36 7C 1D 72 EE CD 16 08 FC 90
 B0 DE 34 4E 0A 6E F2 4D 32 0C A6 AC D1 7B EA 11
 06 9B B1 83 89 F6 77 11 E2 01 6E FA 42 5E 42 55
 19 5C E6 BF 2A F4 64 7C D2 8A 6F 84 11 84 2F 13
 DA 71 E2 C7 80 9F AA 68 8D C5 AA 5B 57 A7 4D 1D
 47 71 5C B8 51 CB 0E D7 AA B4 DE 33 7E 05 BA 67
 06 02 6B 2A 6C 22 11 E3 BF 68 3B 0F 7A B7 2F FE
 18 CF 67 01 E9 2D 66 40 B0 66 C1 41 41 7A 02 0F
 98 06 F2 53 A1 B4 4C B2 F3 67 BC 56 2F CE 42 83
 78 D0 84 86 3D 25 0E 2C A6 BF 27 F1 58 F8 EC CB
 6F E2 D7 8E 46 CF C0 7C C2 BE F5 72 CC FE 61 13
 D0 96 70 85 7E 98 31 6F 0A 31 05 49 6D 88 5C DE
 B4 A6 E3 35 73 E4 4F 04 46 D5 5C D5 B7 E0 3C F3
 DC 30 55 CD E9 6D 2A BA A8 75 33 86 7C A9 97 C8
 7A 47 07 EC DD 6F 26 A6 53 99 DB 48 63 7C 60 9A
 5E 84 AD C1 BF 3B 1E FC CC F3 80 C7 18 E0 DC 39
 66 F2 A6 AD 6F F5 9D D3 97 DF A8 94 00 C8 56 9D
 D6 63 C1 24 02 A4 DB 3E 24 A0 F4 A1 E8 8D 0D 25
 F7 FE 1E 1E 32 EA 42 2B 28 66 5A 74 04 3D E0 09
 DA 87 E1 07 08 3B EF 77 56 32 B8 48 D5 4B 0C 7F
 49 22 2B F6 72 B3 8D 1B 41 67 B2 FE F0 20 DC 0B
 05 85 4D 95 F6 4A ED 35 C6 0B 3C 56 13 72 D4 47
 10 64 15 FF 3D 95 6E 99 4B 84 93 2C 4E D5 4D CF
 F6 F7 19 3B E9 B3 8C 7D 89 8D 98 C7 12 1F 3B 7D
 61 00 8D A0 C1 F4 DA 72 D7 78 CE 25 B4 FB 3E D1
 70 D3 67 8A 21 A0 00 E0 EF CA F9 33 06 1E 68 EF
 20 12 52 32 D6 35 51 F4 12 6B 0F DE E9 CA BE 76
 09 80 2F C3 E7 5A CA DE 0B 68 E3 61 FC 6B DC 27
 EC 50 72 EB 9F C9 80 78 C3 BD 6A 98 8B B3 91 89
 D1 3A 00 12 69 3F 2C 8A CF 20 89 39 52 69 72 3F
 9B E3 23 A5 0F C7 48 A4 95 B6 34 75 3A FC 8F 37
 B6 69 50 76 67 CE 56 91 B5 44 D5 B9 E2 C4 49 DD
 4D B0 F5 AE 57 D5 5B 81 DB BA 59 27 C3 F9 E5 9D
 88 D4 DC 2B 7C F7 C4 BD 4D 3E CF EA D1 6B A4 1A
 49 18 56 D3 27 CD AF 62 ED 91 9A FF 99 8D 1C 09
 2C EA BF F6 9D 8A 91 EC 21 86 1D 7A 9B 03 5B D4
 AC 1F E9 13 7C 0D 2C 3C 1A EB 8D D2 43 C6 22 61
 DC AC 43 B5 EB 26 0F 83 C0 7C 54 1C 7F 7F 6B 93
 AC F7 0B F9 91 D3 CB E4 AB E4 48 1D 31 D1 19 7E
 7F ED 88 EA 16 3B 19 92 06 EC 8F A3 F4 78 9C 9B
 EC 54 4F E9 25 19 18 3E 06 39 85 54 19 1E 28 7A
 3F 0F 0A CA EB BE 95 CF 9D 25 94 3A DC 92 94 6A
 E5 53 38 11 84 89 4C 9A BA D1 8A DF 3B 98 E4 69
 2A D7 61 B1 4E 2D 4C 16 97 CC CF 1F D5 9E 9F 7E
 97 CA 3F 88 A8 B5 07 8B 5F 2C 70 C7 0B 9F EA 05
 05 B7 C5 AE 2E C6 F2 60 B8 FB D7 72 7C 6D 66 0B
 96 7F 53 C6 B7 41 2F A7 00 E5 25 4A BC 57 D8 0F
 47 3C D1 F5 F9 C7 28 A3 65 21 6E AC 59 4D E1 5B
 EF 24 98 B2 8B 77 EB D0 94 ED 9C DB 05 B7 32 AD
 0C 07 17 A3 38 81 2F FA A6 0B BF 93 40 E0 16 A4
 3D C5 FF D6 B4 49 68 E4 FF 92 D2 00 4B 08 B6 63
 C0 B0 E8 E3 E9 82 51 2C 01 62 CD C8 8E 4B CF A8
 C3 9F D8 AC 16 79 7D 91 37 22 26 8F E9 E6 E7 05
 DE 46 A2 50 46 B4 80 D6 59 10 5F 30 12 12 39 C8
 AB 33 6F 5B C8 E1 09 86 4F 28 83 A3 8B 7C 14 34
 13 BA 00 06 51 AE 6F 17 10 78 E1 1F 49 47 EE 03
 6C AD F9 D8 00 D6 F9 0E 9A D3 E4 2A 86 45 B8 19
 6F BB BD 85 88 66 B2 8A A0 5F 73 EC 58 BE 13 08
 EA 9E 0F F3 1D 14 C0 F0 6C 0A 66 80 79 EC A3 99
 97 58 12 8F 1F E7 77 BE A8 1B C2 CC B4 76 AA C4
 0C 2A 8F 00 B5 63 B0 81 40 C5 37 8A 54 E5 FB 2B
 F1 EE 03 69 B8 FC 3C 39 8A 64 D8 F5 16 67 1E B6
 C9 22 DD 7F 9D D9 D5 DE A0 FA B7 54 F4 20 93 35
 D0 ED CC 7F 0F C6 57 8C 11 CE 12 86 A0 DC 1D FD
 6A 58 A0 59 24 33 29 A9 A3 7A FF 74 99 DA 6B 5A
 FE 20 EC 31 93 9D 4C 6A 14 10 9E F9 E4 91 91 A0
 CB 63 98 58 8F B5 0E 11 08 72 1C D9 4E 3B D2 5F
 F9 7F F6 D2 70 94 40 78 88 FC C2 39 C0 B5 BC 11
 06 52 DC 57 97 1A 6F 53 67 D2 A8 13 96 FD A1 61
 DA 38 84 33 50 A4 00 ED 33 69 B3 67 CD 4E CB CA
 79 24 05 16 4B 67 17 17 28 13 DB 45 36 72 D0 C9
 7E 90 D8 91 31 59 44 48 D8 D1 A0 75 B2 45 BE A5
 42 67 ED C0 0A 0E 8A 54 10 DB D7 33 CB F8 0D B5
 26 CF 85 35 D5 C4 88 7D 08 38 79 1D 2D BC E4 66
 5F A8 78 BA 3D 28 13 B5 B2 C5 B7 1D 87 1A F3 AB
 F1 5D B9 AB 84 0E CD A7 40 ED A5 A7 EE B1 88 B4
 18 6B 56 FD A2 4E 25 2D F0 4D E7 F6 32 96 37 22
 29 DD 46 41 FD E3 F4 B8 B5 16 74 23 70 C4 E2 6F
 D7 2F 58 E4 82 AD B3 02 4E A0 34 E7 8C CC 99 B9
 8C F4 48 4D 27 BF B4 DE 24 39 FF BE 14 E1 DE B1
 EB 40 04 79 96 CF BF CF FD F4 C7 57 DB 8C 81 89
 5B BB 67 FC FE F1 C9 30 D6 8E 80 AE 07 30 1D C4
 4B 92 FD 76 80 84 3A CB 4C 64 A9 7D CE AA C9 7F
 B5 69 94 C1 98 1F 62 63 A2 3A A3 CF F5 0C DE 4B
 A5 57 4A D3 7C E2 B2 69 2A DD 8C 8A BE BB 06 DA
 52 D4 F9 CE DD 3C 99 D6 53 59 CC 54 1A E2 9F 2D
 E9 BE ED 04 BA 9D 77 A2 52 CD 99 CD B5 03 E8 3C
 D8 D6 87 0D BE AE C8 C5 AB DC 1D A0 EB B4 23 71
 45 A2 72 9D 9B C4 DF 34 C0 DC 16 70 73 E4 CC 32
 F5 C3 EE D4 F5 F4 6E 46 D2 DB 11 6E 4E 02 E2 5F
 19 2B 3D 2C A8 1F D2 E2 A0 74 63 80 E1 2B 7C 00
 B6 4E 8F 23 E7 17 B4 36 F0 8B 83 53 27 DD ED 5F
 EA 4A C4 F3 53 24 03 00 6C B8 D4 F6 AF 7A 81 E8
 78 B6 15 8C D3 0D 06 5C 18 BD 2B 07 FF 2E 66 C6
 3F 85 EE 6E C1 72 DA F0 A6 17 D7 08 E0 B6 86 3C
 EB E0 5F EB BF 3B F7 32 95 BD 09 D6 BD 67 64 A7
 AC 13 3E 73 1C 35 85 C0 BE B6 8C 1E A4 56 1E 85
 CF 8A 61 D1 DF 03 A2 88 60 35 13 0D 22 A8 95 C4
 7F 10 F5 2A 54 91 E8 CA 66 A6 E2 AE 8B 95 4D B8
 32 8A 9B 82 6D 7D A1 58 78 EB 3E A2 4A 9B D7 1A
 F8 09 BF 1C F8 C4 F7 F8 A1 EC A4 6B 9F A0 33 FB
 F7 FA E3 D6 1A 15 42 A5 70 A1 D9 0F BF 14 02 4D
 FB 3D EF E6 50 55 DD 7C E8 8F 48 72 3C 37 C9 C4
 DB 5F AF 61 88 05 F7 8E 42 49 BD 3B 35 AB 67 D2
 1B 08 66 00 E4 E0 46 41 A0 30 ED 00 7B B1 33 8A
 0B 0E 46 83 86 2C 8E BF E6 FB E5 1C B6 B7 1A F8
 EC CB C9 20 F3 12 91 58 34 DF 8A 96 89 40 15 7A
 FB A6 17 53 EB 78 3D 87 23 D0 62 06 2C 47 B7 F1
 2B F2 27 C4 B1 70 E2 B0 6D 13 5B 78 FD EF EB 02
 F3 F5 4E AD 06 0E DF 5B A6 D1 7C 02 50 3F BB 43
 9C 8F CF 92 7A BA 81 37 AE 30 7E 5C 3A 87 DE 05
 74 66 63 F5 4F 27 93 1B 4C AD 4E A8 A5 C3 34 7E
 7A 37 5B 66 69 22 D6 47 FB 85 B2 FD 88 67 92 A3
 41 E4 83 A4 B1 90 41 1D A1 B5 85 29 A2 E7 A0 1D
 B1 A6 0A FA 2A 25 49 21 CD 39 DB FD 75 BE 92 A3
 28 23 97 FD 2C 33 83 0F D8 23 4B AF 17 96 C1 EE
 C0 4B 07 A8 B2 85 12 17 C8 BB 7D 08 B6 38 B9 10
 A2 B9 9E 7B 76 5D 32 20 AF 95 AA 3F 06 22 DF 2E
 99 A2 77 82 13 1A BD C6 6C 89 F2 C8 82 E9 9C 22
 14 BA 32 1F CB 43 56 55 17 A8 57 4C 4B 0A EB C6
 71 09 99 A3 65 4F 8E 95 42 B3 F7 9F 07 A6 4E E3
 5D D3 26 92 25 C8 60 56 E1 A8 F9 28 3A 1D FD AB
 92 34 E9 FB 5E 5E F0 78 34 98 0C A5 87 CF 6A DB
 45 07 00 EB E1 4F ED 58 0B 85 EA 05 CB 4A AC 9E
 7B 25 29 7A 3B F5 8B E9 98 5D 9C 1E 3C A7 10 63
 D0 08 1E B4 34 14 43 40 51 36 FA 9D EC DF 96 B9
 70 54 4F 99 C3 45 D7 C3 F2 53 BF 50 1E 0D 7E 4C
 80 2D 27 B1 5E 74 03 95 A1 7C 6A 61 06 2E 01 9C
 93 DA FB 82 F9 1C E8 BF 62 56 89 9C F8 90 D9 55
 CB E7 58 33 E6 B2 CB CA 68 38 D9 AD 63 D0 86 2D
 E3 24 AC 4C 31 AB 82 D2 2B B8 11 6F 3D 1E E2 5C
 5B CF 8E 15 ED 05 67 62 7C BA 2B 9B 31 A9 D8 BD
 29 A6 28 1F AD C4 A8 17 5F 2C 3A FD 7D 8A A7 1E
 76 E0 7C B5 6F 4B A8 AA 39 17 DC 85 4B A2 51 5A
 BB DD F5 EE 9F 28 D7 DB 10 FB 1D D6 43 3C AB 26
 3B 35 0B 55 11 74 C3 65 34 33 B7 D6 5C D8 59 C9
 C3 F0 55 1C 8B CD C2 0C E5 35 45 7A 2D DD 4E E2
 A7 50 D7 A7 B7 4F AB F3 77 B9 85 5C E7 D9 B2 60
 E2 77 73 58 4B 88 AF C3 96 94 84 5C 56 AE 64 D4
 EE 69 E2 83 D9 76 1F E1 C8 3B 73 EC B0 37 B7 41
 12 22 D2 8C 06 21 EB 77 5F AA 0A E0 59 7D C9 45
 D1 92 C9 B1 68 2C 42 BF 63 AC 18 A6 DF DB 0D 03
 DD B0 49 EC 5C FD B4 C8 6B 8A A4 67 74 DF 4D 6C
 9B 08 5F CF FA 29 93 AA D2 F4 DD 02 F1 12 47 01
 FE 76 6E 89 84 08 5D 40 A3 E4 EB F5 C3 FA DC 53
 DD 05 1B 54 D4 6A 1E 61 CA 7A A8 F6 25 C9 2B 40
 F7 B1 03 59 68 E6 B9 82 D3 DF E6 E4 9C 51 0F F9
 88 92 26 24 36 C3 F1 2D 07 AC C0 09 86 7D 00 3E
 E8 56 EE E6 7C 39 38 0A 40 3E 28 93 F6 FC 79 39
 C5 B6 DF 91 59 4E D0 27 7B 57 0D 84 9B BD 79 5E
 32 7D 00 F4 78 4B 56 6C F0 EA DC 82 58 10 EC 79
 36 FD C4 0C 88 21 81 3E E1 83 B9 0A 29 01 2D 2D
 47 AA 99 CE 8B 20 7D 05 67 B2 D4 8E 6D EA 6B 63
 44 68 82 BF 94 06 C9 81 7A 3F 15 D0 4E CD 23 DA
 0D 77 D3 F5 48 25 D4 72 48 10 FC 2C 6D 9D 6C 01
 2A 53 5B A3 2E E9 B1 CA FE C7 C5 75 20 5A EA F9
 CA B0 C4 0A F7 5F 09 2C E6 5B C8 CE 0D BE 96 75
 CD 61 13 D0 01 06 2F 16 1B CE 87 59 E9 C2 C9 94
 50 FE E0 6B 93 00 F4 DC 38 61 CB B1 DA E1 7E C3
 D4 31 59 59 23 BC 50 D6 AD 87 1D A1 21 38 E2 0A
 E9 B1 DA 4B BC F0 07 D8 CC 7F 5E FD 6E FA 7E F2
 AA 46 5C FE DB 09 56 FA 19 0D 1B A1 DF 24 9E 94
 2D 56 22 BD 61 32 AB 66 91 91 C0 EF DA 08 1E A9
 B3 29 AF 0E AB 72 D8 E6 6C CD 60 3B B6 0A 27 91
 62 15 51 1E 11 F5 D9 50 1A CA 70 7A E8 0E 1E E9
 37 DD 4F 35 13 F3 6C BF 09 5A 70 CA 73 C5 06 20
 3E 1B 2D EB 17 04 2D 20 C3 42 B2 64 83 3A 6F B8
 70 16 AB 5B 54 2E 35 DD D2 CD 64 DD D5 26 11 F6
 3D A9 A2 A5 48 90 CC 50 55 71 6F 82 D5 8B 99 6D
 E8 4C 29 17 76 81 EB B6 A9 58 09 86 87 6E 61 0A
 2D ED D0 A0 79 1E A8 B9 F8 C3 A4 71 B3 E9 17 57
 E4 7F 0F 0A 44 2C E4 B6 0B 0F C8 E1 8F EC C4 39
 3A 7B 7C 9C F9 DB 65 65 CE 75 56 D2 94 7B 79 55
 63 22 A4 68 05 EF 04 E7 D9 50 B6 D0 80 05 06 89
 50 13 46 66 EA 0E D2 AF 74 56 15 60 0B 77 93 C6
 42 B6 69 0D 59 3B D8 92 97 AD F6 7E 0B AD 2A 15
 C2 08 D6 D7 11 05 D3 8F F6 92 5B A7 FA 01 E2 42
 53 C8 49 9E BC 40 CE 46 E3 8D 81 81 07 C0 E8 47
 65 B4 9D 9C D5 AA 27 ED 15 9C 75 FD 0F 05 8F FA
 61 FB 5A A8 51 83 8D C2 97 70 E5 FC EA E6 84 DC
 4A 79 43 AE D6 0F CB 9C A9 99 31 D7 46 CB 4C 01
 86 6C E1 AB 1A 16 2A FD 86 EE 55 FD 75 59 F6 47
 41 2A DA BB 30 C2 A5 2A E5 FD 8E 2C F9 69 F6 A9
 F9 B9 42 13 27 A4 0A 74 57 1D 47 F9 16 16 4A AC
 CB B7 0A BD 56 AB 94 0C E8 1C 25 AD 3E 15 8E BF
 5C 4F 05 B3 13 A6 78 D3 BA 07 93 D4 50 82 03 C9
 FC 17 41 79 31 56 43 B2 DE B0 78 1E 29 19 5C 8C
 AE 8E BA 18 23 A1 AD 72 35 B3 D7 45 66 D0 C9 0F
 DC 82 90 D7 91 C1 C6 A3 2F E6 47 57 1B DF 51 74
 0B 4D D8 0C 02 9D A7 7B 6E 30 CE 1F 2B 69 6F 63
 63 E4 4C 83 51 B7 EB 68 28 6C 75 01 DB 2A A2 CE
 34 37 D1 39 D0 FE 08 27 81 AB 8D CB 12 B9 55 CE
 A4 7F CD 2E DD 81 7A 65 10 B7 4A 29 0D B7 5E 3A
 C1 E2 F1 8E 35 A8 17 F2 2F 8C 30 32 81 E8 0B 5E
 44 2B A3 67 0D 10 58 CC 63 70 D7 AD F4 5E 75 81
 AC EF 2B 49 4C F7 48 95 B2 34 D7 37 17 E5 97 7B
 4F 5D 7C 63 EE 08 18 AE E1 E4 EE 8A 96 D1 F8 3B
 F2 DF C2 1C 57 E6 94 A3 0A 6D 7B 1B 77 A0 05 CD
 62 AF 46 27 2F 9B 58 D8 BF 0B 18 0B 23 0F 62 44
 10 FD 44 89 35 57 9D 4A 1A EE 67 90 9B BC D8 49
 F1 DE 35 CA 09 4B 91 31 AA DD B5 85 CD 17 A8 9B
 D2 23 A0 16 87 1E C3 C1 2A 88 26 B3 5F 50 D3 99
 9C 86 AB 2B 37 0E B6 D3 E2 71 26 D2 AF EE 9C A2
 2E FE EC A3 D0 C8 76 49 79 E0 77 ED 3D 1B AC 76
 7F 6C 2F 29 39 BF 2E C1 CE DE B8 7D 12 BD 59 0C
 E1 7B 5A E1 1B F9 21 E5 A1 7B 8E 27 EC 12 FB 35
 C3 48 3F 62 E0 D1 34 E9 6C 29 53 0E 06 63 B9 BB
 FF 73 93 2E F5 08 19 FC 1A F0 AA 15 25 0B 5E 65
 56 CD 4C 9B 05 66 3F AC 64 50 E6 29 14 AA 78 02
 71 49 BF E0 26 7C 02 84 00 CC EA C6 95 29 B6 CD
 DA A9 3C 3E BA AD F9 29 5F 2E 5D 0D C5 12 5B 02
 9B AC 39 4F 6E 6A D2 A8 33 E0 FE 13 A0 EA E3 F7
 F2 CC 8D D2 73 4D ED E8 10 BF 98 18 FF 7B 92 7A
 64 69 56 E1 D7 CE F5 4C B4 13 F3 0B A1 DA BE C3
 C1 86 A2 53 75 37 C3 E0 76 38 2C FF 4C FE B9 46
 3D 4C A0 AA 60 34 74 04 0A 9C A6 97 B2 7D D0 49
 3F A9 11 72 6B 6D F6 1E 35 09 F0 3F CE A5 90 E1
 F5 22 F4 BC D3 E4 2C EF 82 13 C0 28 9D 94 D1 2B
 B4 C6 B8 10 59 CA 3A A7 8F B6 6A 1D 72 65 8B 4F
 29 E3 8A C3 FA AD 61 31 F8 43 59 EB 8D B8 AF 23
 71 9E 23 00 53 5C 6C 15 25 64 B9 8B 68 E4 75 E2
 46 7E 3F EA 7A 0C E5 CD 71 0F 9B CE 70 14 47 AC
 FD 16 4A 4C 68 CC 35 83 A2 40 F5 C4 59 32 5A D1
 EB CE F3 D2 57 C6 04 CB A4 F4 C0 35 09 44 EE 40
 11 0D 58 10 5C C0 6C E7 4C 3D E9 FB 9D 6B 5B 16
 74 78 67 28 27 79 C7 DF F6 E5 3E 3A 9A AC E8 0A
 BF 90 8C 3D 85 8C DF B7 78 95 77 9B 08 65 AF 67
 CD 8A 53 66 F7 6F 3F A4 B6 53 7C E3 F8 9A 41 D2
 A9 F1 D5 0E EC 98 A5 C0 4B 8A FA A2 C0 6C 47 7E
 BD 0F A2 FB 79 B8 3C 8D 5E 5E 22 C3 04 C0 BF 61
 04 BB 59 86 4E 0B 3C C7 71 53 7A 88 DB 26 98 5C
 E8 1A 7E 4A C1 A0 0F EB 31 C1 05 EA 3A FF 47 B5
 88 FA 22 7B F0 33 3D 9F 3E 28 B4 0D 44 4D 4E 37
 6C 51 B9 CF C2 5E 1A 5D AF A0 D7 1B 50 42 51 92
 2D 52 BC E3 17 5E 69 02 A4 8F B7 46 41 C0 D8 95
 75 AC EF 5D DA 5D 2A B4 08 7D AF E3 DF 75 02 A8
 57 A6 5D 45 31 71 60 12 33 41 5E 14 3A 1F B5 B3
 F9 54 AB C1 64 90 ED F4 C8 5F 6F 17 E3 07 B7 43
 74 2F 15 52 0B 80 3C 23 CB DE 86 DF D9 65 E3 B0
 F2 04 78 46 E5 E8 15 B5 EC B4 E6 08 55 D9 57 D9
 C9 D0 5C A6 F9 7F 0A 60 80 93 C5 D5 1D 8B 34 D7
 91 A8 0A B5 24 60 F4 BE 09 88 56 7E B6 E9 F0 23
 1A F0 0F F2 4D 8A A9 E9 2D 96 BC D6 6A AF 57 21
 28 8B E4 19 46 F0 0A F3 63 27 AB E3 FA 7F 62 6E
 62 73 DB CD EF CD 85 70 FB C2 B2 1A DF F3 83 29
 4F 4D 06 14 5E CD 34 6F 87 E9 5C AC E7 90 2C E4
 09 5F 38 19 B4 26 23 4B DB B8 23 3C 99 A8 6F F8
 9A C3 C4 CD C1 50 91 3D 2B 88 50 AE 9C A7 0B 55
 08 E4 72 04 75 58 ED 8F DF FE 55 8F BA B8 2B F1
 CD 60 93 03 00 8B CC F0 4C 06 D1 45 8F F8 45 23
 2F A7 26 AA 72 48 AD F7 9B 7F 79 47 7B 4F A7 C5
 9C E0 25 11 34 57 C6 27 11 B0 BE 44 D3 57 17 6B
 7C 6B CE 65 17 90 00 83 4E DC BB 3E 76 8B 78 13
 E7 47 B1 33 61 80 75 DD CD 2E 93 0D 54 F2 2A 59
 DB C6 F4 01 C2 9E 10 60 EC 56 C9 F0 EE 3D 7D B6
 30 1B E4 F6 17 0F C6 07 5A CC B7 84 0F CE 09 8D
 74 37 97 F6 E4 BD AE 57 47 D7 98 95 D2 88 31 C8
 F1 A2 E5 25 C9 45 5D 6A 0D CD DF AA 96 EE CF 62
 B4 0B 57 0A 71 26 DB 53 32 25 8D 2B 88 8E 76 19
 96 28 F7 7A 0F A8 D5 B2 17 45 E7 06 5A 28 ED 93
 3F 1E 8D EB 06 40 A1 7E 10 6B F9 7F 6A 52 2D 09
 F3 4E E9 CA A0 28 28 12 E5 63 6A 16 09 BC 6D 89
 25 06 F6 00 42 5C AB 1B 6D 1A 18 1A B6 9D 8C EC
 13 AF 4E 7F F7 0C 1F 3D 65 6F 56 85 01 9F CE 11
 92 4B E8 0A 65 98 F9 49 89 9A 18 CE 86 5F 82 32
 57 F7 0D A1 99 57 86 6E B8 F7 C1 61 5B 3D 2C D3
 FC 9D 53 63 CE 72 24 CE D0 92 99 7F 4E 01 AE 17
 DB 96 01 4D 0C 66 CA 33 CB 5D FD FA 11 0F E2 D2
 6C E5 67 F0 54 60 82 8A 06 A9 95 95 B7 D5 42 20
 EC 2B D3 22 0C 48 22 58 C0 3B 71 5F 9A C5 43 9F
 A3 92 E2 79 9C 29 4B F5 16 C7 DD 04 84 95 3F 40
 F2 EF 3F E8 61 DB F7 C2 88 5A BF F3 46 81 EE F5
 81 8C E5 A3 CB 8F 52 4B C0 BB AC BE 85 54 8E 19
 2E 1C 52 76 4F 36 D7 AE 3B 3A E2 CA FB 0A 12 08
 3F 0D D4 C0 75 2C C4 4C 1F 88 6A 56 5B 70 71 4E
 9B C3 97 7A 55 0A 2C 0F 2B D2 26 0D 1B 96 D8 9C
 DB 70 D8 E7 48 AF EE 80 A8 9A 84 41 4E 45 03 82
 E2 A0 1D 81 46 81 92 C2 77 60 F8 55 BF B7 F2 50
 DE 8F D5 2E 2D 55 D1 A1 8C 45 A9 9B 69 37 AA 5B
 7E 93 2A E2 2A DD BE 93 E4 E4 DA E2 71 3F BF C9
 6A 45 9C 30 03 2F AC A6 AE E2 0B 56 BF 99 39 C3
 CE D0 F5 AF 45 93 FA 4E B6 E2 31 61 66 A1 5B 3F
 A2 AF 75 12 17 FA ED 45 09 95 74 2C CE 2D 89 84
 E4 30 4D B6 0D 4E 46 5C 48 13 D1 D0 FA 4B AB 74
 19 4D C7 36 46 F0 14 9C 8A 1D CF F2 F2 F1 C4 27
 D6 9E D6 13 78 AA 6E 30 B4 6C C1 E3 25 61 D4 16
 43 B3 B3 DF 97 8C 3F D9 AA 9E BF 60 20 AC D2 08
 1C 46 64 31 BF 20 96 26 45 AB EF 3B FD FD 87 E2
 CB 74 0E AA 03 DA A0 71 E3 A5 CB E6 35 75 13 F7
 24 BB 6E 08 F6 43 08 E1 34 9F CC EE 32 5D 2B 56
 D0 F6 A4 4D 17 76 BD 95 88 39 03 0A B9 F8 EE A3
 9B 42 75 15 6E 66 46 2B 58 E0 D3 E9 4D CB B1 F3
 70 1F EB A5 7C F6 C7 FB 49 60 D7 30 CC 60 9B 60
 DE 53 FB 46 15 5F 81 8A 34 90 00 F9 D3 64 6F C8
 75 68 96 0B C7 41 66 6E 11 16 3A B7 23 E9 1D E9
 C9 EE 5D CB BE E7 67 44 BE 2D F1 A6 63 D3 31 42
 7F 95 17 45 DB E5 AF 44 C6 E8 DC E4 06 CE B1 A7
 B7 36 B3 32 00 E9 4C 3B 24 3A 10 59 B8 62 FA 63
 1B 02 9A 14 EC C0 77 8D 36 26 8C 49 78 6B 6E 62
 60 89 D2 B2 39 14 E4 FB 98 0C 70 0F DF 52 82 D4
 2E D9 29 43 7F FC FF 4A C6 7B 08 57 57 14 93 A8
 E1 E5 90 35 C8 EF 80 EC AA 45 62 2C 49 E2 8F A4
 95 0D C1 C5 98 EE 91 06 AE 44 DC 4F CA 5A EE 41
 E1 77 D0 56 21 6C 4A 32 BD 2F 72 DA 75 0F 0A 45
 E7 3E 3F 56 24 4D C2 06 82 D0 B4 20 01 55 08 EE
 F7 65 0B 96 A4 B5 57 24 9C 46 3D 70 5A 09 5A 04
 94 4C 6D 43 AA 76 F2 8D 9D 7C 51 CA 22 65 F5 AA
 BA 2A F4 16 05 03 A7 40 9B 13 28 15 7B 85 0E 59
 CF 48 31 21 35 7A DC FB EC 19 9B D4 0F BB C3 4C
 71 84 34 91 20 FC 43 B2 B9 4B C2 B7 64 F4 FD 5B
 98 9F 82 CD 7D 6E 9A 05 32 A3 9C 54 F0 93 F8 3F
 8F A2 D5 E0 9A 9D 3B 4B D9 19 B0 30 9E 2D 7D 9D
 4E 7B 2F F9 3A 84 05 96 4D 82 24 01 F8 A8 15 95
 EB D1 EE 69 7E F7 55 66 DE 32 2B F6 83 59 0D 63
 26 79 B9 36 F2 89 51 92 0B 6B C8 22 74 27 5D 89
 7B 06 4E 3F B2 40 CB C2 18 93 10 08 10 C9 BA 67
 F8 C4 A8 DA B9 02 92 96 C8 3A 7C 48 14 B0 F4 2F
 47 88 81 C8 CF 07 9E 74 C9 E3 46 FD 19 7A 9B DB
 D9 05 32 1C 68 4C 01 95 D4 EC DB AB 36 17 1C 99
 0F 12 60 6C D5 47 B8 78 58 4C 64 67 FE FE 50 2A
 AD 25 8D 26 BF AC 3F 86 5C 29 E3 4F B5 3F D0 D1
 CA EC BC 5E DE 87 99 9E 44 25 7F C0 C7 08 27 9E
 37 DF 65 60 57 91 3F E9 B9 11 FA 7E CD 92 DA 62
 6E B4 92 C7 BC B7 E9 DA 30 8E D2 E5 D4 64 DE 07
 14 1B 7F 2A ED 5D FE 3F FE 32 16 6D DF 7B DE 4F
 3B 75 4C 0C DD 15 83 47 B9 8A E4 43 BA C1 91 0D
 A5 B1 F6 E1 D6 48 82 0B 41 E2 E7 72 1B 31 10 25
 C1 2C 79 41 0A 1D BD B1 90 73 4A 10 70 B7 8C 55
 1E DC 7B 05 62 8D B3 36 AE 8D DD BC ED F0 EA 94
 3B 7A 87 42 52 96 75 17 1A DE 4A C5 C6 E1 3C 89
 97 D1 AB 30 E6 6F 39 56 6A 3B 4D 6A 10 06 F9 9E
 49 28 2E 2B CE D6 D0 02 39 4B E2 14 3C 98 66 AE
 25 65 C0 C2 C8 0E 8B 49 C8 40 16 EB 1A CA AB 47
 33 98 DA 55 A6 5D C3 EE A2 3D 61 01 0C 52 66 BF
 BA B1 39 3E 3A F7 CC 9C 56 9E DC F6 AF B2 41 94
 28 72 D7 BE A5 93 2A 89 B7 D3 98 BC 91 FE 28 DB
 04 96 0B 2E 1C A6 3A 0D DB 21 FC 67 E7 8E EA B7
 67 18 20 88 60 88 97 2F 6B 6E 0D E1 20 8F B4 1C
 5E 48 89 77 1A 11 CC B6 C4 AA 58 4E 31 C1 CD 39
 27 2C 0A C2 6F 0A A8 5B 5B 73 5F F3 41 A1 C0 7C
 E6 BF 42 BA 39 AB 77 35 F3 CC 7B 6C 09 4D 4C 34
 2E 11 17 1F 2B B8 00 64 44 EC B8 9D 33 90 6E FB
 06 A6 B3 2C 86 DF C4 97 CB CE C8 CE 4D 1C 57 F7
 48 36 0A 08 28 36 B2 47 67 E5 60 29 67 9A A6 8E
 2A D1 3B CB 7B AF FD 28 76 67 7C 19 BB 6A 82 41
 A6 D3 27 9C 27 A9 54 F6 3C 34 D3 AB 99 8D 60 06
 D9 D7 96 5A 42 38 A5 A7 1A F5 E7 FF A7 0B 3B 5A
 3D 98 52 9C 51 38 AF E9 77 83 6D AF 9C 21 CA 75
 F7 B3 66 9B F1 CC 83 3A E1 7F 5F BA 45 87 3F D6
 07 B0 3C 08 67 74 61 30 91 AC 51 AB B3 2D 53 CE
 8E E3 84 14 48 53 B3 49 E9 6C 68 48 AD 7D 33 20
 6E C7 B1 FF FC 90 94 D5 B7 2F 29 39 5C 9F 55 A1
 35 88 68 1A B9 55 6C CF 93 6B AC 9E BD 89 8B F0
 13 22 78 EA 2A 46 9A 37 6B 7B EC A1 BE B4 D1 2B
 DB 62 1F 16 3E 32 9A 14 97 33 F6 37 1D 72 76 CB
 32 D4 15 44 9D 50 F7 FF 3B E4 F1 30 C6 54 FE 77
 B3 A3 19 FD E0 B1 CC 3C 65 92 87 3F DC 23 4C 9C
 0B F4 7A DD 18 21 36 F5 42 C7 28 27 5F 0D 89 E8
 DB B4 AF 4D 62 30 83 05 E0 62 F9 B7 C4 52 49 7C
 12 9B 3B 9D 99 89 EF 67 B8 E9 8E ED CA 75 BB 79
 97 41 06 4B A1 4A 43 8C 09 DB 7F 2B AF 49 23 FE
 9B A1 35 ED 31 00 22 2D B9 5F 8B 71 9D F1 2F 7B
 43 42 24 38 86 3E 06 56 DB 35 85 87 E2 51 63 4C
 29 AF 69 A9 1D EB D9 A1 02 42 63 C1 61 B6 CF AC
 DD 2B 78 76 3B 0E 7C A0 D7 71 44 FF 24 0B 36 50
 47 10 CE 1E E1 BB 3E 8D 43 F7 D2 8E 47 69 91 40
 DD 5C D9 4C 4A DD EA C6 B6 1B 17 83 C6 DB CD 8E
 B6 9D 6B E3 26 BB 55 29 B0 C0 9E 27 C4 CA 74 67
 EC 75 E1 B2 C3 8C F7 A8 2A 79 7C 8F CE F4 49 CF
 BE C2 B8 8E DE FF 4A C7 15 C5 06 7E 88 B2 C9 DE
 7F D8 98 9E E0 5C 64 80 3B 6B 00 A1 D2 74 76 D3
 9B D1 CD 61 59 47 86 C5 D2 1D 2C C9 7A 6B DE 30
 AE 73 FB E9 0D CC F7 E7 85 C8 2F 32 0F 4D BC F8
 39 49 F7 ED 3D D4 BC 7F 81 3F 28 56 A6 D7 F3 CE
 58 59 CE B2 1A B4 BE D5 63 5B 69 E6 AB CF 0A C3
 95 D1 5E AD 0E FF 6D 56 AC AF 97 4E 06 18 30 AA
 C9 2B DD 2D 4E 7B 72 D5 A3 93 E1 EB 92 1E 66 DC
 82 EF E7 A2 16 65 BA 1D E7 80 D3 6D 2A E8 28 EE
 AB 0D F6 3F 9C 44 A6 27 E5 21 A1 25 11 CE 25 64
 2A DA 6E 2D CB 96 90 4A 6E EA BD 2F 96 4C 8B 6A
 12 5E 64 E3 BE 9B 4F 9C BB C9 89 DE AF EB E4 92
 DE 29 2E BC F2 B1 65 EB BF FE 2D 8E 9E C6 63 74
 7B DB A5 F8 1E 92 EF 43 4A C0 6D 83 1F B0 A3 2C
 9F B0 34 E6 89 26 72 95 19 36 1E D1 1A C4 6E 58
 16 B0 C3 B7 DE 91 01 41 EC CA BC 93 12 C5 9F 6E
 B6 38 2B C3 0B 42 37 D3 74 B2 7E EC 48 1D 76 35
 5F B0 6D AD 49 3B 8A EB 8C 8D E2 DC E4 1E D4 F5
 55 69 7E E9 26 55 99 A1 0D 56 38 8C 73 76 79 1A
 39 C4 AF 87 B6 57 7E EC 77 12 CB 9B 1F EB A4 D3
 C0 2A 9C EB 4D 77 E0 1E B8 C2 5F 06 E4 6A 9F 7A
 32 B8 79 41 E4 A2 D9 96 B6 0B F7 B9 A3 18 07 2C
 30 E9 B4 2F EF 11 39 05 04 D7 E3 3C F0 C8 80 7A
 4E D3 93 F4 4A E1 24 E1 7D 89 AB FA 9E 9A 97 A6
 1C F7 58 C2 8A DB 9D 46 41 FF 3F EF 11 60 BE 37
 8B CC 95 56 D5 16 7D D9 88 5D 0F 8A FB 4E 33 C4
 85 B9 4C EF 55 FB 61 21 CF 45 28 8D 33 90 8A 5D
 17 7D 78 FB 47 3E 63 29 0F 01 64 72 E0 97 FF FB
 DD FE FC 50 F5 D1 D9 5E 50 8E EE 7E 65 DE 4D 40
 4D 9B 8C 52 0E 43 1E 33 CD 58 42 8E 87 47 37 53
 2F 4C 47 4B A7 27 7F AF 11 7D C6 32 2D DC 9F C7
 2A F6 69 2C 15 2F CF 24 AA 04 4D A7 8D 8D D2 60
 25 F1 7D B9 6C 2A 41 3D CD 59 3B C1 FB 30 73 3A
 6C 73 AC 22 54 06 66 71 96 82 3F BD 76 C0 0E 81
 C4 C0 41 0A FD FE 3E 8A 0E 70 BB 28 A5 C7 0D 85
 DF 24 00 BA 58 2E B7 67 E7 62 BF C1 39 7D CD 29
 D0 6D 74 8F F5 2F 83 64 13 1B 73 B5 72 7A 59 0D
 10 13 A0 4A B6 1C 1B 86 41 AF 60 D1 3C 7E D9 C8
 D3 1B 12 77 83 FB 00 6D 82 D3 A7 D8 BB E6 C5 EF
 7D 97 79 24 EE 1E 11 68 30 56 A0 50 A0 FB 9E DA
 57 D2 11 07 07 16 D1 E1 F1 75 70 89 EA 3E ED 41
 CD 97 63 2D 25 0B B6 39 BC 40 3D 54 93 16 71 A0
 10 17 7B A5 C6 1D C4 D3 6D 6D 15 ED 80 E0 1C C8
 9F CA B6 31 17 AB FC 7A 16 9B F6 8D C9 5F C7 EF
 28 E0 C1 6D 75 9A 88 6B 05 C0 64 14 FD 81 37 5A
 50 E8 56 25 7D 9F 91 E6 8C DE A5 3B BE 55 43 85
 07 9D EE 76 9E 3C 80 80 B4 C4 DD 4A F3 45 2B 01
 58 51 DD E3 C9 AF 35 A9 76 84 BE 03 C5 31 7D DC
 7E B2 9A 41 27 15 37 F8 93 8A 7C B4 0C E9 41 83
 E5 D3 EC 7D 03 CD 6A 99 52 05 67 79 F5 3D 7F 64
 E8 B4 DF E4 DC B9 DE 83 0E B8 E5 59 67 98 BF A5
 19 B6 C4 D9 E2 06 54 52 3E 95 5E 6D DB 4B F0 90
 D5 82 52 43 FA 70 C0 87 B6 F4 E5 E6 43 49 1D 8B
 02 5E 34 A8 CC 56 4E 4F 90 A0 85 ED D7 69 AE AD
 65 72 9D 48 64 60 A5 1E 45 DF CD 3D 77 D2 68 96
 EF 06 0B 73 30 D9 DC C6 92 E3 12 AF F1 6D 98 DA
 5C D5 A9 DB C4 6B 0B A2 A0 42 64 A9 8A 5B DA 5A
 A9 81 19 35 95 D0 9B B7 5F 4B D9 3A 13 88 A1 E8
 55 88 C4 77 BC 72 05 33 B1 78 67 41 17 93 48 CF
 3C D3 B2 62 05 B6 EA A2 E0 20 90 74 9D 59 94 4D
 AF BC CF 97 46 A4 83 79 50 C2 19 08 E5 9E 00 BC
 7E FD C5 CE D1 26 8F 11 0C B0 EF E2 00 9D 3F 10
 B2 ED B3 13 4C 48 61 BB 05 27 8A EA 24 79 1C A2
 93 15 8C CB 26 F0 C2 26 BF 82 FC E4 29 1D F1 1F
 92 37 F3 15 84 C7 10 64 CB 45 C2 2A 0C 8B 34 94
 C4 97 08 3B 72 07 F7 4F 8E 39 D3 27 4B C6 A7 9C
 F3 A2 CC 6C 17 C0 59 96 2B EE 15 6B 19 93 AB 0A
 B2 6B 81 FF 58 DB AF 34 46 BA 18 C8 2D 0A FF 27
 42 78 01 93 20 D0 1D 30 1E B1 EF 81 9E 65 C4 95
 EB 72 A2 DA 3E 3C 7D 3E 12 B6 11 FA B6 51 F5 36
 FE 91 FD 05 8E 86 9C 30 2D 6F 0E 58 05 D2 59 13
 86 62 D9 57 4F EC DC A9 93 ED 94 15 CB EA 68 21
 F5 E9 E7 CB 51 65 C2 D0 98 F8 D2 C2 A1 94 E3 E4
 36 1A 2F F7 E3 AA D8 E1 13 C7 87 F0 AE D0 64 FF
 09 1D AB 22 EF F1 E0 6A A5 78 DA 88 80 06 6F 1F
 57 44 9F C2 BA 9B BD 83 78 8C EE 79 12 3A 77 49
 04 65 CB 6B 8E 5D D5 34 D3 31 61 95 71 82 55 80
 C2 42 F4 70 C2 30 30 6C BA 54 2C D7 19 B6 F5 6F
 53 57 8C AF 49 2F D2 CA 4B B2 6D 22 1C 5D F5 C4
 43 AD 96 73 3C FA 66 38 B6 23 B4 4D 1D CC D3 C9
 95 33 66 9F F5 6D 10 98 BC 9C 5D 62 BA 93 3A CA
 0E AC A8 73 E2 1F 58 72 16 EC 40 E4 75 CD 17 B2
 0E F7 FF 72 1C C4 C6 18 11 61 98 1A 72 84 F7 5C
 8F 26 C5 F7 63 4B 20 8B F2 47 EB DA E4 38 E5 E2
 8A 34 E8 A4 AC D6 96 FB 71 60 B6 D0 14 93 19 C5
 06 FA 48 D9 D1 39 8D 15 4C 4A B9 DF 16 62 02 06
 02 DF 44 78 0B 32 DF 15 BF C8 6F FA 17 03 E0 72
 7B B8 C1 4A F9 E8 1E 67 5C B4 F1 2C AC 72 FA A9
 CF EF 89 B4 FF 13 56 74 5A D4 AA AA 56 A7 6B 26
 91 B2 F4 52 07 37 81 0E 37 D4 94 58 08 2D 65 27
 45 CC E7 FD 37 5B 67 02 33 21 96 E2 D2 FC 95 C9
 C6 00 96 AF B3 EB B4 33 79 EA 59 53 45 A3 E2 D2
 63 2A AA CB C6 8C F0 8C AC 34 58 37 E4 C4 74 73
 E0 5C B8 50 32 7D F9 29 7D AA 25 D0 72 8A 35 E4
 AC 3A 9B 40 EC 07 07 7B BE FD 22 D0 19 79 8B 9C
 E3 8C 3C AB 86 CD 5A 83 BF B8 C0 62 99 C3 79 47
 B7 C8 35 76 C3 5F 5F 09 F0 2A 58 05 9B BA 01 BA
 79 F7 6F 60 A0 2F 6C 7B 92 5D 66 F5 16 55 5B E0
 83 37 22 91 F8 B5 05 FE F9 E5 04 6D BC CB 27 CB
 DB 38 82 09 E8 C1 49 23 74 AA 82 E9 F2 33 B0 21
 9B 76 E0 9C 3D C4 AA 4E 06 37 73 34 FA 96 01 7B
 DA F5 3C BC F6 34 69 C5 13 A7 B3 65 05 1C B8 D6
 19 A5 80 BF B8 88 35 ED FB 39 F9 28 55 ED FF 56
 71 B4 D2 97 D5 8C 84 60 CB 6C 12 07 0A 8C 77 68
 2B 4B 71 83 5C C7 2F 5E 6C 51 0A C0 AA 01 01 1A
 87 58 97 AD 8E 59 E0 11 49 B6 3C E2 58 71 2C 5C
 7A CF 82 84 AF 2D 3B C9 67 9C 7F 06 25 5D 08 17
 C0 AE 3B E5 DF B0 B8 A2 31 C0 DB 6E 8D F2 70 57
 04 A4 48 01 DA 8C FA 56 C6 B7 FB E0 AF CD 15 E0
 77 C1 DE 4A DF 62 CB FF 9E F8 37 A3 C1 A4 6F 6F
 18 FC 0B 40 22 EA 33 07 F0 C2 B2 45 EB 27 D2 61
 B1 CC 90 BF 14 83 B2 FE 3D F5 EB DA 22 EA 4F A9
 4E 49 8C 68 E1 04 AC 9D 06 22 02 D3 9C 77 4B 02
 A4 CB 0D 9B 50 32 75 87 26 66 1E 17 E5 0F D5 D2
 C6 27 77 61 04 96 E3 6B E1 F1 5B D9 C1 7F DA 8F
 04 34 7B 3C 0F A4 20 64 20 2B ED 87 32 A3 58 1D
 78 DF 72 23 F7 9E C8 92 89 37 90 8A 69 55 DD F4
 49 79 FB 7A D5 D2 81 AA 2C 3F 13 34 7A 26 9B 27
 35 45 0B C6 06 7D 84 2A 7F 87 0E D4 AD 81 E7 AE
 53 7F 57 02 BB 2D BC 7F 79 B2 C5 46 18 90 0D AD
 E7 5F 6B 46 B3 6C 4C 4B 90 F1 C2 A3 AE CB 40 B0
 F2 93 EF BC F4 44 CF 40 57 77 D6 C3 43 C4 FE 77
 60 B0 BC 58 95 45 80 4F D1 19 EC 77 6D C4 2A D7
 AB 73 83 22 DC 55 E4 C7 D0 AA B1 C2 0C 3A CD DC
 55 82 19 83 EE 8D 80 B5 91 08 39 61 34 47 2E 04
 AD 16 10 EF 62 67 C8 7C 22 C5 87 5C E2 6F C3 CB
 1E E5 72 16 AB 14 DA 43 D6 20 D4 9A 3E 4E 24 D3
 70 B0 94 87 3A AF 5E 79 3D 5B 81 17 3B 02 50 FA
 92 C9 98 57 2B 54 DB 5E 05 63 D5 F5 8A 8F 63 1D
 B0 8F 1F 5D 27 5C 94 93 E0 4C D1 4E 60 D5 C5 84
 D4 5A 1E 24 C4 C3 E2 30 73 3A D4 97 E3 FC B8 22
 D5 73 5C F1 27 34 AF A0 B8 F9 82 58 0D A4 E1 78
 E7 5C E8 18 CD A0 D0 CF 2E 02 17 03 59 85 17 8E
 EA 28 00 E7 20 98 30 47 AB B9 F4 AD 42 DC ED D3
 87 71 8C 42 EE 54 8A EA 73 B4 4E E4 4D 1C 30 4A
 71 B2 60 3B 74 9D E2 22 F8 95 FE 39 76 4D B6 27
 C0 49 7C 9F 16 58 92 A1 5B E5 CA 87 20 2F 63 C4
 C8 C9 17 33 D8 9C 1F 18 06 B2 99 8B 51 EB 2A E3
 48 7B A6 E6 63 23 CA B4 ED A8 B3 90 B5 D7 40 B2
 70 E9 03 FA F4 19 DC 27 26 23 54 5C F1 A8 62 86
 E7 F6 6E C2 F5 08 C7 AF FF 56 41 A2 64 0F EF 85
 C6 E7 96 38 55 F0 7E 08 E8 F5 49 6C 04 2B 48 2D
 E3 67 CE 5F 4C 00 28 6B 01 79 17 65 D1 E9 2B 78
 3C E2 A2 03 AC 96 B9 BD A8 E8 66 E1 F0 AF 1F 1D
 4E CD 08 21 AE 31 63 D8 FB EC DE 9F 26 75 70 F8
 20 EF 0D 97 14 81 2C 25 8C 76 88 6A 25 C2 E3 33
 61 BF 91 41 2E E1 13 E8 9E 73 E6 02 46 5D F7 73
 69 16 91 72 78 21 83 A8 20 E0 9D 05 C5 7E 40 E7
 97 67 48 FF 46 C4 3F 0B 09 8D 3C A5 D8 EF 31 E2
 40 2F 09 6B 4E 8C D5 DC 74 36 EF 3A A4 E9 23 96
 2C D1 F7 8B 03 60 97 BF AF 95 4C E2 64 9C 61 75
 E4 04 C1 6D F2 E5 92 07 98 E1 FD 5C C7 11 73 F3
 E5 FF C1 F0 A2 C4 F9 86 9C BE AF 1E 57 32 AA 35
 9A 50 6B 08 C2 54 09 40 3B 89 92 96 43 A0 5D 28
 4E D3 68 29 A3 48 70 33 20 0D 35 5B 10 4D 4E 8C
 8A 82 5E F6 C7 BD C3 C8 87 EE 25 38 C9 E5 79 87
 EE C0 6F 61 BC 19 92 EE 9A 7A 58 05 94 88 69 B9
 50 7B 84 C0 0C 61 9B EC FA E9 DD 41 AE D6 02 F5
 45 B9 5B 0A 7D 0C B9 62 0D 25 39 25 E0 C0 DC BB
 A1 CE E9 66 7C 11 5D 64 46 1F 0D 48 F1 95 14 9F
 16 B3 1A C2 EA 39 F8 15 B8 B2 5C E6 97 77 D8 1F
 20 6F FD 94 8B 4A 53 F9 E4 80 AB 9F 2F 7C 20 59
 71 80 DB AD C9 DF 85 D1 3F 81 AF E5 54 68 E9 64
 92 D9 6F AE D5 6F 0E 70 A0 2E 3F 9C 77 71 C4 89
 DB 5E 3C EC 83 65 BB E2 B3 51 5F F4 C3 2C 1C FC
 0E 86 65 A0 2B DF 3B B2 60 73 7E 7C C0 D1 8F 3B
 B3 7D 26 86 DD 42 D8 7B C2 9D B7 87 A1 F7 52 FA
 2C 98 12 1D C5 EC F8 5C 47 62 08 04 5A 51 7F EF
 A9 32 ED 85 58 7E 34 4A 15 80 D2 46 7E 06 84 44
 23 83 B5 9A 85 C6 6D F3 5A B4 20 31 B7 C2 CD 57
 C1 1B 13 A6 23 AD 83 E5 F3 3E 59 D4 F2 78 E1 EF
 1B 3F 48 03 E7 50 1E E8 00 21 61 F7 B8 8B C7 7F
 76 00 CE 4E 7A BE 03 B5 50 14 0C 6B 1F 36 1C C5
 91 58 2F 99 5A EC 45 31 54 18 C2 83 C0 2D 36 18
 CB 08 74 1A 7C 93 5D C7 B6 37 87 5B DF 3A DB 25
 B4 9D 17 62 57 76 87 64 D0 3A D2 35 67 56 96 F6
 AE 8E 6E 4E 60 25 6D 40 46 59 02 FC 52 FD 51 1C
 DB FB 65 CE F2 F0 F5 36 B8 8E 71 BE DF 0F E8 DC
 33 DF 3F 60 0A 39 FF D6 7F 35 D2 90 AD 12 2D 84
 8E DD 35 38 4C 07 15 FA 97 B1 30 D0 77 45 58 D5
 26 B0 9E 46 F1 1B C1 14 DF EE 35 DD 43 1B E5 04
 9F 85 82 27 45 43 0D 06 0B DD 77 3D 54 34 E7 E2
 F7 89 AB D7 87 B1 24 CD 67 90 27 D7 B2 2A F6 27
 1B 5C 03 B0 4B B2 FF C2 DD 3C C3 CE 26 23 8C 42
 9A 4B 05 8E D1 8A B0 58 1E B3 A0 4C 76 6E CB 7E
 85 79 9E 7E 15 AC A7 E3 33 BD F4 C4 D0 2E 94 03
 73 6E 0B C0 8B B2 0C 6B 1B ED A5 96 14 39 3E 06
 1A EF 09 D4 E9 0C 50 99 67 D0 75 DC CB 7C D1 19
 9D 9F 60 63 31 7C 09 65 E2 CE DB A0 9B C1 B0 95
 EB FD 68 E6 0B 73 11 CE 86 B4 CE 23 D4 91 A7 C9
 CC BB 62 73 E8 80 22 84 16 47 0E 5C 3C B5 B1 BB
 BA 73 49 00 D8 18 54 7B 64 4F AA 9B 33 5C A5 0E
 19 17 6A 0E C0 B4 0C 94 4F 03 D3 33 FD 7B 2C A6
 CB 8B F1 AC EB 9F 28 44 01 99 D2 9F F2 71 A4 3A
 2C FD 44 E4 9C CE 82 3E 19 50 DB 3E 9C 21 5B E1
 F8 71 3E 30 BB 5D 6F BD 38 F7 F3 F0 5A F8 2F E4
 CC 18 6F F5 01 5D BE 0A CF 2A C5 5D EA 23 FE 61
 61 98 07 53 51 DF 5E 02 DF AF 6A 70 8C B6 17 23
 AC A6 2B F3 F8 EB 9D F1 8C A7 66 B8 61 73 A8 19
 9F EB 1E 94 9F C5 F3 BF BF CA A0 2A B7 E7 94 22
 C3 55 2F C4 E4 66 D1 64 EC F6 59 E6 41 DF EF 56
 A0 53 CB 7F 38 F4 24 89 61 74 AB BA 4A 57 45 8C
 1C 96 C2 29 3F 4A DB 66 C8 01 3E 7E C8 26 D4 02
 27 8F C0 48 CF 09 BE 28 D6 22 72 40 44 8C 62 A1
 0D FB 41 76 93 AC 23 4D C3 87 B6 BF 7D C6 F0 DA
 D1 B8 75 C9 FA C6 A9 76 64 7A 2A 0D 3C 43 7E DF
 D9 D5 46 B0 AA 29 1B 34 0D F5 EC C2 E4 8E 55 14
 16 ED 3D 41 BF F5 77 17 E7 A0 20 0B 17 70 4B B8
 41 4E E1 FD CD 25 A9 54 8D 57 8E A1 F2 87 79 C0
 47 0B 86 58 10 5D 89 48 FD 6C 00 72 85 D6 F5 82
 27 F4 CF AA 68 7A DF 5C AF B8 80 E7 75 92 04 18
 09 92 3E 18 5F BF DC A1 AD A7 CC 89 D5 E9 A3 96
 A4 7A 67 EF D9 B2 D5 C9 48 A6 C0 3B BA E6 9C BE
 0D 47 DB 13 07 45 7D B9 CD D5 C5 A0 0D 13 FD 1F
 13 51 AE 8E D3 7E 8F 85 F0 76 4F 8E 6C 82 D3 DC
 11 A5 33 0F 0C 19 E8 20 B9 98 96 F8 D2 49 0B 25
 7A E6 5B 21 04 CB 8A 38 45 85 1C D3 7A A9 48 21
 37 48 A3 6A 81 C7 29 49 5D 3D B5 65 35 3E 58 8F
 38 0F 7C 3B 52 47 40 F1 FC 3C D4 BE B4 26 24 2B
 C5 91 3A B6 7E 4C F8 CC E5 84 29 37 C0 EF 05 30
 32 8F 9B 6F E2 1F AC 48 A0 2E 73 59 D2 8B D1 41
 74 97 B2 3C 58 E3 3D 79 DF 5D E5 9A B5 9D B9 18
 5C AC 81 CC 29 30 D9 B9 F2 60 12 07 B3 C8 B7 DC
 AF 69 D5 84 98 01 0D 9C CE 07 43 E2 10 89 9D 39
 3A 2B 49 11 72 A9 E9 E5 97 45 AB 3B 57 BE 2C B0
 A0 9B AA 1F 75 AB F3 89 D8 C1 54 86 65 49 7C B8
 18 AC 5D 50 86 1E 1E 62 27 E9 A7 22 4B C8 FC 9F
 B6 73 71 CD 8C 11 29 2D B6 E7 D1 50 80 DF BE 25
 F1 A5 9E 79 B6 64 C7 86 AD 50 85 03 75 97 00 13
 12 1E D9 02 D3 81 2D 82 3F 5F 90 71 C0 1C B4 63
 C6 41 A8 1F 90 41 16 37 4B 5E E6 6D 77 E9 81 2C
 20 D3 18 73 37 BF 47 D2 2F 26 61 5E 7F 60 3A 62
 CF DE BF CB F1 02 B8 F0 0A A4 0C 9C 3F 05 5D E3
 BE 5A A6 54 46 81 E1 D0 E7 6F FF 4F 80 39 0C DC
 3D 85 72 70 E3 F1 1C D1 F1 77 A1 1B E2 7E 23 78
 18 05 59 06 C6 1F CF 8A 6C 00 05 E7 EE 4C F8 1B
 32 10 FE 2D BC 96 7F 50 79 D2 E9 CE 5D 79 F8 98
 19 DB A9 4A 88 03 69 A8 67 D1 BA B2 23 35 05 EE
 02 3E 0B 66 F6 B0 B3 43 C4 78 18 44 CA 86 54 22
 57 2A C8 B3 78 18 95 0B 5C 97 03 2D 07 C6 00 B3
 C2 49 E4 53 3E 2E 19 5D 41 FB 86 AB F6 58 A6 5A
 3C 75 DD 1F 39 3A 74 C1 E1 31 0B 00 63 7C 52 D1
 22 ED 2C A0 34 22 68 46 25 50 13 66 44 7D 05 C8
 B4 58 81 16 C9 30 CB 38 4C 77 0D A3 37 E6 79 64
 55 62 17 4B 57 21 88 59 5F 4D 5B 02 D1 6E 5B F9
 6C 49 BA 70 01 52 94 E5 5A 7E 85 C8 63 88 1E 33
 9F A8 88 D9 B1 73 7E EE FE 4F 0B 85 E7 71 00 2F
 CB 8A 23 74 FC 64 99 AA C5 34 32 CC B4 D3 6C 57
 59 03 A4 A3 3F 5B B6 4D C9 21 FE BF 08 A5 E4 4B
 CA 0D E8 42 A2 33 4A 10 A3 5C 4C 40 3F 56 3E E7
 D5 F4 49 42 6D D2 81 C9 C1 1E 9B 99 3B 98 C0 8F
 E6 D2 CA CC 5B 38 5D A1 D0 90 D8 E4 3C BF 56 B3
 D4 DA 93 CC 6A 97 AB 2E D8 DE AC 6F 24 A2 82 53
 C5 4B C4 B2 98 CF 49 F6 45 6A B8 05 7F 14 2F 9B
 87 28 7B 67 0F 2F 2E 68 D0 0A 99 2E 84 06 43 06
 56 F7 6D 57 E3 1A 8D 0F B1 36 A3 AA D8 EE 97 BE
 A3 FD 6D A4 B9 FF A9 22 64 F1 B9 35 7A 89 A2 6F
 9A A5 69 EF 4B BC D8 B5 4F 89 32 F1 B7 17 F2 8F
 5A 8C 70 44 F1 B3 93 11 E0 A3 ED 91 71 D3 E1 FE
 66 14 4F FF 72 C0 75 90 F0 93 D7 34 97 67 EE 1A
 34 03 F2 91 74 04 71 41 15 FE 5C FD D8 28 98 E6
 C2 7D 42 C2 9A 85 02 7F 24 A0 48 6A 69 4C F7 6C
 60 16 A3 89 3C FB 0E 0D 99 1F B0 0A BC 42 78 64
 B1 A9 47 F7 7C 93 F5 87 40 25 97 28 93 97 93 79
 E4 85 F1 55 D0 EB 85 4F 2C A4 53 4E 9D D8 96 80
 B7 68 61 E9 F0 43 25 BA 13 AB 6E DF 47 83 1A 21
 A0 86 92 6C 11 11 F2 64 C9 A1 97 F1 07 E7 60 B1
 34 07 9D 8F 24 3A 49 E8 32 05 95 12 C0 82 15 45
 59 BD 62 57 C2 B8 DB 1A C5 E8 0F 8D CC 2E 42 61
 8C 51 7A 15 C3 38 81 8D 54 48 E0 0E 1D 9D BD 54
 52 A7 30 4E 8A AB A6 8D 67 4C 1E C4 1C 80 4D E7
 4A AF AC 5F 58 19 9A 2C 37 7F 4B 6A E5 E0 4B FB
 E3 C8 69 8A 4F 64 1B FF F7 CA CE B1 72 9A 92 22
 46 CE 1B D4 CC 7B 7D E5 64 C4 F5 BF 98 07 DA 61
 AF 4C BA D3 B0 C5 74 50 69 83 6E C9 CE C6 BD CB
 AE 65 42 C7 2C 97 30 E3 D2 46 F3 2F 83 BE 91 B4
 8E 59 D9 2A AA E7 08 29 70 A3 C3 EC B6 33 D3 8B
 F8 C9 6A 9A F6 68 23 B1 20 7B B9 98 25 26 B4 48
 40 D3 68 CD 6B 92 CE 04 A8 09 9B 7D DC E5 0F A9
 D6 79 FC 05 B9 F9 D7 57 DB BF 64 C0 C5 F7 2B 00
 73 E8 69 15 DC B9 DD 9D C8 C6 F3 E5 BD FB 92 01
 D4 6A CB A7 0B 6B 93 53 E9 60 EE 5D 30 44 EE FB
 57 7D 65 19 91 66 39 97 81 58 BE 2F 80 83 1B E6
 74 E9 B6 BE C1 71 42 62 74 93 AA 4B 25 19 42 34
 47 A3 82 D6 5E 77 28 A7 08 01 45 75 8C F3 EB 81
 EB 5D 79 F3 C1 BB 90 A5 B7 B8 22 62 58 4A A3 CB
 60 73 EF 99 95 80 22 FB 7C D1 E8 1B 84 5A 0C BF
 2C 09 2B 46 3D F9 CB 6F 52 75 43 1C BF 33 F2 FF
 12 D2 10 E7 2D 1D BF 8B 4F E3 29 C5 E3 79 B6 9B
 DD 8A ED 28 37 E8 18 16 99 63 E1 02 31 63 3E B5
 B8 9E 0E 6B 7A CB DE 68 2C 76 BE 09 F7 00 36 48
 11 F7 AA F8 1A 7F 20 F5 9B 17 70 22 2D 57 C2 29
 58 27 91 43 14 B3 08 E7 71 53 BF CD 0A 47 3C 17
 82 40 ED D0 49 12 C2 D8 69 07 9C A7 5B 81 E5 70
 73 69 69 13 61 5E 81 15 CC 49 0D 8D 16 4D 87 66
 8E 9A 45 5E 48 E5 23 6E A7 F2 F3 B7 A2 C2 65 A1
 BE 9E 9C 53 8F F5 BF 72 9A F6 F0 CF DC B9 05 B2
 AE DA D1 D8 82 DA 19 C4 9B 43 46 7D 40 B2 4D C5
 91 24 EC 0A 5C 91 9D 51 3C 09 FB EF BB 92 50 8C
 BD 09 51 A6 90 C9 83 BB 58 EE D7 0A A1 85 F8 E2
 5D F7 E9 59 B6 C0 84 D4 0E EB 8F CA 4C 47 96 56
 8A 9D 6E 85 9F 7E 62 C0 48 9C 7E 48 8B E0 1D 4B
 FC 9D 68 FD 00 74 72 AA D4 06 82 86 3E 53 4D 5F
 4A 1F 69 2D 31 E3 30 6D B8 72 E9 CA 2F 3E C4 14
 0C FC 28 0A 29 9C C7 94 4E 87 58 12 4B 0B CB 9E
 81 05 F0 D3 01 BA 3C 93 5A CC 72 EC 1A F9 FF 04
 49 98 C2 3A 80 70 34 B7 5B 24 05 FA 57 EF 93 A0
 E1 DC AD A2 FB 71 04 AA 0C 83 E2 B5 08 B5 B3 5A
 01 18 B9 11 0B 9E E8 C1 ED 06 87 32 65 25 7B B3
 77 5E 3D 29 50 C2 E7 83 1D 7C D9 60 00 28 63 05
 B4 95 7F 76 00 38 66 45 78 43 79 FA 8F 52 51 14
 C4 E2 76 4B 87 7C 27 A2 DE 49 DE A5 CC BD 86 2F
 5A 7C DE 19 6C A2 67 20 E3 43 F8 0D 62 4A B7 49
 56 D0 B1 98 5B C8 D5 93 69 41 1F 01 87 E5 86 85
 DB EB 22 8C F2 AE B9 FC 82 E7 92 D9 9B FE F1 55
 F9 5E 0D 24 4C 4D 75 36 CB 4F 9D 6C 1B 2C 8E AF
 B5 88 C4 38 B3 D1 83 75 A7 B1 B1 D7 80 E1 C5 FB
 37 E0 3D A3 BE F7 B5 84 72 43 40 BC AE 2C 5C 1B
 53 16 2A 08 B8 61 C0 00 D3 39 CB 61 15 A6 9B 24
 31 D1 8D 6E 3F CC F4 70 02 C1 CD A5 C5 D9 E4 2C
 F3 50 E4 AC BA DE 61 09 7E 8C 57 B3 C0 BD 9D 10
 49 3E 41 F1 CF 04 FB F1 3A B7 3E CF 67 37 B1 8A
 88 0D 41 6D 39 B8 EF 92 44 59 EE 05 6A A2 72 B6
 CA C8 AB DE 79 B4 2B EF 2B 6F 7B 2C DE 5E 78 AA
 07 B9 DD 95 4D B6 50 09 DA 58 D7 2C B9 3F 40 15
 DF 54 F6 1F C8 CA 8A 89 05 49 21 78 20 6E 1C 56
 57 14 13 5F AA 8E 54 89 1A 9F 68 04 E2 ED DF 22
 13 84 08 66 6D AD 24 BF 5A 6D FF 80 7A F1 15 A2
 CE 2B 16 28 AD 4B 18 70 0F DE E0 2B CE 53 97 60
 D3 1D 7B 9B E2 8F 19 81 F5 26 7F 5F C4 28 7A 43
 79 1A EF E0 0F AC 97 1D 24 4F 6E 91 54 02 56 5D
 19 A9 54 01 F1 EB 2C C9 46 2E 11 28 B3 99 1B A8
 5D 53 94 52 6B 40 B0 D3 00 AF 90 17 85 CD 5F A8
 F4 1C 34 E8 B3 8A F6 36 75 65 E6 C4 34 96 42 44
 7A 21 62 28 CB 36 49 7B 60 37 4B CD 4B 18 82 39
 EF 49 DC F8 61 48 5D 33 E8 08 D1 50 6F 19 4C 65
 71 A5 F6 BC 5F 7B CB 4C 55 39 7F 8F 7E 1F A1 6B
 FD E9 AC 25 E0 A8 CF 83 B0 97 59 FA A8 32 8C 5D
 6F 28 B7 58 FB A6 02 27 1A 4F 05 6A E4 F0 81 F6
 46 E4 AD BC 95 93 1B 69 11 6D E1 E0 D1 38 CE A2
 B8 BE 86 11 B7 0A CE E2 4D 7E FA 9E D3 D7 D6 F1
 88 AB E2 52 8F 2C E7 9B 24 A8 63 F0 49 C0 6A F4
 0D 5A D1 06 B4 44 A2 34 B9 70 A6 EE 61 7E 62 6A
 C0 F6 55 88 F6 56 CC 72 B2 5A 23 D3 93 59 CB 96
 15 E0 42 34 DA AC F6 61 A6 12 C9 E9 DD 67 84 5E
 26 F8 13 36 00 DB AE 5C 0C 4E 52 C1 95 6A 47 D5
 67 C7 7C 5E 5D DE 9E 1C 6C F7 34 C3 D0 27 A5 7A
 05 3E 26 00 CC 11 86 1B D6 8B FD FE FC 17 3B BB
 61 22 B0 09 51 DF 3D 87 BA 48 47 93 AD FF 38 56
 B3 70 BC AE 75 BF 81 3C BE D1 EF 5E CF 6C 38 7A
 1E 4F DC 4D B0 CE 40 6D 6B 92 96 B6 98 A2 51 7C
 29 D5 96 4E 45 DB AE 2E 18 87 5F 37 C8 0F D5 71
 D6 09 8F 51 64 7B 63 ED B0 D3 DF 26 97 34 F4 1F
 BE CF 81 0E 85 58 F5 7D C0 8C A6 FF C8 EE 49 F2
 A1 66 A2 B9 CE 80 8A FD 5B 27 28 F7 06 9E 37 44
 17 2C 1E 34 7F 41 93 E3 1D BA A8 D0 D8 F3 74 99
 DC 83 4F 80 8E C8 85 9E 0B 92 C0 02 0E B8 09 6D
 0E F5 28 70 DB 93 20 19 5B F6 45 9A 6E 9A F2 6E
 4D 69 45 FC 8A E5 31 96 F7 9E 03 C6 02 B6 BA 68
 C4 11 37 4B A8 68 61 DD 2A 6F B2 BC 36 54 62 47
 C8 63 D5 13 25 22 3A 08 76 CE 63 5A 1C A8 D1 A3
 B8 34 6C 0C 0B 08 F0 F2 DE F9 78 3A 9A 6F 6F 32
 E1 01 C6 45 C6 A4 C5 30 BA 19 9D FE 28 8A DE 29
 0A 90 E8 43 D1 B7 BF CA 28 38 C9 A3 7F AB 95 1B
 8E 47 52 53 01 7B 5A 98 AE 39 46 79 B8 3B 7C FF
 63 15 C3 CA 2E 12 0C 08 B7 67 29 74 34 3E F8 4C
 DD 0F 76 3F B6 B6 62 D9 D7 40 B5 E9 74 72 7D 73
 57 7B CE 3F 1E 96 98 99 E2 45 20 3A 44 6B A3 29
 E1 AD B0 4E C7 1B 0A 51 A4 2E 2F E1 FB CC 23 5B
 39 B6 AC B0 4F 58 34 1C 24 B6 FC 17 65 38 A6 57
 84 C9 8C 9E 7F D3 B6 96 1F 6E EF E1 56 63 60 62
 F8 DE 5D 09 5B 00 66 13 25 06 D7 2D EE 2A 71 C3
 C7 66 1E 18 CA 4E 6C 23 B0 6D 40 C6 75 4B 0B C4
 2D 7D FA B8 3F B0 4C 49 DB DC 1C F6 04 BA 94 10
 FF 6F 64 74 B2 A0 5C 62 A7 70 AF FD 88 06 B2 A1
 0C 8D 0B A1 0B 72 98 97 AB 1F 18 A4 DA 5B 99 B3
 C5 77 8B 88 3F 99 8D C2 1B CE 05 DE E6 20 90 14
 D0 ED D9 54 D0 6A AF E1 7F 6D 8D 2D BB CC F4 BB
 A7 2F 80 38 D4 AF 7F 8A 78 63 35 0C C9 D1 2D DD
 72 F0 69 F5 8F 8D 07 0C B6 A0 DA 9E ED 98 B7 E1
 34 47 AB 59 F9 49 40 08 75 A0 45 1A B2 8F 1D E5
 96 F7 64 4F 8B F9 BB A9 55 D9 3D C9 D6 45 88 DB
 1C 9C E7 69 31 8D B9 F0 3A 4B B9 DE 54 CE 87 14
 70 FE 15 B3 9C 84 3A 4E DF C6 6F 26 79 60 BE 66
 E6 01 5E 59 48 9F 89 34 BE F8 B2 AA 85 3D 31 A4
 5F 58 24 A6 68 EE FE 15 49 CD 8D 6B ED F4 1C C4
 2F A9 CE 0A 4B CA 6F A2 91 BA 93 B8 03 AE 7D E7
 9C 00 18 03 43 EA 01 B9 EB F2 40 0D 6D 51 80 A2
 42 70 6E 5D 9A 4D 52 97 B7 53 41 02 7F 67 BF 6C
 E9 CD DB B6 1C 8C 0F 7D 78 D9 0E 08 27 DB D7 F1
 BF 31 C3 FF A2 E2 BE DC 03 13 39 79 14 C3 FE C9
 00 C0 19 6F 74 19 77 AF 94 95 DB CD 35 EF B1 37
 EF 47 2E 9C F5 C0 05 C5 8F E0 FD CE E2 BA 19 D1
 08 A3 6A 31 F1 6C 68 54 27 A7 93 5C 29 B6 2C 49
 D1 0E F6 FA 0A A5 F8 66 6A 3E 92 FF 33 FB 7B B0
 0C B6 96 56 85 AC DE 69 5E 86 77 23 58 11 24 45
 91 40 F3 11 D5 D2 24 BB FF 05 3D 37 5B 92 95 31
 AE 28 DF 92 B2 8D 30 A2 0A E3 FD 49 E3 96 61 41
 19 AF 26 6C BF EA 3E EE B6 FB 8C E4 CF EA 24 33
 EF 64 A8 98 75 69 BC 1C 16 9A 99 56 F6 D5 35 F6
 F3 71 06 C1 2C 78 B3 F5 1B 29 87 45 92 0D 0C 59
 3D 26 76 B5 47 1A 7C E8 E2 F1 F9 44 6E 85 A0 DA
 0D 41 48 A0 89 17 D4 D5 6C 6A 20 7E AD 30 17 12
 C9 2B 6E E1 D1 DB 3B B8 DB 9E B2 92 3D E5 83 8E
 4D 8C 3B 95 E4 EC 6C E5 6C 7D 0D 07 D6 B1 42 75
 C8 9D E4 BC 1F 82 0D 76 FB 02 3A 65 C7 78 D4 B6
 3E AB ED DA D6 A5 AB 9D 26 5E C9 64 F3 70 9D 79
 DA EE 04 75 44 A9 6B 7B E7 10 CE 0C D5 5A F6 C3
 BD 85 0F FC CC 36 27 08 0F 1A 6F 3B B5 2E 9E 5C
 DC 3D 1B 33 C3 B5 DE A9 03 D1 0A 78 40 9C 04 AB
 6B 7C 83 F1 47 08 45 A3 48 DD B4 53 33 BC 34 0B
 9C F4 4B 59 9B 11 3E F5 22 EB AD 36 B0 41 B7 D7
 97 B6 F0 DE CC AB AA 6A 8B 53 A5 D6 0B BC E4 47
 98 FA 90 8B 9E AC 3B 10 46 5E E0 D3 42 78 D3 A0
 D7 32 60 E0 C7 24 EB 2C B6 29 4F AB 1C 96 6E CD
 7E BD 3F 02 59 31 BF 46 44 BD A1 65 64 D9 37 83
 12 E9 01 E4 2D BF F0 8B 8E A4 CB 0B 18 8F E1 FD
 DF D7 F3 03 8A 63 66 07 AF E4 12 38 E7 55 AA EC
 7B 5B 2E 5F FA C9 C9 78 A4 DD 60 DC 99 46 9B 4F
 45 D7 B3 80 A4 1B 2B 49 FB 23 F9 D7 F7 04 9F 4B
 53 45 15 33 16 41 F2 41 D7 E3 86 22 D4 62 BC 19
 D3 36 FA 04 67 54 D4 5A A1 5C 85 37 93 E4 28 2E
 B5 E4 D3 35 EB D2 E6 3D 82 02 74 F9 1E 1B 70 7E
 3F 5B B5 58 47 1C 4E 33 32 35 ED 06 98 35 98 A9
 8D E8 99 2F 5A D9 95 75 28 0C 3B 58 E2 D6 F6 CA
 FC 50 A8 0A BD DB C7 AC 83 A6 A6 BC 8F 74 36 D4
 AF 4D 70 39 58 53 7C 55 49 36 14 F1 94 5C 38 28
 2E 45 9D FF 89 DB 81 91 C7 04 37 C1 FF A7 E5 87
 91 3B 76 42 CB 36 12 95 82 1F 24 96 8A 43 E2 F7
 45 57 72 67 0F 69 D1 AD 37 91 F8 C7 2A 2E C2 B7
 3C 35 50 2C C0 AE 63 29 D8 D7 07 DE 40 5E 2B FC
 72 F9 BD E3 0E AE AD 66 DC FF 4E 11 AE 3B B2 F5
 1D 6E 73 8A D2 96 48 3B C8 44 51 73 1F B7 7E DE
 7C E2 34 B6 27 5C 24 6C B6 EC 1D B7 D3 BC 7E 22
 04 A2 B1 FD 6E 7C 36 74 F8 07 A1 0C 82 6E EB A5
 48 AB AF 6C 94 6D 6D E0 5C 27 3A 72 BA 23 19 60
 55 4F 7F 58 39 5E EC 91 41 D8 E8 16 15 AF 0D 6D
 88 99 7E 52 25 DA B6 E0 72 45 ED 59 17 92 6F 2F
 11 8E 83 E0 65 98 8A 87 4C 2E AC 01 57 12 98 C3
 42 AF B9 EA 90 B4 1C 92 89 19 CF 7B B1 E4 B1 76
 DE F6 69 23 32 88 0C E6 48 8A 43 56 17 C6 8B C2
 CB 9B 00 B3 07 E2 F9 C9 53 C7 D3 28 66 DB 77 1A
 51 93 1E C5 50 37 35 F8 90 1C CF 69 26 D7 00 9E
 70 10 76 97 B4 E3 1C 1A 17 09 08 32 A1 27 CB 49
 C9 EB 3D 83 02 49 D3 12 18 29 22 4D 76 ED 17 00
 81 2C 70 60 A5 57 A0 B0 51 4F AE E6 3F 34 98 08
 B8 C0 71 32 91 8C 21 DD 15 D5 7B FD 5F 5A D5 ED
 14 A2 94 FB F3 10 2E EB 55 A0 83 42 6A 42 1B 71
 E0 A5 B2 DA 6D 75 0B 5E 26 37 9F 38 97 48 AF FC
 18 09 02 25 03 64 6A A1 D5 13 1D BB 88 1F 6A BB
 43 CD 19 0D 83 E7 25 86 40 3B 74 5B 9C 3D A4 B8
 C9 75 29 34 06 E4 BD 48 6B FE ED 35 7C E3 40 A4
 5D 4D A4 6F 1E D0 95 FC 85 7B FB B5 54 4E AD 26
 DF E0 41 1D 74 28 DF 50 9B 79 E5 FA CA CA 8F 07
 55 95 F6 A7 EB 68 F7 2A 57 FC 4E BD B9 D1 FD 49
 0D 88 84 53 5D 8B 9B FA 45 26 0B 08 15 3E D0 03
 C0 B5 45 03 1C 68 E0 E5 58 97 1F D4 84 FA 1C 82
 3E 1C 83 AF BA 5E B0 FD 02 07 C5 C9 FA 4D F9 EC
 D4 2E 2B B1 73 4B F9 10 BE FB E2 69 43 83 AB F1
 BF FB 66 EA 9E DE 45 CA 05 14 E4 DD DB 4D 47 4C
 B5 C1 7F E9 15 9D D3 94 C5 AA 8D 02 8F 01 84 51
 C0 D8 38 EE 64 56 35 D5 24 2F 84 A4 B8 78 1A 5E
 76 78 CD AD BE 51 65 FC 4D D8 9A B7 26 47 45 DD
 B0 70 EF 08 09 E2 66 71 30 C9 0E 2A EB 8D C1 E7
 50 BE 6B AC 8C FD 43 94 85 F9 47 DB 28 3E 62 87
 0F 1E 3F 0E 78 E9 62 1E FA BB D8 71 4C 01 61 34
 63 24 16 06 FF 6A A2 0A 2B 9E 60 74 B1 99 B9 95
 F5 E0 FD 1F 0A 43 9B F3 13 FA 11 8F C4 BC D2 97
 4E F2 48 D8 6C 70 0C A4 7C 45 BF 6E A2 F1 37 75
 83 0D 7E 0E 02 4E C9 66 7B 88 DB E4 64 26 84 8F
 76 D6 90 1C 74 6D BD 39 57 54 14 B2 AF 2E AF 24
 08 FB 6D 1A EF 5B AD 1C 58 B2 1A D5 33 AF 74 E8
 CE 10 FF 54 16 D5 2B B1 05 5E CB 9B 8C 5F 0F 7A
 A2 78 A2 D4 28 45 FB AB 61 BF 58 CE 1D 75 48 7D
 1B 0B 7D D4 AB 32 BE 43 DD C2 9B 6D 52 0F 03 92
 05 93 12 C4 34 FC 13 61 4D 99 96 20 26 23 37 E5
 0F 7B 51 8A A7 E2 DF 36 FB 68 7E 1F 46 54 EC AC
 53 B5 2B A2 47 C0 CF 5B 19 D8 3C 40 4C 7E D8 75
 3F C7 5D A5 10 49 B6 77 07 49 10 38 D5 92 F6 02
 AF 48 11 08 F0 3A 4C 75 3C FB 55 4F 59 CA 72 C5
 E3 D2 31 3A B6 47 FE 66 FB 74 4E DC DE FC 67 EA
 9D 94 BA A9 4C B3 D8 C9 2E 20 24 7D F9 4D 4F AA
 A7 5D 9A 76 76 8D E9 17 01 86 9B 71 53 15 0C 6B
 D9 E2 15 ED 72 A5 11 39 82 80 5D B3 F3 2E 82 85
 A3 F4 4D C7 F2 97 54 C6 01 2C 92 0B 5E 28 44 6F
 98 18 82 E7 02 85 07 AA 92 E0 A8 33 29 09 66 BE
 6E 75 94 45 6A A4 F1 72 BC 32 AB E0 21 3D 6D 77
 50 A2 EE 59 33 5A 63 D5 19 12 9D EC 92 C5 5F DD
 BB 4D F0 27 0E 0A 7C AD 98 FB A9 83 CD 31 DA C4
 19 8F 6C 95 27 85 B0 30 0F E2 68 C8 91 E0 23 CA
 BC F4 8B 4E 65 0A A8 CD CA A4 65 55 CE 8F 27 3F
 7B 80 D8 2E 3F 88 06 B8 FA A6 9A 55 FB 51 CF 59
 CD 0C 1C F5 DD E7 47 F0 35 33 AB 2C 57 49 35 AE
 40 D8 8E C9 82 0A 4D 61 DE E1 43 9D 52 CE 21 AC
 FE 6A 3A 6B 45 58 C8 EB 93 E4 DC 85 47 DC 68 C4
 37 AE C7 1E AE A5 31 EC D9 9A 44 94 A1 66 5B 15
 D6 C5 FB E8 DD CB F6 10 BB 85 46 8B 35 0E F6 65
 A7 F6 31 25 E0 33 F2 CF 1A 68 09 86 BD 24 46 58
 C3 6C 62 5C 02 1F 40 46 5D F2 87 C4 D3 43 F8 C1
 B8 95 80 DC 46 3D 34 E9 A5 CB B0 F1 F2 5E B4 D5
 80 C9 2A 2E C5 FC 81 3B 3E B9 FC A2 39 45 09 5C
 1C 4A 8F BD 50 ED B2 30 F0 BA 5C DF A0 45 A0 74
 B9 8F E5 87 16 44 CB E1 AC B8 5D 66 5A 3E 61 8F
 88 70 4C 9E CA 36 E8 23 57 5E DE FC E1 D7 A3 A9
 8D C9 E3 16 64 B3 14 47 49 53 FE 61 F8 B0 81 78
 17 C3 92 2C 9E BF AD 57 70 DD EC E0 2A BA 80 C2
 3B DA A4 59 9D E8 7D D6 9B 3D 3F 7D 8C A7 5B 53
 C5 88 9E B2 3E FB EA 35 FC 42 DD E2 4C 4D 0E 19
 4D 1A EB 57 DB 65 2D 37 76 B4 E6 3F A7 45 1A 9C
 3D 11 3B D4 4D AB 5B A8 21 AC C6 22 AF 12 D4 08
 36 D6 80 D9 FA 68 13 AC B2 B6 46 0C C9 7C 6F BE
 B7 FD A8 26 7E 65 8D E1 36 78 F5 0F 3A 01 EC 73
 8E 10 67 B9 F8 26 3B AA EE 98 25 75 1A 27 0A F8
 F2 2C 0F 66 8D 3A 8A F6 05 B9 B7 DD 54 56 DD F6
 48 20 FA 3E CF AA C7 45 79 78 B4 B4 50 68 DD F7
 72 9C 97 98 B0 65 E9 54 5A 2D 69 85 B5 81 7E 38
 9A C1 8C 0F 8F D5 EB BB C1 92 56 D0 61 6D A1 E4
 2C A6 07 77 73 5E D7 10 A3 A2 1F 97 7E 6E 83 D3
 17 87 E4 89 32 23 31 EB DD EC E7 50 5F AC EB 6C
 DA BF B9 9C A5 4D 61 98 A5 ED 4C 42 95 6A D6 05
 62 0C 7C 94 CD 8C 9D DA 65 9D 33 FF AC DA 21 96
 63 EB 71 01 9B 48 3B A6 A6 7D 8F 76 FC 51 31 22
 88 CA 42 63 6C C3 F3 DE 3C D2 E6 7F C7 6E F6 F4
 64 FE 69 9E C2 FA 12 38 42 74 B2 80 34 59 DD 2F
 CD C5 E8 34 DD 49 11 38 36 55 A0 4E 0A 23 A0 3D
 3E 14 38 64 C2 F3 A1 36 0F 6E 48 75 B5 ED 48 8C
 A0 58 D2 01 6B 8B 20 A9 6A 43 45 42 45 D0 F8 54
 34 DD F8 6C F7 5F 39 59 24 EC 5E 36 58 94 B4 A0
 B0 2B BD BD D5 5E F9 F5 48 25 9A 9B 3E CD 19 1F
 2F CB 3C D4 66 73 0E FE 8E 97 62 BC 61 43 AA DE
 CA 31 1C A7 B2 2C 5C B3 2C FD D6 27 1D 5C 7C D9
 38 CB E5 14 70 42 6B 21 9D 11 59 CD 6E 48 E6 08
 82 5B 34 81 D2 A7 3C 45 6D 80 92 4C 5F FB CF 7E
 73 37 31 89 66 2F 37 67 42 51 FE 48 3B 1B 7A DA
 F8 7A 46 EE EA FE 02 2A C3 5D E2 B7 2A 7E 90 3F
 16 90 02 9B FB 8D F8 E2 30 FB 8B DF EA E2 86 7F
 D7 1A 8C 29 5A 04 E8 94 AD 5B 19 C2 92 F8 37 C0
 43 76 09 74 E1 FA 00 E0 67 81 73 FE B3 74 2E C2
 F1 73 B0 A3 8A E5 96 AC 8F A3 8D 9B 65 75 79 4F
 55 C4 DB CE AF AC CA E2 7B 79 9E 02 CF E0 F4 BB
 97 70 FC F8 08 A1 E8 44 08 7B 1D 6F 08 AC 9B CE
 12 B4 F4 8C C8 59 A5 8B 3D 19 49 DA B0 77 D1 C3
 FC 75 A0 1F 97 01 C1 65 16 43 53 91 FD C8 CF 81
 FB 3A 1B 6D AF AA 66 CB 70 DE 2D AC 78 D7 E3 46
 68 DB CF BE F5 53 23 C6 B8 23 9F 18 6E 28 FA DA
 76 F3 B0 83 26 0B 2F B3 3F F1 D9 71 A9 84 31 84
 E8 81 53 3B C2 4C E2 09 82 9B 36 2E C1 9C CF 44
 0A 3A 31 CE 2F 50 D9 14 80 C0 AE 2B 5C DF 9D DD
 16 CF 4E 58 75 17 8A 84 E1 6C AD 98 34 2F 52 FE
 78 A3 14 BC FC 35 91 6C 9A 19 39 47 BF 40 D6 D4
 49 44 A0 DA 58 76 42 BB CF C0 1F 76 AD 50 24 42
 57 AF 8B 90 DF 56 27 2F 62 F7 F1 1D 98 12 C8 F5
 8C 14 D6 8D 07 C1 82 88 A4 37 21 0D A8 45 9E AB
 E9 D6 C6 5D C2 A7 D7 CB 47 93 AD 70 8B A2 AA 28
 DB 5D 0F 32 7A 0D 28 48 F1 C4 FF 3E 8A 71 97 FA
 AD ED 5C 9C 64 73 D8 22 4B B7 72 DB 56 85 FA A6
 6C 47 A0 8A E5 D1 B2 7C DC 78 C4 D9 6B BA 80 6F
 96 3F 7E E5 0F CF B8 90 C4 D5 FC 9E CC 1E 77 53
 2D B8 CD AD 04 40 A7 B2 98 AF 5D 20 79 70 73 53
 BE 1C 4E 83 06 F3 E5 3E F9 86 C6 B3 88 24 74 14
 C2 2A F7 AF CA 13 71 3E CC F3 D5 4B 07 AF 2D 7B
 F4 85 CD D2 04 BA 38 7A 67 0E BD 58 DF 25 29 E5
 6D 9A B1 8C C9 B1 18 A5 6B A8 C3 08 7F 38 20 6E
 00 DA B8 4F E0 3A C5 DE F4 6F 3A 1A E5 72 52 24
 4D 8E 8B E8 F4 EA 47 3E D8 09 84 9A DC E9 15 79
 EC A4 A9 D6 98 BC 39 1F BB 14 A9 2B 83 AB 97 13
 39 C2 10 08 FE 74 A3 7A A5 16 BE 8E 26 71 FE C8
 0A 1F D8 4D D7 43 B8 4B 99 ED 10 EE CD 6F F4 76
 44 B2 57 72 4B 38 AC CC D3 B6 71 59 82 E4 E5 B0
 BF 97 8E 15 8D D3 00 58 D1 62 7B 5F 79 DF 3B 60
 38 4E C4 6A 05 8A B2 A7 87 91 98 32 0D 99 8A 8A
 ED 01 63 85 B8 8F F6 51 91 2E 9C 41 4B 07 74 28
 BF B6 30 E7 C6 8A 1D E2 EE 7F 3D 19 11 93 6E 4C
 04 79 0C 87 C7 B7 B3 79 09 A8 F0 CE BA 6D AB FB
 A1 13 30 72 C1 95 93 0F BF 55 6E 2C 4C 2D 3C 79
 EC D4 EA 9B AF F6 91 8A 40 AE 50 12 C0 CB A6 09
 EC A9 0D 63 AE 1D E0 57 42 26 EB 0F 1D FF BD 0E
 22 18 11 66 AA AE 54 C7 87 C9 A4 10 28 80 C0 B7
 6D 3E 63 E9 E2 7B D1 01 B2 AA B5 BD 61 44 E4 BC
 06 13 F4 38 82 28 9B D3 39 5C C8 AA 75 59 4A A0
 95 96 CD D2 C9 4F 75 08 F2 31 F1 8C 9E 7E 3C 2B
 7B 33 BD 86 85 3D 3B FE 44 FF 01 26 63 D5 0D C5
 B5 0B A7 59 D2 24 4F ED AD 1E C6 B6 20 6F 7F 4B
 E3 9F 14 9B 6C DA 06 E2 D8 AB 9D 0A 2B 7A 26 E1
 95 3D 51 9A 75 F9 1E 93 28 53 52 00 DC FC DF 07
 FF 8F BD 24 28 46 24 F1 B2 FA A3 D8 C8 CF C6 8B
 63 6D 8D 94 29 AC 22 D6 75 F9 56 B3 C6 2C DD B3
 F4 92 74 31 D2 4A 7D 20 74 9C 36 F8 A5 40 A7 3C
 40 72 63 C0 99 56 BB 43 B4 BD 54 1F 2F 30 DD AB
 77 F7 B4 67 1F 4A 02 59 54 00 1F A3 48 CE 2B 03
 09 34 40 5A 9B C8 1D 1F F2 8E 3B 08 8B 5F 1C 27
 95 1E FD AE C5 2D 90 72 C4 82 34 F3 B0 F5 FD D8
 6F 4C D9 FB E3 01 51 A6 60 60 6D 50 65 0B 0A F4
 33 F6 6E 29 D3 95 3A 8A F6 EF E8 5D 97 96 58 E8
 69 98 FE 19 49 38 AB 46 47 99 A8 B1 35 86 30 4D
 C6 B1 74 A1 23 75 C5 A4 A5 0F 22 08 9B 6E 2B 0C
 E2 F5 EA 98 40 60 E3 A6 78 38 BA 2C C6 91 A9 77
 4D 8F C5 A3 04 8C A5 06 F8 31 31 B3 FE 27 CB 35
 3E C3 61 8F 38 BA 9C B7 44 C9 28 51 F2 22 07 49
 8E 5C B8 C7 55 06 14 98 83 C2 24 E9 CC 00 67 D4
 5F 2B 79 72 16 5C 4E BC F1 2E F5 7B 3D 41 26 DA
 D6 C4 E9 C9 F5 41 FB BE 2C 27 A5 0F F9 D4 19 F6
 1A 7B 76 71 CF AD BF C1 70 8F B5 0C 06 E3 48 5C
 3E F7 BB A1 0F B8 E4 FE F2 00 EF 8A ED E5 6E 6C
 DE 1A 76 EC FD 2D 37 88 15 1D 55 61 5D E5 2D 0C
 C7 FA DF 3F 39 20 91 5E FA C8 B6 3F B9 E6 EF 4A
 D6 D1 FB A9 C8 0B 29 48 EB 2D 55 51 88 B8 ED 2E
 28 F9 F9 BC 37 B7 55 50 A9 AD 27 1D A3 3B 17 97
 96 40 63 DB 7E 98 31 FA B2 77 86 BD FE 6D EC 59
 CF 2C A9 12 89 9B 43 91 BD 69 2E 9E 1D 09 7D 5D
 93 61 E3 1D 36 40 BE A7 63 9C 8F 5B AF 2D 67 E6
 F7 A5 4F 34 7F A9 13 35 AE F5 3B 86 CF D0 5B 16
 7D 09 6B 31 80 74 0E 69 99 A6 23 AB C8 FE B4 51
 E6 BD CE 4F 3B B3 23 7C 6E 6E 3B DF 08 79 29 E9
 42 52 7A A1 F8 88 05 DB DB 83 CE C1 31 A4 7D 9E
 C7 E1 D5 9D 0D BA 0A 90 FD 9B 7A CC 92 21 BF 92
 EA B9 45 00 F4 35 EB C2 19 4C F5 81 F0 23 02 3F
 68 B0 A9 60 35 83 41 6D 23 34 53 F8 4B 57 D6 56
 44 79 7B 64 90 D0 00 B1 20 D4 81 D0 FF CD 46 90
 D0 6A 14 55 9A AE 2E 03 30 32 8D AA 17 1B F6 CF
 BD E5 EE B1 B3 F7 CE 71 49 EA B8 A2 7C 37 26 E3
 AB 9E 17 7B FC CD 25 8A 6B FD 58 D0 E6 89 DD 1B
 2B 0A 12 CB 49 51 48 5B 4E 67 92 75 B7 41 2C 35
 A2 AF 4F AC 07 78 B1 8E 6F A7 F6 1F BC 15 C5 B0
 34 6F 95 33 D7 46 8D 19 E4 A3 2C B1 B7 82 44 AC
 37 DA 34 86 17 1F 2F 59 37 0C 6A 2A 8D 64 D4 DF
 30 F0 F9 0A 79 7A 16 BE 43 1C 67 86 EC 66 2A F8
 D1 96 F2 57 72 FD 84 82 FB 06 70 A6 91 B9 01 1B
 C0 5C BA 69 8D 3A FB 5A 2D CC 35 19 44 7F 2B 17
 10 4E BE F2 53 9C F2 25 F7 CD 3A 86 68 8E AF A7
 66 15 3F 16 21 12 64 1E 88 C2 CB 10 0C 98 49 E8
 EE 38 02 DE 0B 15 EF BA 6F 5D 08 F4 AF 76 98 35
 6E 83 44 83 C8 C1 64 65 10 75 67 4E 3D 9B 86 7E
 F0 68 D5 B5 45 B8 8A F0 71 09 86 59 AE BD E8 0F
 82 DF D5 45 0E 16 F8 C0 AF 32 35 63 7B FA C0 00
 11 BE 2D DA 1A 17 93 37 6C 32 0E 80 E6 92 38 10
 8B 65 65 92 A3 54 AA 36 D0 58 E1 F8 7A E4 48 A0
 9F 52 5C 90 B7 D3 CA F7 1B 40 DB 97 BF 87 19 1D
 84 D3 15 B1 40 EC 48 5A 53 1B F6 78 67 1D 77 DC
 39 A0 BA E4 42 93 A9 53 78 6C 9C 51 0B A0 15 71
 65 1F 6B A8 2B 6E 4D 4C 42 E9 3B 49 83 47 8F C0
 3C 1C 56 19 B5 A7 6B EA BE 4F 64 15 49 6F B8 4B
 7D DD E1 8D 24 4E FB 64 C2 3F 15 42 A6 5C 7F 33
 37 6B 8A F8 89 52 79 0D F9 12 AE 9A 2C D7 71 E2
 B6 B1 02 74 C8 03 BA F5 98 DD EC 1B C0 AF 86 2B
 D0 F5 5E 56 2F 75 19 19 67 18 B4 66 7A E1 DF 6A
 EF 16 4B CA 0A 73 4C 83 B5 4A B2 E7 3D 43 FC DA
 12 E0 5E B0 0E 9E 2A 11 B9 80 94 20 D8 C9 D4 1B
 95 1E 60 4E AB B0 13 BB 0C B9 13 44 C9 C7 89 91
 19 06 06 7B 3F 63 EE CA 7E 69 70 AD 21 E0 37 27
 7C 6E 96 DD 69 2A 84 CD 94 B7 25 BF 78 AB 76 FC
 60 9D 10 2E 15 2D 65 65 AB A0 32 16 E0 2D CA AE
 D6 6E 0F 56 2F 4E DF 4F 43 4F BA 61 74 8E FC 01
 3F B5 FB 6C B9 53 3D 38 C0 BE F4 DC F4 F2 65 BA
 67 53 2C 8D 36 CA F7 B5 77 07 25 68 2A A6 09 D2
 D3 D9 FF 0F F6 1E 08 3C BC 06 36 6F 2C 7B 38 7B
 C7 6E 60 F1 40 F6 D6 27 11 E8 3F 6A 3B CD 9F 1A
 EB 3C A9 FC 9A 38 E9 B3 E3 45 43 34 D9 94 1C CC
 95 EA 76 DB C8 F6 9A 76 2B F9 0D 38 DB 81 08 BB
 23 A6 08 09 8D DB 80 FF 27 33 60 85 1A 73 E9 F2
 A6 1C 14 6D 05 79 93 59 6C BD 26 23 79 93 5F A7
 22 83 A3 FA 7B 21 45 BD 68 61 9E 84 A7 EF BB 16
 25 04 5A 2F 1C 2B 46 3E 47 C2 58 57 51 EB E6 51
 73 85 90 9D 5A 74 5E C9 F4 B8 59 34 4F 6B C6 0E
 DE BC 63 F7 C3 DC 42 01 74 CF 66 AD 4F 0F 18 A9
 A9 EC F9 76 3F C8 ED 62 DB E7 DB 14 68 9C 23 83
 3C F6 57 45 8B EF C4 32 C0 61 E8 EA 08 4E 46 0F
 79 3D F8 D2 94 0A 09 9F F6 F9 47 6B 7F 33 B8 90
 A9 80 BC 4D 91 FC 6B 0B 6B BD 84 C7 EE A6 99 6E
 2C DD A2 29 27 89 26 0B 20 8D F6 8B 65 F8 83 86
 4F 01 F9 FE 0B 3E 4D A0 C2 90 06 94 5F 7A 9C CE
 53 FA 65 0C 9F F5 2D 1A 82 4D AE 08 4C F5 71 B6
 11 10 4B 6F F4 CB 0C 52 4B B7 C7 08 BA 43 9F BF
 4E B6 34 0D CD 86 67 00 04 F3 6A 90 9B 86 FF 26
 6E 6E 9A 00 DE 8D 0A 92 2D D4 7A 55 79 1A 00 AD
 90 E7 ED 08 29 AF 15 FD E0 AE A3 0C E3 CD E7 A8
 E7 55 C6 30 9A 66 A0 00 B3 CC 9F B4 3D FF 8E 39
 35 0E 1B 99 2D ED FC B9 D9 94 B5 D1 7F C5 B2 4B
 0B 62 98 3F 06 23 2A CF 60 C7 D9 93 9F F0 BA CC
 0B A8 4F B7 BE 7F A2 84 2F 50 AF D1 65 0B CF 87
 5B B8 7D D1 DB 01 0A 83 86 38 9A 17 2B 15 C1 8F
 D6 E7 20 DF 89 19 2B 0D A0 97 CA C2 FA F8 CB 29
 45 DD 44 53 06 A2 9D C3 78 E4 70 49 0C 75 BE 0D
 74 F5 CF 71 7E 94 F4 96 E7 6F 3B 28 63 25 BF 75
 9D F6 DC AD B0 24 80 94 2E 86 3E 8D EA 39 D3 46
 E4 06 91 D2 0B 80 9C 2D F4 20 53 93 19 6C FE 6A
 3D 60 77 5C A2 40 04 D1 4A 8F A9 80 F9 02 FB 65
 00 4C A0 B5 8E EF AD 59 0B DF 0B FA 04 56 13 95
 EF 9F 99 7A A8 C3 55 3A F0 86 5B 22 61 D0 D9 4E
 90 DD 35 0B 89 A7 61 42 32 D8 43 74 DC 85 CF 27
 26 CC 61 2B 79 43 8E D4 D1 7E 6B F7 CE 2D 06 5F
 13 D6 4A F9 3A 46 96 57 77 E6 BC E3 92 17 1F 9B
 99 60 48 3A A4 85 86 4E 26 03 F3 25 A5 69 19 F2
 8D 50 96 22 7F 03 A3 D8 03 B6 15 74 93 A7 B5 AC
 FB 29 70 A3 0E 9C 9D 14 E4 A8 7E F7 57 46 90 4D
 77 D1 8C 17 5C C7 55 A3 C3 F2 0A B3 DC 0B BA FF
 0B 2A 32 56 84 C4 31 D8 7F DF 3A 91 2E 92 57 88
 9E 56 16 8D 27 09 D2 55 62 4C 6C BF 8C 75 22 41
 A4 09 63 0F BC 59 1A A9 95 0F 61 01 7F E5 89 7A
 CA 24 74 0C CE 36 6B 2D A5 A0 00 62 A6 99 D4 0B
 29 C4 06 8A A9 34 7C 8E 69 96 88 8D 22 A5 1C 5A
 15 3A 43 34 D6 F8 74 82 02 9F 9B 07 9E C7 D3 57
 31 EA 78 A6 D0 95 8D 3F 29 38 6E 12 E8 2D 63 64
 32 92 EF 5E BC E0 8D D5 57 28 38 AD 14 EE B9 AF
 F0 53 3B 71 71 AD 4D 41 35 DB 52 7D F7 F5 39 4C
 3D 39 34 F9 90 8C 38 3F BE 70 5A 81 99 03 F3 0E
 90 DC B3 32 41 C9 37 64 51 7E 71 38 B5 7F 85 4C
 00 89 63 E6 F0 4B DD 69 DB 77 A1 DD F1 55 2A BA
 13 45 90 6D 01 5A 30 FD 2A 6E 4E 6A B6 D2 35 05
 FD A2 DA F8 13 57 99 4F 86 BB C0 BD D0 93 69 86
 08 D5 82 CA 5E 08 3C AF B6 4D 55 B0 23 61 2A 6E
 48 DA CE 8C 7F C8 AC 98 63 15 67 AC 89 CA B3 BD
 C4 E0 D5 0B 0A 67 92 BD 49 BE 5B 07 79 3B 6C A6
 06 2A 96 51 75 3F 2E 51 ED 7F E1 9F 8C 20 F5 55
 18 E2 08 BE 52 5E 36 55 0A 4C 49 A9 F0 6C 4C 1D
 31 63 E3 CE 69 13 D4 27 0F 08 8E 91 3F 30 0A 02
 93 1B 7C 06 BA 5C 3A D8 B7 CE 4F AB 94 11 57 B6
 2D 1D 3E B9 2D EF 50 58 CB 69 78 83 62 26 BB D9
 57 4C F0 8B 19 CB 73 61 38 08 1C 2D B0 54 B8 AF
 13 CF A8 94 56 BA C9 2E F2 7C 84 B6 B5 91 76 2B
 FD 4B 76 5D 5B 25 62 9C 4F 8C 0A F4 93 44 68 68
 38 80 0F BF FE 27 9A 01 9C 4A EE 75 3A B3 26 30
 6A 24 2B E1 04 82 EE 0C 35 94 00 E0 63 34 64 CC
 73 D7 B3 B1 4A 12 CD 6B 4C 34 5A DA 4E C7 0B 02
 45 C2 B1 95 AE 2E 1A 68 C5 4B 2C 6D 89 23 1C D5
 BA 43 3A 3B FC 04 D0 73 7F 82 4C 22 66 EF B3 E5
 49 BA 10 40 14 D0 36 5E C0 25 FB CE 2A 79 AC D6
 DE BB D9 91 AA 03 26 BB BB D9 29 8D 15 0E 79 ED
 DA 60 2D 94 E9 CB 1F 71 10 EF 00 E5 1F FE 1E B3
 6D 27 7F 69 A1 16 88 DB 2B 7A C2 5E 69 80 DC 70
 90 A4 39 7E E9 82 B4 1F 87 6D 7A 4D 72 80 B9 DF
 D1 16 8B BE DA FF A2 F9 E0 14 A5 F9 69 29 D0 C9
 AC BB 74 B7 F0 18 98 04 B2 1F 85 2C 84 DD 4C F1
 CF 07 20 7F 44 79 4A 13 F7 9A C4 AA 72 88 26 2D
 AA D0 1D 96 96 44 AA E4 07 4C DB EF 81 C0 40 02
 88 1F DE E6 95 FB 8A 93 13 11 D2 CF 45 BE 96 7D
 26 DB 6E A3 DB 96 63 5E CC EC 27 50 7D C7 DD 4B
 58 00 F4 E9 28 41 EA D1 08 B3 17 03 F6 2F CF 8D
 49 43 2F FA 9D 08 DE BC F1 1F B6 8D DD 92 99 B0
 AA 77 A2 9E 64 DE 46 F0 63 2E 14 43 17 88 48 4F
 9D EB 6F 78 5A 35 BE D3 E2 07 F1 6E 93 7D C7 B1
 62 92 67 D3 82 77 55 10 14 2B 1A 11 3B 25 60 E9
 F7 F9 AE C4 82 15 74 83 E7 06 70 8D C0 96 C0 4F
 14 B0 9C 62 66 45 C7 17 D5 70 3B 78 C4 74 6C 74
 D1 37 01 E3 39 F5 3B 34 9E E0 89 19 10 F5 9C F0
 E4 03 18 60 76 4A 37 C7 4F EB 1E B4 30 A1 49 69
 50 9A 14 F1 F1 0D 9E E6 C6 C6 1E 72 69 E3 A2 2F
 92 7C 77 A8 61 E7 0D BE 57 24 B6 42 7D DF A9 E6
 19 14 6D 1A 60 79 5F B4 2B E9 4B 0D ED 8F 2E 9C
 7A DB 93 5E BD F2 1F 09 8D 19 12 92 3A 58 FC BF
 A3 A6 67 6B 9B 33 A4 84 A0 9E FB E1 53 B0 5A D0
 89 8B 37 1E E8 F5 60 0E 63 37 E3 9B 23 88 84 7A
 58 F2 E7 A2 6E 3C 93 2A AA 49 5D B1 C5 64 C2 6F
 B8 67 89 7D A9 B7 8E 61 EC B7 59 A8 2C B4 7C 88
 24 C1 23 90 E9 2F 24 75 34 61 E3 C3 9C 1E 6E 30
 D4 C3 5A DD 1A 7A 32 3F 75 F3 07 A1 C1 FA 39 AA
 00 19 1A 88 11 9A F1 AF FB 2F 0A 1E 2C AD 60 34
 85 A4 AE FE 82 8D 5A A5 54 9B 33 1D 01 42 05 44
 36 A0 66 E7 C9 87 51 3E E9 25 02 4D 46 38 F8 46
 6B 83 7A 42 70 C2 5B 0D B6 8A 62 F2 D1 C1 91 3D
 D1 64 7E BC 60 52 85 51 B5 C1 C0 10 3A 14 30 2A
 56 8E CC B8 CE 21 71 3F AA 01 80 C4 EC 34 9A 1A
 09 FF C5 05 27 37 85 54 7D 74 3C EA C3 A6 FB 2E
 6F EA D5 BC FE E6 6B 59 1C DD 98 C0 EA E7 BE 2F
 F3 81 C8 AE D0 7C 0F E9 E5 7A 45 AC CB 82 51 A6
 B9 AC E5 7F 2C C1 01 92 15 7C 1D 94 8A 74 46 34
 0B EA AE 36 13 03 42 0E 97 7D ED F7 3C DA 83 DE
 96 BA BC 77 DA 31 34 F6 B8 6D 63 E8 8C E1 CE 24
 76 80 DF 91 73 4F C1 F3 A1 62 8B 3F 5B 2D 00 95
 4A 19 1D 74 15 87 11 5B 98 18 93 E3 A3 FA 10 0F
 15 48 7C 14 26 9F 8A 12 9B 45 12 90 09 51 EE 33
 1D 06 EE 05 50 9E 40 41 C6 F0 7B EC 77 33 89 75
 65 A1 1F 43 04 B9 A5 38 AC 56 6C 4F CF FB A5 28
 D9 D0 CE 30 98 B3 26 47 0B E8 C9 01 5E C6 D7 81
 EB B9 FE F6 D0 A1 2E 63 57 E1 AB 1D 6F 95 B4 AA
 29 30 E2 1C 58 7A 8E E8 CC EB 4F E5 7B AC 9B 93
 81 17 17 37 9F C6 47 39 DB 99 E9 ED 3F FC 06 FD
 58 F6 94 E0 C9 AA 3B D8 F7 B5 B3 50 E3 9B 1E 5B
 1C F0 8F C3 E3 4C 41 A9 75 B4 89 D6 98 E3 A0 36
 4E C8 A7 A9 B6 C4 02 FB 37 F0 CC 21 22 AD BF BC
 9F EC 21 40 D3 32 01 97 A4 90 7F 8A 67 41 78 FB
 0E CA 51 3D 96 93 7C EA 86 7D EE 83 6D FF F6 0E
 A3 67 5C A7 7E C2 F6 2E DF 49 6B 3A D8 5B D4 27
 DF D6 53 A8 4E BA 54 15 A8 6A F6 AE 7D 1B B8 84
 6A 3E 81 AE A3 93 27 E5 B6 8B D6 BE E1 37 11 F1
 89 04 3E 76 30 35 A0 DF 29 1B F5 0A B9 D8 F4 B3
 1D 5E FD FE 87 A9 07 E6 11 15 7E 8F B4 D0 BB AF
 E3 85 8F 19 81 5E E3 55 40 10 0C 3E 76 6B C2 36
 74 DB 3C 76 50 46 23 57 50 42 ED 34 A7 86 B1 F6
 E0 90 56 5B 22 DE C7 21 9A E4 72 77 38 56 4E 7E
 C7 B5 6B 4D FC 2A A4 06 50 09 59 A4 12 C2 E3 9B
 54 44 7A 6D 1A FD 8B 52 CF E5 7C B3 58 D7 95 5A
 ED 98 C2 B6 41 BD 3C 6A 8B 92 40 14 26 63 58 53
 3E 51 85 F7 2A 47 93 5F E9 E9 31 46 84 E4 B6 68
 56 2C 6B F1 F9 0F A4 F8 B9 4B B1 06 3B D1 5A 94
 C1 6E 28 D3 67 AF 3A 0B 48 AA A6 98 44 C7 AA 57
 3A C5 57 BF E0 C5 65 DE 06 AD FA 5B 84 FB C9 35
 C1 89 4B 18 84 17 7C B9 48 0D 2D 45 F8 AB 99 D4
 72 45 52 AA 12 55 28 92 32 64 81 CB 6C F5 6D E5
 53 CE 19 54 AB E5 2E AF D8 54 32 25 7D C4 1B 2A
 BB D8 7F 60 97 4E 7F 79 86 85 17 77 0B C8 C2 09
 0F D0 F1 08 96 3A 8F C1 00 B2 32 EA FF 4F 1D 0A
 A7 3F 68 85 B9 20 72 76 4D 55 46 4A 6B 58 94 8F
 8D D9 74 06 DF 0A 46 30 3A 8F 78 F3 14 0C 40 ED
 C7 80 AE D6 69 FD 3C 69 A8 68 CB 3B 4D A0 CE 94
 30 C4 22 63 5F 2E 82 BE 97 E7 C5 24 66 F4 EE 44
 35 AC CD C5 42 68 9F CD E8 E1 A9 8E 64 D2 98 22
 06 7C 86 EF 65 A2 FA 32 82 84 1C 71 87 2D 4F F3
 E5 D0 F4 B7 EA 65 12 C6 DE 70 6D E0 5A D2 6A 68
 5D 1B 35 D0 DB F3 88 B7 D9 A6 E2 B7 A5 26 2C 9C
 4D 65 D8 F3 4C 49 33 33 EE 1A 41 A5 E1 2D 0F C8
 2E E7 38 DB A1 97 D7 6F 66 8E 55 32 57 85 43 E3
 2C 1C 72 28 BC 3C D0 EB AF 7F D5 70 3A 21 F4 0C
 A9 04 58 F1 A1 8B 9E 8E D7 6D F8 33 59 33 30 64
 FC 7E 49 F3 12 24 7F 3E 8D F7 93 09 FE B3 A6 78
 63 CC DF F6 FB 20 59 0E 90 AA CE 64 3F 1B 45 5D
 14 10 86 AB F1 34 33 2F A2 56 F1 AB 29 F1 33 9C
 02 69 32 6B 8C B6 05 D5 D8 2B 1D 34 64 5F BB 51
 CB 81 07 C4 4B BA 69 C5 D7 7A 4C 2A 1F FC A2 E6
 79 52 07 7B 9B 55 9A 6C 29 70 47 93 F3 8C 92 17
 1F 98 CB 2A 90 6C 56 0E 53 89 3B 03 8F B4 9A E9
 47 4F E8 2E 74 07 5F BA 9C 22 C4 32 BE 66 C2 2D
 A7 52 54 4F D6 70 37 15 F3 5A CD 0F A5 12 56 1C
 B7 EF 09 69 8F 94 BA 72 C3 6A 6B 6B B2 72 E8 D6
 24 3C 7C CC 61 C5 DD E1 44 95 47 16 DF DB F5 13
 22 31 7D ED 55 93 09 4D 32 B8 FC 5A 48 FC 4A 5D
 22 47 8C CA 89 63 B5 6F F8 B7 79 A6 4D 71 17 1A
 6D A0 F4 8A 0A 57 59 BD D0 69 E4 3A 57 77 AB 5D
 07 44 34 C2 4A BE C6 35 99 EE 21 77 A4 E7 44 EE
 43 6D 22 2D 5D 05 4A 0C 4D C3 A4 5E 3E 97 A6 92
 AA 73 13 FE DF FA 9B B8 C9 F6 33 52 A1 B1 5D 72
 BD 1D 5C 63 79 5F 5A 89 B2 FA 10 30 49 FF D9 19
 8F 55 DF 44 29 F3 81 90 5B FA B8 83 67 BA 66 AC
 DB 69 E5 96 0C CE DE BB 61 2C F0 DA C7 8D 0B BC
 6B 9B 3D 06 D8 DC 4D 24 50 CF EC 3C 78 BB F4 A0
 2C 28 32 A4 68 F5 3A AF 8D 1E 9D 44 E4 4B 8A 50
 87 7A 9B EF 02 2B 1D B2 B8 38 AB 78 B5 F6 64 64
 A9 E0 40 87 2E 81 6C 0B 22 3F 41 E4 57 DF 27 5D
 7D 21 D3 83 74 55 4F CB A3 2A FB 71 80 64 22 F2
 5D 07 DC A5 DF 0E 29 CB 7B B8 AD 4B AF 9F 03 1E
 B3 67 46 EA 6A B7 D9 2D CA B7 CD B9 DE A5 51 D4
 07 BA 95 7C D2 94 15 E3 1A AC F0 0A FC 2A FA 21
 37 A7 20 23 4D 9A 59 2F 79 62 38 82 63 B4 95 83
 F8 6F E1 B0 75 F0 45 5B DF B3 BF B4 AC F8 30 0E
 5D 4A 2B A3 7B 35 6B 81 62 CF 2C EF BA 59 7E 60
 5A A3 12 33 B9 3D 17 BC 03 3F 40 ED 12 B7 46 6B
 27 9D 39 7C 5E 18 3B 75 79 8D D1 61 37 6C 35 AE
 45 B5 18 2C E3 46 72 0A EE 4F 3F F6 BC A6 F6 D2
 7F 0C 56 03 3C 78 C0 7F 30 93 BA 9E 85 7E C1 24
 45 97 D1 41 EB DC 2E 00 D8 03 EE 35 2A 6D CC 1C
 60 F7 AD 57 5F DF 4C 65 A6 B7 B6 2E D9 EC 67 9A
 C4 EF 93 A2 2C 7F 00 B8 15 49 B0 56 52 79 9C 02
 83 81 E6 D7 C7 E1 47 58 00 8B 21 31 12 52 D6 75
 BF 6B D7 56 1D 2E 46 F9 42 B9 8D 4F D1 07 9A 16
 6B 18 83 CD 97 D0 8B 53 3B 88 A2 92 FC 4D 10 10
 70 0F CC F1 6A 68 FD 4E 00 42 7C 8F B2 8F 9A C5
 9E 0A 91 88 31 23 54 C7 F7 AF 26 2C 37 61 8D B6
 5A 1E B7 E0 BF 5C DE 07 18 00 DA 32 FF BE 79 4C
 43 34 D4 41 FC 1A 0D AA 5D 46 6D FE AF F6 78 F9
 B1 BD 89 CA A6 DA 0E B8 69 01 AC 6E 26 3F C9 E7
 1F AA A7 8E BE 66 ED 7A E2 D0 28 44 42 2C 6B A2
 7F 38 EA B3 7D D2 E6 49 59 88 3C 7A B6 59 05 D7
 0E 17 63 1F 7A DA C5 B1 E4 AE 5C 81 35 54 18 34
 E3 47 B9 1D 86 6B FC F0 DF D0 75 40 89 7B AD B6
 B3 FA 10 B2 8A 67 E0 32 24 5F BE 70 42 81 FB 15
 0E D9 D9 EA 3B 3D 1F A7 AE 16 0E 4C 68 6D 5D 6A
 6B DB 44 10 F1 11 06 9B D5 4F 80 33 CA 0E 5E 1D
 A0 EF AE BC 04 E9 73 1C 43 53 FD A2 B9 E6 CF 3E
 C6 4F DC 9C 52 D5 BD 5C F1 A0 3F A0 B6 92 71 B1
 3B C8 FE D4 46 36 F6 52 1A CB 0F 69 17 06 67 47
 49 DD CD 49 CE 52 19 36 72 0C 34 A4 CE FD 8A 5B
 CB 77 60 FF CB BE 8F 60 AC 64 94 9E D4 D3 0F B6
 75 CB 91 4C 43 F3 5F 9D 7A C3 9A 3B 16 66 C1 F6
 69 3B 47 02 AE FE C9 B7 47 DC 5B 85 EA 39 6E 0D
 3A 30 79 D0 BD 69 C5 17 C7 5E 31 51 78 A4 D8 88
 88 83 AE 57 58 AE 12 67 B7 F5 85 3E 92 65 64 50
 0C 11 0A 12 8B 96 F8 58 9D 79 3A 3E 1F 54 A7 3B
 7E F1 C6 67 6D 29 52 7A D8 17 2D 71 F8 95 83 83
 CB E8 82 7E AA AD 92 8F 28 27 79 19 E8 E8 F4 35
 EE 75 21 7E F5 3B A2 CE 9F 91 78 82 A9 5C 3E DC
 84 06 CE F4 54 54 9C FD 60 08 13 23 A8 25 2A 89
 E7 31 FC 01 A0 49 87 F2 D4 49 9C BD 10 B9 B1 B9
 6A 4F B6 E5 55 3D B7 C0 56 1A BB 5B 76 31 F2 D3
 D6 FA 70 97 E3 D9 F0 19 BA 2A 05 A6 88 AA 55 ED
 70 0C 63 70 CD AB 5F D7 C8 C9 9B 01 16 4B 9D ED
 FC 30 97 7A 73 35 31 3A A7 FF 17 81 E0 59 DE 6A
 37 4D E7 F6 C4 DA A3 E5 E8 58 60 0E 2D 08 BF D0
 0F F1 49 64 CD 84 83 08 29 38 AB 18 A0 37 A7 46
 35 67 05 ED 0B 4F 42 94 31 2E 76 A3 B1 34 F9 9F
 4A 4D 58 FE 44 15 98 F0 DC FA A2 49 D0 41 66 4B
 F9 F7 A7 D5 FE BF CD 9F B4 A9 73 74 FC BD CC F0
 24 1F BE BF D7 07 0E 41 B5 EF 09 1D FF 0A 24 11
 DB C4 1B 91 59 E6 04 3E B0 B4 83 5B 4E 6F 76 91
 35 88 CF 8F 59 17 9A 19 55 F0 A7 60 43 85 39 3F
 8A 64 5C 67 DF 5A 3B F5 ED 3D 9C FB 19 50 9F EC
 B6 25 B7 40 3C BB 41 6C FC 6C AA B6 6F 6E 78 B3
 C5 35 FD 77 8F 85 7D EB C5 01 12 0F FA 76 47 97
 7A CF 55 E9 97 85 8A FC 45 34 73 13 29 03 C3 FA
 AB 99 07 7B B0 E7 A4 C3 75 CF 23 5E A7 D0 EB 84
 C6 5F 6C 4E F3 19 4D 9F 7B B5 D8 38 43 29 8E 3A
 5A CE 52 4D 08 49 05 8F 54 5F 13 AE 4D 88 FC AA
 71 AD 86 80 8C 80 07 C8 FA FE C7 18 C4 C3 F4 26
 BA 7E 44 E1 6D 3E 60 9D 20 0D A4 E6 92 46 0F 4F
 1C BF 73 37 03 72 02 DB 9C 69 D2 67 2B 05 72 25
 93 72 F9 1B 9E 3D E8 17 03 3C 5E 2E C7 A9 CC 4C
 9C 08 FB 65 C3 A3 60 47 8A 52 C3 F0 F3 02 AB B8
 37 69 EC CF D8 DB 6F A7 6E 42 7D DC 91 E4 12 A5
 EA 26 43 50 19 88 67 CB 29 04 E4 2F 53 E4 12 50
 C0 D2 17 57 1A 95 45 FE 0B 2C 66 B0 B1 D0 FB 20
 F2 E6 22 66 E3 5C 34 D5 11 35 2E AD EF 4B 54 A5
 FC 57 9B 6C 36 2C 62 54 55 B9 86 C2 86 42 91 2D
 AD A2 8B E8 B0 94 E0 92 09 CC F8 07 0D C5 B6 18
 74 84 14 B0 6C 8F 1F 68 C1 F6 4F 75 36 58 E1 8A
 7F 97 3C 5E 04 25 6A 87 37 0E 56 06 8E 37 3C 88
 50 F4 3D 60 8D FF DD A1 8A 69 47 94 60 F5 E0 47
 34 24 B3 15 47 9E 52 5C F1 91 D3 D8 72 AA 5B 24
 84 57 16 B7 10 51 00 A3 A3 D2 FC 6A 8C 19 D9 AB
 37 51 C0 55 F7 DF 06 EE 59 3E 0D 4D A8 E2 35 3C
 B9 90 4D 0B B6 CF 75 0A 3E C6 E3 F5 B5 1C CD BC
 63 80 5A E5 D6 1D A2 21 24 B5 8A 4E F0 D4 CB DB
 34 6D 2A 21 5F 86 92 0C BF D7 17 A1 E0 34 F0 B7
 74 2D B7 54 BA E1 A3 5C 14 B8 00 40 D3 81 4B D3
 C7 F3 5A C7 4C 26 62 46 71 43 68 A4 43 3E 75 09
 15 71 84 24 C7 2A D8 51 08 55 DF E3 B1 D5 A6 9B
 6B DB 82 33 0F 51 EF 9B 6E 6E 99 6C 52 00 B3 47
 68 6A 79 50 48 E6 F6 1A EA A4 79 36 02 B5 8F 99
 A8 42 87 44 21 A3 80 CE F1 A7 9E 7B 3B B9 4E 2A
 4D A4 42 C6 4A FB 8E DA A2 0A B6 35 E2 75 47 37
 31 33 55 96 B3 CB 60 DC 02 E8 AF 53 EF 5E 48 CE
 33 6C 44 78 80 84 67 DE 85 B5 A7 44 C9 D5 EC DD
 49 AE F2 90 5F 2E A2 EB D2 70 39 34 65 EE CF 0F
 91 EB 48 BB 94 14 B5 49 31 48 94 52 9D 78 54 AE
 89 1A 80 0B 7A 08 9F FA 21 59 84 40 41 AE 4A A4
 24 68 8D 33 B1 97 F9 E2 00 95 B1 A2 9B 00 BC C9
 C3 F4 04 18 83 0B 18 39 22 C1 AD E4 4A AC 5E 7D
 91 A7 29 4F 41 7E 52 F4 12 4D E6 8C 9F DD F9 86
 13 43 8B 71 71 DD 36 03 2E 30 B5 25 36 1B 43 FE
 A0 2E 6B AC 62 CB 23 79 41 A2 F4 9A 42 25 19 B8
 EF 0B EE 23 F3 BF 61 1C BA E6 9D 3D C5 F9 09 A2
 24 E8 DF 88 4E DA 48 7A 23 BB 1F 26 24 8A 73 6E
 65 45 CF 39 5B E7 8C F0 40 FD 4A 43 94 AA 29 78
 7E 26 72 82 94 75 E7 0A DB CF 17 9D EB 16 40 B6
 C1 33 A3 24 B1 F4 85 5A 6E 24 16 78 B7 4A A9 30
 8A 05 CD 3B 38 16 ED D6 05 F5 3D 46 6D 36 B5 27
 6F 34 D9 8B 0A D3 09 84 E8 2A 96 8B 4A 79 6F A5
 42 1F 4F D1 44 56 CB A1 22 8D 31 56 87 3D F7 39
 DE 9E 89 2F B6 96 48 BD 51 FD E4 00 57 B0 C8 14
 F4 EF 2D 0D 00 F5 0A 8F E3 FF 0D DA 8E AD 53 1D
 29 17 32 32 8B E7 B4 C1 66 BE 3D 0C 0F 8F 93 94
 BB F8 C7 13 3B D2 C0 BE 1F 04 76 84 3D 0C FE 6B
 46 06 23 9A AB C5 95 02 E1 61 B9 1F D4 DE 45 18
 37 25 EC 9E 20 91 36 09 63 22 52 CB F2 5C 6A AD
 AB 9E 93 C6 D1 7F 75 A9 94 A4 BA EE E1 5D 96 60
 3C 32 C2 53 1A 39 39 02 F9 9F 72 7C 16 80 B6 80
 10 77 7B 87 54 DB 8C 71 C0 50 00 9A F4 BF 21 7F
 2E 56 1D A0 0E F6 CE 2D 9F 73 07 18 B3 F8 82 E9
 11 96 38 D7 02 DB 9B 12 3F D3 BC A2 49 93 40 C3
 12 B2 FC 16 AD 6A 41 A1 E0 56 6A AE F7 36 79 0F
 AA 53 01 0B 0A 3D CC D6 A8 D5 98 6D 52 B2 DF 8B
 6B ED F8 16 49 1F 61 79 1C 64 44 1E 1B 48 1F 50
 DE 7A F9 93 CE C4 12 05 31 F4 6F 6C FF 3B 4C 54
 FD A4 E5 63 8A B8 83 5A 00 2B 41 F2 E1 73 72 4C
 57 3E 22 3A 4F CB D3 56 65 BF 33 7A EC CE 5A AA
 38 A4 77 61 97 CF C4 4D 98 29 93 C9 D6 90 16 D4
 87 E3 DA 01 79 FB AF 12 C7 05 B0 7F 6F 92 D9 98
 90 02 D8 89 BD 3A 84 55 C9 05 B7 C2 D6 0F 5D F6
 31 81 67 D9 B3 5D E7 0F 10 87 05 6C 83 8B 0D B1
 EC DE 26 DB 45 B3 93 94 EF 3A 8B 7A AB 47 E9 98
 CD E4 71 7B A0 A0 27 13 10 56 C3 0F FD 8E BB B9
 B6 DF 63 BE DD D3 F1 92 44 21 8B 13 F0 84 7D 4F
 07 50 C0 0C 5F 2F 7F 62 59 02 3D 99 F6 26 94 91
 5A A9 4A BD 1C 57 AE BE 40 7E 5C 40 D9 CC 8E 4F
 C8 EA 52 F2 D7 D7 98 0F 9A D4 5B B6 70 C5 2D F2
 E7 C9 5F A9 AF B7 FA C4 BF 9C 4F C1 25 2D B3 9E
 8C E2 7D 14 47 80 D9 AC B8 01 B2 87 66 89 91 9F
 C5 0D 2F 46 D1 68 4D B1 F2 B2 A8 CE FD 00 99 DB
 2F 99 28 02 9B 54 09 6E CC F0 9A 24 CA DB 2A 5E
 B3 11 1D 15 95 25 D2 F7 9D 9B 67 B5 ED 90 BD 00
 96 57 42 ED D9 E8 BB 7A A8 99 9D 26 F5 63 22 25
 3B 55 85 7F 5F 10 6C FF 7A 13 BB 30 BE 48 17 15
 A9 FE 70 71 76 53 0A C9 9C B3 D1 F4 C8 82 DA E2
 EB 49 17 06 FD DC 0B 83 68 A8 3D EE 72 48 F7 89
 D1 A3 D5 82 C2 DB EB C0 D0 0D D0 11 21 8E 74 B4
 13 90 E1 45 4A 8E FD 0F A0 8D 3C 1E 93 97 A8 DE
 F6 DC FF D2 91 E9 9D 4F 78 4E 73 94 CA FB 27 32
 E6 04 E2 43 81 3B 55 A5 CC 86 A0 D5 68 04 CD C9
 F3 50 8A FE 19 AD 4E D2 64 23 30 48 64 19 0E DD
 53 E1 59 A1 57 B3 69 2A EF EA 2B D0 E8 08 B4 35
 B0 E9 09 A0 2C 4C 83 99 D7 DD D3 EC 66 35 36 16
 68 3A 76 8F 25 3F 0F AF B3 B6 E5 89 1E 1D 4E 01
 35 A5 ED 6E 15 EF BF 41 FB 28 65 79 F8 E0 84 45
 89 E5 70 AA 62 77 3A 19 F4 9D 9B 57 D4 1C A7 61
 B2 73 31 A4 D2 D4 52 FD 04 82 EF 78 33 15 64 82
 36 DC 7D 30 B9 16 E2 82 07 F8 8F 46 1A 3D 8C 6D
 C5 71 47 7B 06 CD 04 46 C0 A8 3D 80 02 0F D8 05
 03 50 B1 3F B4 88 C0 40 EF 39 2F A5 46 C5 65 2E
 F7 24 2A 41 D6 45 8C 0C 4F 76 A7 6B 29 C0 B3 96
 01 E5 25 55 84 85 9B 04 FD 91 20 C5 B4 D2 1F 63
 75 00 4A 63 6C A5 6E 60 2D B5 25 B2 FF 00 8F 08
 B4 86 7E E0 08 CD 21 05 A1 C7 FE FC 81 BA A9 28
 AB 76 1C 09 83 BD 90 C6 CD AC A4 AB 27 2A 67 2F
 9F CB 2A 67 C1 A4 AB CD 3E 0C D6 22 75 85 50 79
 76 3C 56 3E 86 56 E9 7B EA 54 3D 6D BE A7 23 87
 E8 94 D7 00 20 49 1D 1E C2 25 BA FA BE 55 8C C8
 31 53 48 0F 4D D3 C1 D9 D8 1E 21 32 D6 75 F8 49
 E7 D6 6E 91 C1 0E 38 ED 26 06 2C 2F B3 B7 2A 65
 5D B6 11 7C 4A EC DD 74 9E CF 87 68 28 61 72 B1
 D7 76 CE B1 E4 28 61 C3 20 17 F6 71 7E D8 C7 BB
 DB 9C 13 28 9A BB 45 40 88 46 A3 2C 82 49 0E E8
 CB A4 8B 3B BB E7 36 17 B9 82 D5 5A 6C B2 4A 1F
 C9 9A 8E 3E B2 46 87 C9 A8 5E 20 9E 72 10 A9 13
 68 26 E9 6B 19 A1 2F 7B 74 B4 92 D4 B1 03 CB 16
 B0 9F 19 E9 18 7A 78 1F AC EE F1 B3 EC 32 38 AD
 A9 85 43 91 9B 7F E8 EB 91 75 F0 37 55 0F 78 EE
 B9 6A 74 A3 72 BD 04 35 54 C7 F9 26 E1 99 0C DD
 35 91 D2 4E 25 6F 72 6F 7D AC 41 DA 47 89 14 51
 D1 E8 A0 17 08 2E FB 0C F6 08 83 4B 6D FA 2C 2C
 FA E9 01 DE EB C1 D0 72 08 25 E1 29 B0 52 8F 85
 9C 1B 86 FB CE 59 FD 7C 41 19 A9 E8 03 5D FE 03
 A1 C6 9D 98 3A 3E 7B C0 C0 35 ED 42 D5 36 7A BC
 39 B1 D2 AA 54 84 89 14 2C 48 52 84 9C 34 5D CB
 B6 7F CD 45 E9 54 51 A7 58 31 B0 04 E6 24 79 67
 3D 57 A1 03 A4 D2 75 FA F2 EA 6F C1 17 D2 9E 83
 AD 28 9C F2 08 61 18 B1 7B 80 AC 58 D6 BC 99 AA
 E9 35 C4 F4 2E 56 5B 1B 45 24 C5 C2 A0 19 F7 73
 35 BC 09 3C F5 1A 38 7D 8B FF AD 1B 67 E7 BA CE
 B6 82 98 C2 C3 1C 10 6B CE A1 EB FB E9 D9 B3 B0
 D9 A8 95 75 93 89 5E 83 2A 69 E9 2B EB 0F 72 E8
 2F 92 23 7E 9E 10 FE A4 71 B9 20 64 83 CF 02 78
 46 C7 93 89 93 BE 64 01 D0 DB 9B 3B 78 D2 AA BF
 80 A5 C8 93 A1 96 68 13 D9 C8 94 93 A7 26 02 EF
 AE EB C3 2C C9 05 F4 23 87 F9 52 15 E5 72 CF 99
 36 60 C9 D4 CE CF CE B7 1F AA D4 29 BE 91 92 29
 BB E4 A4 D4 9D A6 8D 4A 67 8D F6 95 D7 B6 3A 39
 28 18 DF 6B 5D E7 AC C9 97 29 5F 6F 9F 32 F3 0F
 AB 06 3B 91 FA 1A 4B 06 D5 CC 2E 2D BF CA 80 2A
 F9 6E 6B 5A 55 3C 5B ED 49 78 C2 74 00 BC 4D 9B
 17 09 BD 0C D4 D0 C2 DC 27 4B 52 07 91 EC 40 C9
 3F A7 5E 2A 22 AF A2 04 75 8C F7 3D F9 95 05 E6
 64 71 CB CC A9 99 BC C1 9D 14 BD DF E2 BB 20 DE
 FF 53 62 56 C7 15 BA C5 5F EE D8 AF D2 48 56 4C
 95 0C 63 A7 08 98 F8 D7 5D CC 54 F7 F1 1E F7 4D
 80 EA 38 89 43 22 19 06 2D 14 1C 87 95 E9 C7 E8
 FE 03 E9 1F 04 97 DD 55 F4 69 2B FC 9D E1 17 DB
 ED BD 3C E2 0E 2E B1 B9 17 56 59 37 E3 A2 49 33
 38 9A 03 F7 85 87 DE EE 37 18 1D C3 19 56 6C D8
 BA 84 CB F9 75 29 F8 87 A1 0C 61 8C 1E 66 00 86
 2D 8B 4B 58 CC AE F6 B6 A9 83 FB 5F 4C BA 01 B5
 E5 4A 22 DE 74 B9 8B BC 2A ED 58 E0 D3 39 BA 29
 A3 4E 89 1A 39 7B 11 EC D6 3A CC 54 8F 85 E8 69
 5C 20 BD E1 C3 EB E5 ED 5A E8 AE 19 EC 10 03 B0
 DD 62 70 F5 B3 CA 7F 6B 06 AE D4 95 2C B6 98 2C
 7A D3 4A D3 1F CF DA 74 55 13 60 E4 6B 82 28 13
 F6 ED 6E DD 19 C1 0A 1E F1 2F 8A 15 6D C2 31 38
 08 38 EE E2 D3 94 CE B0 BE 60 1B 9E 7D 03 BC DF
 8F EE B5 81 33 9A E3 60 6D EA E8 16 B9 FB 57 BE
 7F B7 CF 9F 8D 3C 31 9F 34 B5 D5 07 3D 57 DA 6E
 03 0E 9C CC 5F F4 66 EE 0D 9B 95 38 BD 83 09 90
 B5 14 12 C3 73 1C 72 13 FA B6 D0 B7 18 E4 46 03
 7A C6 A4 EA 48 86 01 D1 B5 95 E5 47 CA 67 70 31
 1C 0E 73 AE E3 B1 60 45 D4 DC 77 4A 73 F4 A7 B4
 2D 87 6C A6 04 C1 3B C8 1C 60 F7 89 3C 38 32 59
 AB C4 1B 86 CD C4 DC 03 AB 32 81 A3 2E C5 E7 8C
 87 59 D9 60 00 BA BB 80 F7 0F F2 5C 63 42 FB 32
 C7 67 01 BB 94 8A EC 56
* End 77536280 4213765698