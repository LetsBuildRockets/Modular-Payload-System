.SUBCKT T521D475M075ATE075 1 8
*Temp = 25°C, Bias = 0VDC, Center Frequency = 10000 Hz
*KEMET Model RLC Tant5RC
R1 2 3 0.0234496109187603
R2 3 4 0.00891980528831482
R3 4 5 0.00891980528831482
R4 5 6 0.00891980528831482
R5 6 7 0.00891980528831482
R6 2 8 2128000
L1 1 2 2.29999996825825E-09
C1 3 8 1.51612903225806E-07
C2 4 8 3.03225806451613E-07
C3 5 8 6.06451612903226E-07
C4 6 8 1.21290322580645E-06
C5 7 8 2.4258064516129E-06
.ENDS