.SUBCKT T521X226M063ATE075 1 8
*Temp = 25°C, Bias = 0VDC, Center Frequency = 10000 Hz
*KEMET Model RLC Tant5RC
R1 2 3 0.0139982542023063
R2 3 4 0.00546912709251046
R3 4 5 0.00546912709251046
R4 5 6 0.00546912709251046
R5 6 7 0.027345634996891
R6 2 8 454500
L1 1 2 2.80000000962843E-09
C1 3 8 7.09677419354839E-07
C2 4 8 1.41935483870968E-06
C3 5 8 2.83870967741935E-06
C4 6 8 5.67741935483871E-06
C5 7 8 1.13548387096774E-05
.ENDS